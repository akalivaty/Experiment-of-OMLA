//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n462), .A2(KEYINPUT69), .B1(G567), .B2(new_n458), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n468), .A2(new_n469), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n476), .A2(new_n469), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n476), .B2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n467), .A2(KEYINPUT71), .A3(new_n470), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(G136), .B2(new_n494), .ZN(G162));
  NOR2_X1   g070(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n497), .C1(new_n474), .C2(new_n475), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n498), .B2(new_n482), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n497), .A2(G138), .ZN(new_n500));
  INV_X1    g075(.A(new_n496), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n467), .A2(new_n469), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n467), .A2(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n499), .A2(new_n502), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  AND2_X1   g098(.A1(new_n517), .A2(G89), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n513), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AOI22_X1  g108(.A1(G51), .A2(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n526), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n518), .A2(new_n539), .B1(new_n520), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n518), .A2(new_n545), .B1(new_n520), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n530), .B2(G53), .ZN(new_n560));
  AND2_X1   g135(.A1(KEYINPUT6), .A2(G651), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT6), .A2(G651), .ZN(new_n562));
  OAI211_X1 g137(.A(G53), .B(G543), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n558), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n530), .A2(new_n559), .A3(G53), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n511), .B2(new_n512), .ZN(new_n571));
  AND2_X1   g146(.A1(G78), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n513), .A2(new_n517), .A3(G91), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n569), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n530), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n518), .ZN(G288));
  AOI22_X1  g157(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n515), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n518), .A2(new_n585), .B1(new_n520), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT76), .ZN(G305));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n518), .A2(new_n590), .B1(new_n520), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n593), .A2(new_n594), .B1(new_n515), .B2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n513), .A2(new_n517), .A3(G92), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n513), .A2(G66), .ZN(new_n600));
  INV_X1    g175(.A(G79), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n527), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n597), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT78), .ZN(G148));
  NOR2_X1   g189(.A1(new_n550), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n605), .A2(new_n612), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT79), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n615), .B1(new_n617), .B2(G868), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n467), .A2(new_n471), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2100), .ZN(new_n624));
  OAI221_X1 g199(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n625));
  INV_X1    g200(.A(G123), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n488), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(G135), .B2(new_n494), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n623), .A2(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(G2096), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n624), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT80), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n656), .B(new_n653), .C1(new_n649), .C2(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n649), .A3(new_n651), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT81), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n665), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  NOR2_X1   g255(.A1(G6), .A2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n588), .B(KEYINPUT76), .Z(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G16), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT32), .B(G1981), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G288), .B(KEYINPUT84), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G16), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G16), .B2(G23), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT33), .B(G1976), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(G1971), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AND4_X1   g272(.A1(new_n685), .A2(new_n691), .A3(new_n692), .A4(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT82), .B(G29), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n494), .A2(G131), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n487), .A2(G119), .ZN(new_n706));
  OAI221_X1 g281(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT83), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n710), .B(new_n712), .Z(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G1986), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(G1986), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n700), .A2(new_n701), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT85), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G29), .B2(G32), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n487), .A2(G129), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT26), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n729), .A2(new_n730), .B1(G105), .B2(new_n471), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n494), .A2(G141), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n723), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n734), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n738), .B2(KEYINPUT88), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n702), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n487), .A2(G128), .ZN(new_n746));
  OAI221_X1 g321(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G140), .B2(new_n494), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n745), .B1(new_n749), .B2(new_n735), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2067), .Z(new_n751));
  INV_X1    g326(.A(G2072), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n494), .A2(G139), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(new_n469), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n735), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n735), .B2(G33), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n751), .B1(new_n752), .B2(new_n761), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n742), .A2(new_n743), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT24), .B(G34), .ZN(new_n764));
  AOI22_X1  g339(.A1(G160), .A2(G29), .B1(new_n702), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2084), .ZN(new_n766));
  NOR2_X1   g341(.A1(G5), .A2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT92), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G301), .B2(new_n693), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n628), .A2(new_n703), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT91), .B(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n766), .B(new_n779), .C1(new_n752), .C2(new_n761), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n703), .A2(G27), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n703), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2078), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n551), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT86), .B(G1341), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n693), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G168), .B2(new_n693), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT89), .ZN(new_n790));
  INV_X1    g365(.A(G1966), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n783), .B(new_n787), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n605), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1348), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n785), .B2(new_n786), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n780), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(G162), .A2(new_n703), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G35), .B2(new_n703), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT29), .ZN(new_n800));
  INV_X1    g375(.A(G2090), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT93), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n790), .A2(new_n791), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT90), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n763), .A2(new_n797), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n719), .A2(KEYINPUT85), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n718), .A2(new_n720), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n693), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n609), .B2(new_n693), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1956), .Z(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n801), .B2(new_n800), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT94), .Z(new_n814));
  AND4_X1   g389(.A1(new_n721), .A2(new_n806), .A3(new_n808), .A4(new_n814), .ZN(G311));
  NAND4_X1  g390(.A1(new_n721), .A2(new_n808), .A3(new_n806), .A4(new_n814), .ZN(G150));
  NAND2_X1  g391(.A1(new_n605), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  INV_X1    g393(.A(new_n518), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n819), .A2(G93), .B1(G55), .B2(new_n530), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n515), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n550), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n550), .A2(new_n822), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n818), .B(new_n825), .Z(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n827), .A2(new_n828), .A3(G860), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n822), .A2(G860), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(new_n628), .B(new_n484), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G162), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n836));
  INV_X1    g411(.A(new_n749), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n737), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n509), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n499), .A2(KEYINPUT95), .A3(new_n502), .A4(new_n508), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n734), .A2(new_n749), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n838), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n843), .B1(new_n838), .B2(new_n844), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n836), .B(new_n759), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n759), .A2(new_n836), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n845), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n708), .B(new_n621), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n494), .A2(G142), .ZN(new_n854));
  INV_X1    g429(.A(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n482), .A2(new_n855), .B1(KEYINPUT98), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(KEYINPUT98), .B2(new_n856), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT97), .B1(new_n487), .B2(G130), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n487), .A2(KEYINPUT97), .A3(G130), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n854), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n853), .B(new_n861), .Z(new_n862));
  AND3_X1   g437(.A1(new_n848), .A2(new_n852), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n848), .B2(new_n852), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n835), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n848), .A2(new_n852), .ZN(new_n866));
  INV_X1    g441(.A(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n848), .A2(new_n852), .A3(new_n862), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n834), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n865), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(G299), .B(new_n604), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT41), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n874), .B2(KEYINPUT41), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT79), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n616), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n823), .A2(new_n882), .A3(new_n824), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n823), .B2(new_n824), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n617), .A3(new_n883), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n877), .A2(new_n879), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n874), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n888), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT103), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n888), .A2(new_n886), .A3(new_n890), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n888), .A2(new_n886), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n878), .B1(new_n875), .B2(new_n876), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(G303), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n682), .A2(new_n686), .ZN(new_n900));
  INV_X1    g475(.A(new_n686), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G305), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n899), .B1(new_n902), .B2(new_n900), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n900), .A2(new_n902), .ZN(new_n908));
  XNOR2_X1  g483(.A(G290), .B(G166), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT101), .B1(new_n910), .B2(new_n903), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n898), .B(KEYINPUT42), .C1(new_n907), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n903), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n906), .B1(new_n904), .B2(new_n905), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n910), .A2(KEYINPUT101), .A3(new_n903), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(new_n898), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n892), .B(new_n897), .C1(new_n916), .C2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n897), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n919), .A2(new_n898), .B1(new_n914), .B2(new_n913), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n907), .A2(new_n911), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT102), .B1(new_n924), .B2(new_n914), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n926), .A3(G868), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G868), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n822), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n921), .A2(new_n926), .A3(KEYINPUT104), .A4(G868), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(G295));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(G331));
  AOI21_X1  g509(.A(G168), .B1(G301), .B2(KEYINPUT105), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n937));
  NAND2_X1  g512(.A1(G171), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n823), .A2(new_n824), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n823), .B2(new_n824), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n823), .A2(new_n824), .A3(new_n938), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n935), .A3(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n877), .A2(new_n879), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n944), .A2(new_n890), .A3(new_n941), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n924), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n917), .A2(new_n918), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n941), .A3(new_n890), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n944), .A2(new_n941), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n948), .B(new_n949), .C1(new_n950), .C2(new_n896), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n951), .A3(new_n871), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n944), .A2(new_n941), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(new_n875), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n949), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n955), .B(new_n924), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n871), .A4(new_n951), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n954), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n953), .A3(new_n871), .A4(new_n951), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(G397));
  XNOR2_X1  g544(.A(new_n749), .B(G2067), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT107), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n737), .ZN(new_n972));
  INV_X1    g547(.A(G1996), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n842), .B2(G1384), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n472), .A2(G40), .A3(new_n483), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n976), .A2(G1996), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n737), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n708), .B(new_n712), .Z(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  AND2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT114), .B(G8), .Z(new_n989));
  OR2_X1    g564(.A1(G102), .A2(G2105), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n507), .A3(G2104), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n503), .B1(new_n474), .B2(new_n475), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n467), .A2(new_n469), .A3(new_n500), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n496), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n995), .B2(new_n502), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n472), .A2(G40), .A3(new_n483), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1981), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n588), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n584), .A2(new_n587), .A3(G1981), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n998), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G288), .A2(G1976), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n998), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT45), .B1(new_n509), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n977), .B1(new_n1010), .B2(KEYINPUT108), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n840), .A2(KEYINPUT45), .A3(new_n1009), .A4(new_n841), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n696), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n509), .A2(new_n1017), .A3(new_n1009), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT109), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n509), .A2(new_n1020), .A3(new_n1017), .A4(new_n1009), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n509), .A2(new_n1009), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n977), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT110), .B(G2090), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1016), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(G166), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT113), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1016), .A2(KEYINPUT111), .A3(new_n1026), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1029), .A2(new_n1036), .A3(new_n1037), .A4(G8), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n998), .B1(new_n901), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n998), .B(new_n1042), .C1(new_n901), .C2(new_n1039), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1005), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1008), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT63), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1035), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1024), .A2(new_n1018), .A3(new_n1025), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1016), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1051), .B2(new_n989), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1044), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1038), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G2084), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1022), .A2(new_n1055), .A3(new_n1024), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1023), .A2(new_n975), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n997), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n791), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n989), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(G168), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1046), .B1(new_n1054), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1029), .A2(G8), .A3(new_n1037), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1049), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1046), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1038), .A3(new_n1053), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1045), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  INV_X1    g645(.A(G2078), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1057), .A2(new_n997), .A3(new_n1071), .A4(new_n1058), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n1072), .B2(KEYINPUT120), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1010), .A2(new_n977), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1071), .A4(new_n1058), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1073), .A2(new_n1076), .B1(new_n770), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1011), .A2(new_n1013), .A3(new_n1071), .A4(new_n1014), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1070), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1079), .B2(new_n1070), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G168), .A2(new_n989), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1085), .A2(G168), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1033), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT51), .B1(new_n1090), .B2(new_n1086), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1084), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1038), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1069), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1079), .A2(new_n1070), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT121), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1079), .A2(new_n1080), .A3(new_n1070), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1077), .A2(new_n770), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT122), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1077), .A2(new_n1108), .A3(new_n770), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1070), .B(G2078), .C1(new_n977), .C2(KEYINPUT123), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n977), .A2(KEYINPUT123), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n976), .A2(new_n1014), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1105), .A2(new_n1110), .A3(G301), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT54), .B1(new_n1114), .B2(new_n1084), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1115), .A2(new_n1054), .A3(new_n1092), .ZN(new_n1116));
  INV_X1    g691(.A(new_n568), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT75), .B1(new_n566), .B2(new_n567), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n575), .B(KEYINPUT57), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n573), .B(new_n574), .C1(new_n560), .C2(new_n564), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n569), .A2(new_n1120), .A3(KEYINPUT57), .A4(new_n575), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n997), .A3(new_n1018), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT115), .B(G1956), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  AOI21_X1  g712(.A(G1348), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n997), .A2(new_n996), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(G2067), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1140), .B1(new_n1077), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n604), .B1(new_n1143), .B2(KEYINPUT60), .ZN(new_n1144));
  NOR4_X1   g719(.A1(new_n1138), .A2(new_n1137), .A3(new_n1140), .A4(new_n605), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1011), .A2(new_n1013), .A3(new_n973), .A4(new_n1014), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1139), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n550), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1151));
  XNOR2_X1  g726(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1136), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1126), .A2(new_n1133), .A3(new_n1128), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1143), .A2(new_n604), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1126), .B1(new_n1133), .B2(new_n1128), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT119), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1153), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1105), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(G171), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1083), .B2(G171), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1105), .A2(KEYINPUT124), .A3(G301), .A4(new_n1078), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1163), .A2(KEYINPUT54), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AND4_X1   g742(.A1(new_n1116), .A2(new_n1159), .A3(new_n1161), .A4(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n988), .B1(new_n1101), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n978), .A2(new_n985), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT48), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n709), .A2(new_n712), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n982), .A2(new_n1172), .B1(G2067), .B2(new_n837), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n984), .A2(new_n1171), .B1(new_n1173), .B2(new_n978), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n980), .A2(KEYINPUT46), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n972), .B2(new_n978), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n980), .A2(KEYINPUT46), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT126), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT127), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT47), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1180), .A2(KEYINPUT47), .A3(new_n1182), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1174), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1169), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g763(.A1(G229), .A2(new_n465), .A3(G401), .A4(G227), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n966), .A2(new_n872), .A3(new_n1190), .ZN(G225));
  INV_X1    g765(.A(G225), .ZN(G308));
endmodule


