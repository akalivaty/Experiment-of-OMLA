//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT71), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n206), .A2(new_n207), .B1(G183gat), .B2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(KEYINPUT28), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT27), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n212), .B2(new_n214), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G183gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT27), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n209), .B1(new_n213), .B2(KEYINPUT27), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n222), .A2(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n218), .B1(new_n227), .B2(KEYINPUT69), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(G183gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n223), .B1(new_n229), .B2(KEYINPUT27), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT69), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n225), .A2(new_n226), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n208), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT72), .B(G120gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G113gat), .ZN(new_n236));
  INV_X1    g035(.A(G113gat), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT1), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT73), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n244));
  INV_X1    g043(.A(new_n242), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n241), .A2(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT24), .B1(new_n213), .B2(new_n209), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(G183gat), .A3(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n229), .B2(new_n209), .ZN(new_n252));
  AND4_X1   g051(.A1(new_n251), .A2(new_n219), .A3(new_n221), .A4(new_n209), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT23), .B1(new_n203), .B2(new_n204), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G169gat), .B2(G176gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  OR2_X1    g059(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(KEYINPUT23), .A3(new_n203), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n247), .A2(new_n249), .B1(new_n213), .B2(new_n209), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n260), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n234), .A2(new_n246), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n227), .A2(KEYINPUT69), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n218), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n273), .A2(new_n208), .B1(new_n259), .B2(new_n266), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT74), .A3(new_n246), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n234), .A2(new_n267), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n244), .A2(new_n245), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n242), .B(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n277), .B1(new_n279), .B2(new_n240), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n270), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT64), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n202), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT75), .B(KEYINPUT33), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n282), .B2(new_n284), .ZN(new_n288));
  XOR2_X1   g087(.A(G15gat), .B(G43gat), .Z(new_n289));
  XNOR2_X1  g088(.A(G71gat), .B(G99gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n285), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  AOI221_X4 g092(.A(new_n202), .B1(new_n287), .B2(new_n291), .C1(new_n282), .C2(new_n284), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT77), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n270), .A2(new_n275), .A3(new_n281), .A4(new_n283), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT34), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n284), .A2(KEYINPUT34), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n270), .A2(new_n275), .A3(new_n281), .A4(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n297), .A2(KEYINPUT76), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT76), .B1(new_n297), .B2(new_n299), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n285), .ZN(new_n304));
  INV_X1    g103(.A(new_n288), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n291), .ZN(new_n306));
  INV_X1    g105(.A(new_n294), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n297), .A2(new_n299), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n297), .A2(KEYINPUT76), .A3(new_n299), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n308), .A2(new_n313), .A3(KEYINPUT77), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n303), .A2(new_n314), .A3(KEYINPUT36), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n293), .A2(new_n294), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n300), .B2(new_n301), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n311), .A2(KEYINPUT78), .A3(new_n312), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n308), .A2(new_n313), .A3(new_n317), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT36), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G1gat), .B(G29gat), .Z(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G57gat), .B(G85gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT5), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT83), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  INV_X1    g132(.A(G148gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(G155gat), .B2(G162gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G155gat), .B(G162gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT2), .B1(new_n330), .B2(new_n331), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(new_n335), .A3(new_n336), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(new_n341), .A3(new_n332), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n246), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n343), .A2(new_n346), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n280), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n329), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n246), .A2(KEYINPUT4), .A3(new_n347), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n280), .B1(new_n359), .B2(new_n347), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT84), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT84), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n362), .A3(new_n359), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n354), .B1(new_n365), .B2(new_n352), .ZN(new_n366));
  NOR4_X1   g165(.A1(new_n358), .A2(new_n364), .A3(new_n329), .A4(new_n353), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n328), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(KEYINPUT5), .A3(new_n352), .ZN(new_n369));
  INV_X1    g168(.A(new_n328), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n358), .A2(new_n364), .A3(new_n353), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n354), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n366), .A2(new_n367), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G197gat), .B(G204gat), .ZN(new_n378));
  AND2_X1   g177(.A1(G211gat), .A2(G218gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(KEYINPUT22), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G211gat), .B(G218gat), .Z(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(KEYINPUT79), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n380), .B(new_n381), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(KEYINPUT79), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n386));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n274), .B2(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n276), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n276), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT80), .B1(new_n393), .B2(new_n387), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n385), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n389), .B1(new_n276), .B2(new_n392), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n274), .A2(new_n387), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n396), .A2(new_n385), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n395), .A2(new_n399), .A3(KEYINPUT81), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT80), .B1(new_n396), .B2(new_n397), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n386), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n384), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n402), .B1(new_n411), .B2(new_n398), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT30), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n403), .B1(new_n395), .B2(new_n399), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n415), .A2(KEYINPUT82), .A3(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n377), .B(new_n408), .C1(new_n414), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G22gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n361), .B2(new_n363), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT86), .B1(new_n422), .B2(new_n385), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n362), .B1(new_n347), .B2(new_n359), .ZN(new_n424));
  AOI211_X1 g223(.A(KEYINPUT84), .B(KEYINPUT3), .C1(new_n343), .C2(new_n346), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n392), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n384), .ZN(new_n428));
  AND2_X1   g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n383), .A2(new_n392), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n359), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n431), .B2(new_n349), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n423), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n422), .A2(new_n385), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n392), .B(new_n382), .C1(new_n383), .C2(KEYINPUT79), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n347), .B1(new_n435), .B2(new_n359), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n429), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n433), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n433), .B2(new_n437), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n421), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n433), .A2(new_n437), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n438), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n433), .A2(new_n437), .A3(new_n439), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n420), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n418), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n323), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n374), .A2(new_n376), .A3(new_n412), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n403), .A2(KEYINPUT37), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n409), .A2(new_n410), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n398), .B1(new_n452), .B2(new_n385), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n404), .A2(new_n451), .B1(new_n453), .B2(KEYINPUT37), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT91), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n403), .B1(new_n453), .B2(KEYINPUT37), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n395), .A2(KEYINPUT37), .A3(new_n399), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n457), .B(KEYINPUT38), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n450), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n384), .B1(new_n391), .B2(new_n394), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(KEYINPUT88), .B(new_n384), .C1(new_n391), .C2(new_n394), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n388), .A2(new_n385), .A3(new_n390), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT89), .A3(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT38), .B1(new_n404), .B2(new_n451), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT89), .B1(new_n467), .B2(KEYINPUT37), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT90), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n468), .A4(new_n469), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n461), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n365), .B2(new_n352), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT87), .B(new_n353), .C1(new_n358), .C2(new_n364), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n351), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n352), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n328), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n482), .A2(KEYINPUT40), .A3(new_n328), .A4(new_n485), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n488), .A2(new_n372), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n416), .B1(new_n415), .B2(KEYINPUT82), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT30), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n491), .A2(new_n492), .B1(new_n406), .B2(new_n407), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n447), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n449), .B1(new_n476), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n303), .A2(new_n314), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n442), .A2(new_n446), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(new_n377), .A3(new_n493), .A4(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(new_n418), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n320), .A2(new_n321), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n499), .A2(KEYINPUT35), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G36gat), .ZN(new_n506));
  AND2_X1   g305(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G29gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n514));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(G1gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G1gat), .B2(new_n520), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G8gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n517), .A2(KEYINPUT93), .A3(new_n518), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT93), .B1(new_n517), .B2(new_n518), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(new_n524), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(KEYINPUT18), .A3(new_n529), .A4(new_n530), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n517), .B2(new_n524), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(new_n530), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n529), .B(KEYINPUT13), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G113gat), .B(G141gat), .Z(new_n541));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT12), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n531), .A2(new_n532), .B1(new_n538), .B2(new_n537), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n534), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n505), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G57gat), .B(G64gat), .Z(new_n554));
  XNOR2_X1  g353(.A(G71gat), .B(G78gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT9), .ZN(new_n556));
  INV_X1    g355(.A(G71gat), .ZN(new_n557));
  INV_X1    g356(.A(G78gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n554), .B2(new_n559), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OR3_X1    g363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G231gat), .ZN(new_n569));
  INV_X1    g368(.A(G233gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n566), .B(new_n567), .C1(new_n569), .C2(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G127gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n566), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n524), .B1(new_n576), .B2(KEYINPUT21), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G127gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n572), .A2(new_n579), .A3(new_n573), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n575), .B2(new_n580), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(new_n330), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OR3_X1    g387(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n588), .B1(new_n582), .B2(new_n583), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT7), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G99gat), .B(G106gat), .Z(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT96), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n597), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OAI221_X1 g405(.A(new_n606), .B1(new_n518), .B2(new_n517), .C1(new_n526), .C2(new_n527), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n517), .A2(new_n605), .B1(KEYINPUT41), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n607), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n607), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(KEYINPUT41), .ZN(new_n615));
  XNOR2_X1  g414(.A(G134gat), .B(G162gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OR3_X1    g417(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n613), .B2(new_n614), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT98), .B1(new_n591), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n598), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(new_n593), .A3(new_n597), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n562), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n566), .B2(new_n606), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT100), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  NOR2_X1   g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n628), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n566), .A2(new_n636), .A3(new_n606), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n627), .B2(new_n636), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n634), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n638), .B2(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n627), .A2(new_n636), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n576), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(KEYINPUT101), .A3(new_n628), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n629), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n633), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n639), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n621), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n589), .A2(new_n590), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n622), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n553), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n377), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n494), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT16), .B(G8gat), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT102), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT42), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  OAI211_X1 g463(.A(KEYINPUT102), .B(new_n664), .C1(new_n660), .C2(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(G8gat), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(G1325gat));
  INV_X1    g466(.A(G15gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n503), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n655), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT103), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n668), .A3(new_n323), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n655), .A2(new_n498), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n591), .A2(new_n649), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n650), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n553), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n377), .A2(G29gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n677), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n553), .A2(KEYINPUT45), .A3(new_n679), .A4(new_n681), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n418), .A2(KEYINPUT104), .A3(new_n447), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT36), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n503), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n303), .A2(new_n314), .A3(KEYINPUT36), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT104), .B1(new_n418), .B2(new_n447), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n476), .A2(new_n495), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n504), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n685), .B1(new_n694), .B2(new_n650), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n650), .A2(new_n685), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n496), .B2(new_n504), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(new_n552), .A3(new_n678), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(new_n657), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n683), .B(new_n684), .C1(new_n700), .C2(new_n510), .ZN(G1328gat));
  NOR2_X1   g500(.A1(new_n493), .A2(G36gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT46), .B1(new_n680), .B2(new_n703), .ZN(new_n704));
  OR3_X1    g503(.A1(new_n680), .A2(KEYINPUT46), .A3(new_n703), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n699), .A2(new_n494), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n704), .B(new_n705), .C1(new_n706), .C2(new_n506), .ZN(G1329gat));
  INV_X1    g506(.A(new_n698), .ZN(new_n708));
  INV_X1    g507(.A(new_n323), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n678), .A2(new_n552), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n680), .A2(G43gat), .A3(new_n669), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(G1330gat));
  NAND3_X1  g516(.A1(new_n708), .A2(new_n447), .A3(new_n710), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G50gat), .ZN(new_n719));
  OR3_X1    g518(.A1(new_n680), .A2(G50gat), .A3(new_n498), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1331gat));
  NAND4_X1  g523(.A1(new_n622), .A2(new_n552), .A3(new_n653), .A4(new_n648), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n727), .A2(new_n694), .A3(KEYINPUT106), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT106), .B1(new_n727), .B2(new_n694), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n657), .A2(KEYINPUT107), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n657), .A2(KEYINPUT107), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(G57gat), .Z(G1332gat));
  AND2_X1   g534(.A1(new_n728), .A2(new_n729), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n494), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND3_X1  g539(.A1(new_n736), .A2(G71gat), .A3(new_n709), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n503), .B(KEYINPUT108), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n557), .B1(new_n730), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n741), .B2(new_n743), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n498), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT110), .B(G78gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  NAND2_X1  g549(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n502), .A2(new_n503), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n476), .A2(new_n495), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n448), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n323), .A2(new_n756), .A3(new_n686), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n652), .A2(new_n551), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n621), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n693), .A2(new_n763), .A3(new_n756), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n650), .B1(new_n764), .B2(new_n753), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(KEYINPUT51), .A3(new_n759), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n595), .A3(new_n657), .A4(new_n648), .ZN(new_n768));
  INV_X1    g567(.A(new_n759), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n649), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n695), .A2(new_n697), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n377), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(G1336gat));
  NAND4_X1  g572(.A1(new_n767), .A2(new_n596), .A3(new_n494), .A4(new_n648), .ZN(new_n774));
  OAI21_X1  g573(.A(G92gat), .B1(new_n771), .B2(new_n493), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n778), .A3(KEYINPUT52), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n774), .B(new_n775), .C1(new_n777), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1337gat));
  NOR2_X1   g581(.A1(new_n669), .A2(G99gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n648), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G99gat), .B1(new_n771), .B2(new_n323), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1338gat));
  NOR2_X1   g585(.A1(new_n498), .A2(G106gat), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n765), .B2(new_n759), .ZN(new_n788));
  NOR4_X1   g587(.A1(new_n694), .A2(new_n761), .A3(new_n650), .A4(new_n769), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n648), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n695), .A2(new_n447), .A3(new_n697), .A4(new_n770), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n767), .A2(KEYINPUT113), .A3(new_n648), .A4(new_n787), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n792), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n790), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n790), .A2(new_n794), .A3(KEYINPUT114), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n800), .A2(new_n806), .ZN(G1339gat));
  INV_X1    g606(.A(new_n545), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n809), .A2(new_n810), .B1(new_n538), .B2(new_n537), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n550), .A3(new_n648), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n644), .B2(new_n628), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n638), .B2(new_n635), .ZN(new_n818));
  AND4_X1   g617(.A1(new_n817), .A2(new_n642), .A3(new_n635), .A4(new_n643), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n641), .A2(new_n645), .A3(new_n815), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT55), .A4(new_n633), .ZN(new_n822));
  INV_X1    g621(.A(new_n550), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n546), .B1(new_n549), .B2(new_n534), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n639), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n820), .A2(new_n633), .A3(new_n821), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n814), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n650), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n813), .A2(new_n550), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n822), .A2(new_n639), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n832), .A2(new_n621), .A3(new_n833), .A4(new_n828), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n652), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n622), .A2(new_n649), .A3(new_n653), .A4(new_n552), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n447), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n493), .A2(new_n657), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n669), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n237), .A3(new_n552), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n838), .A2(new_n733), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n497), .A2(new_n498), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n493), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n551), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n843), .B1(new_n237), .B2(new_n849), .ZN(G1340gat));
  OAI21_X1  g649(.A(G120gat), .B1(new_n842), .B2(new_n649), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n649), .A2(new_n235), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n847), .B2(new_n852), .ZN(G1341gat));
  AOI21_X1  g652(.A(G127gat), .B1(new_n848), .B2(new_n652), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n839), .A2(G127gat), .A3(new_n652), .A4(new_n841), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(G1342gat));
  OR3_X1    g658(.A1(new_n847), .A2(G134gat), .A3(new_n650), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n842), .B2(new_n650), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n709), .A2(new_n498), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n844), .A2(new_n493), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n551), .A2(new_n333), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT120), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n709), .A2(new_n840), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n838), .B2(new_n498), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n828), .A2(KEYINPUT119), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n826), .A2(new_n875), .A3(new_n827), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n874), .A2(new_n833), .A3(new_n551), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n621), .B1(new_n877), .B2(new_n814), .ZN(new_n878));
  INV_X1    g677(.A(new_n834), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n591), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n498), .B1(new_n880), .B2(new_n836), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n871), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n333), .B1(new_n883), .B2(new_n551), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT58), .B1(new_n869), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n825), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n826), .A2(new_n875), .A3(new_n827), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n875), .B1(new_n826), .B2(new_n827), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n886), .A2(new_n889), .B1(new_n648), .B2(new_n832), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n834), .B1(new_n890), .B2(new_n621), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n837), .B1(new_n891), .B2(new_n591), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(new_n498), .ZN(new_n894));
  INV_X1    g693(.A(new_n872), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n879), .B1(new_n650), .B2(new_n830), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n836), .B1(new_n896), .B2(new_n652), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n447), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n870), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n899), .B2(new_n552), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n883), .A2(new_n901), .A3(new_n551), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n900), .A2(G141gat), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n869), .A2(KEYINPUT58), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n885), .B1(new_n903), .B2(new_n904), .ZN(G1344gat));
  OAI211_X1 g704(.A(new_n447), .B(new_n895), .C1(new_n835), .C2(new_n837), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(new_n648), .A3(new_n870), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT59), .B1(new_n908), .B2(new_n334), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n648), .B(new_n870), .C1(new_n894), .C2(new_n898), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n334), .A2(KEYINPUT59), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n910), .A2(KEYINPUT122), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT122), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n866), .A2(new_n334), .A3(new_n648), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n899), .B2(new_n591), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n866), .A2(new_n330), .A3(new_n652), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  AOI21_X1  g718(.A(G162gat), .B1(new_n866), .B2(new_n621), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n650), .A2(new_n331), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n883), .B2(new_n921), .ZN(G1347gat));
  AOI21_X1  g721(.A(new_n493), .B1(new_n731), .B2(new_n732), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n742), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n839), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n203), .A3(new_n552), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n838), .A2(new_n657), .A3(new_n493), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n846), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n551), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n931), .B2(new_n203), .ZN(G1348gat));
  AOI21_X1  g731(.A(G176gat), .B1(new_n930), .B2(new_n648), .ZN(new_n933));
  INV_X1    g732(.A(new_n926), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n649), .B1(new_n261), .B2(new_n262), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G1349gat));
  OAI211_X1 g735(.A(new_n930), .B(new_n652), .C1(new_n216), .C2(new_n217), .ZN(new_n937));
  INV_X1    g736(.A(new_n229), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n938), .B1(new_n926), .B2(new_n591), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n209), .A3(new_n621), .ZN(new_n945));
  OAI21_X1  g744(.A(G190gat), .B1(new_n926), .B2(new_n650), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n950), .B1(new_n924), .B2(new_n709), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n323), .A2(KEYINPUT123), .A3(new_n923), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT124), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n893), .B1(new_n892), .B2(new_n498), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n906), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(KEYINPUT124), .A3(new_n952), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n955), .A2(G197gat), .A3(new_n551), .A4(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(G197gat), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n928), .A2(new_n865), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n552), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n957), .A2(new_n960), .ZN(G1352gat));
  NOR3_X1   g760(.A1(new_n959), .A2(G204gat), .A3(new_n649), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT62), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n955), .A2(new_n648), .A3(new_n956), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1353gat));
  OR3_X1    g765(.A1(new_n959), .A2(G211gat), .A3(new_n591), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n591), .B1(new_n951), .B2(new_n952), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n907), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  INV_X1    g771(.A(G218gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n973), .B1(new_n959), .B2(new_n650), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n955), .B2(new_n956), .ZN(new_n976));
  INV_X1    g775(.A(new_n953), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n907), .A2(new_n975), .A3(new_n956), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n621), .A2(G218gat), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT126), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n974), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g783(.A(KEYINPUT127), .B(new_n974), .C1(new_n976), .C2(new_n981), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1355gat));
endmodule


