

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U557 ( .A1(G651), .A2(n628), .ZN(n640) );
  OR2_X1 U558 ( .A1(n687), .A2(n982), .ZN(n690) );
  XNOR2_X1 U559 ( .A(n582), .B(KEYINPUT15), .ZN(n988) );
  AND2_X2 U560 ( .A1(n525), .A2(G2104), .ZN(n877) );
  NAND2_X1 U561 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U562 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U563 ( .A1(n690), .A2(n689), .ZN(n696) );
  INV_X1 U564 ( .A(KEYINPUT32), .ZN(n733) );
  XNOR2_X1 U565 ( .A(n734), .B(n733), .ZN(n742) );
  INV_X1 U566 ( .A(n767), .ZN(n750) );
  NAND2_X1 U567 ( .A1(n772), .A2(n774), .ZN(n725) );
  XNOR2_X1 U568 ( .A(n686), .B(KEYINPUT89), .ZN(n772) );
  NOR2_X1 U569 ( .A1(n777), .A2(n776), .ZN(n808) );
  NOR2_X1 U570 ( .A1(n628), .A2(n535), .ZN(n638) );
  NOR2_X1 U571 ( .A1(n530), .A2(n529), .ZN(G160) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U573 ( .A1(G113), .A2(n879), .ZN(n521) );
  XNOR2_X1 U574 ( .A(n521), .B(KEYINPUT64), .ZN(n524) );
  INV_X1 U575 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U576 ( .A1(G101), .A2(n877), .ZN(n522) );
  XOR2_X1 U577 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U578 ( .A1(n524), .A2(n523), .ZN(n530) );
  NOR2_X1 U579 ( .A1(G2104), .A2(n525), .ZN(n880) );
  NAND2_X1 U580 ( .A1(G125), .A2(n880), .ZN(n528) );
  NOR2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U582 ( .A(KEYINPUT17), .B(n526), .Z(n885) );
  NAND2_X1 U583 ( .A1(G137), .A2(n885), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U585 ( .A(G651), .ZN(n535) );
  NOR2_X1 U586 ( .A1(G543), .A2(n535), .ZN(n532) );
  XNOR2_X1 U587 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n531) );
  XNOR2_X1 U588 ( .A(n532), .B(n531), .ZN(n644) );
  NAND2_X1 U589 ( .A1(G60), .A2(n644), .ZN(n534) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U591 ( .A1(G85), .A2(n641), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n539) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NAND2_X1 U594 ( .A1(G72), .A2(n638), .ZN(n537) );
  NAND2_X1 U595 ( .A1(G47), .A2(n640), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n538) );
  OR2_X1 U597 ( .A1(n539), .A2(n538), .ZN(G290) );
  NAND2_X1 U598 ( .A1(n638), .A2(G77), .ZN(n540) );
  XOR2_X1 U599 ( .A(KEYINPUT67), .B(n540), .Z(n542) );
  NAND2_X1 U600 ( .A1(n641), .A2(G90), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n543), .B(KEYINPUT9), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G52), .A2(n640), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n644), .A2(G64), .ZN(n546) );
  XOR2_X1 U606 ( .A(KEYINPUT66), .B(n546), .Z(n547) );
  NOR2_X1 U607 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U609 ( .A(G120), .ZN(G236) );
  INV_X1 U610 ( .A(G69), .ZN(G235) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n638), .A2(G76), .ZN(n549) );
  XNOR2_X1 U616 ( .A(KEYINPUT74), .B(n549), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n641), .A2(G89), .ZN(n550) );
  XNOR2_X1 U618 ( .A(KEYINPUT4), .B(n550), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT5), .ZN(n559) );
  XNOR2_X1 U621 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G51), .A2(n640), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G63), .A2(n644), .ZN(n554) );
  NAND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G168) );
  XOR2_X1 U628 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U631 ( .A(G567), .ZN(n674) );
  NOR2_X1 U632 ( .A1(n674), .A2(G223), .ZN(n563) );
  XNOR2_X1 U633 ( .A(n563), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U634 ( .A1(n641), .A2(G81), .ZN(n564) );
  XNOR2_X1 U635 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U636 ( .A1(G68), .A2(n638), .ZN(n565) );
  NAND2_X1 U637 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n567), .Z(n570) );
  NAND2_X1 U639 ( .A1(n644), .A2(G56), .ZN(n568) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n568), .Z(n569) );
  NOR2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n640), .A2(G43), .ZN(n571) );
  NAND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n982) );
  INV_X1 U644 ( .A(G860), .ZN(n595) );
  OR2_X1 U645 ( .A1(n982), .A2(n595), .ZN(G153) );
  XOR2_X1 U646 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n573) );
  XOR2_X1 U648 ( .A(KEYINPUT71), .B(n573), .Z(n584) );
  NAND2_X1 U649 ( .A1(G79), .A2(n638), .ZN(n575) );
  NAND2_X1 U650 ( .A1(G54), .A2(n640), .ZN(n574) );
  NAND2_X1 U651 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n576), .B(KEYINPUT72), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n641), .A2(G92), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n644), .A2(G66), .ZN(n577) );
  NAND2_X1 U655 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U656 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U657 ( .A(n581), .B(KEYINPUT73), .ZN(n582) );
  INV_X1 U658 ( .A(n988), .ZN(n598) );
  INV_X1 U659 ( .A(G868), .ZN(n660) );
  NAND2_X1 U660 ( .A1(n598), .A2(n660), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G91), .A2(n641), .ZN(n585) );
  XNOR2_X1 U663 ( .A(n585), .B(KEYINPUT68), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n638), .A2(G78), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U666 ( .A1(G65), .A2(n644), .ZN(n588) );
  XNOR2_X1 U667 ( .A(KEYINPUT69), .B(n588), .ZN(n589) );
  NOR2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n640), .A2(G53), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(G299) );
  NAND2_X1 U671 ( .A1(G868), .A2(G286), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G299), .A2(n660), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n596), .A2(n988), .ZN(n597) );
  XNOR2_X1 U676 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(n598), .A2(n660), .ZN(n599) );
  XNOR2_X1 U678 ( .A(n599), .B(KEYINPUT77), .ZN(n600) );
  NOR2_X1 U679 ( .A1(G559), .A2(n600), .ZN(n602) );
  NOR2_X1 U680 ( .A1(G868), .A2(n982), .ZN(n601) );
  NOR2_X1 U681 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U682 ( .A1(n879), .A2(G111), .ZN(n603) );
  XOR2_X1 U683 ( .A(KEYINPUT79), .B(n603), .Z(n605) );
  NAND2_X1 U684 ( .A1(n877), .A2(G99), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U686 ( .A(KEYINPUT80), .B(n606), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G123), .A2(n880), .ZN(n607) );
  XNOR2_X1 U688 ( .A(n607), .B(KEYINPUT78), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G135), .A2(n885), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n947) );
  XNOR2_X1 U693 ( .A(n947), .B(G2096), .ZN(n614) );
  INV_X1 U694 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U696 ( .A1(n988), .A2(G559), .ZN(n656) );
  XNOR2_X1 U697 ( .A(n982), .B(n656), .ZN(n615) );
  NOR2_X1 U698 ( .A1(n615), .A2(G860), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G80), .A2(n638), .ZN(n617) );
  NAND2_X1 U700 ( .A1(G93), .A2(n641), .ZN(n616) );
  NAND2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G55), .A2(n640), .ZN(n619) );
  NAND2_X1 U703 ( .A1(G67), .A2(n644), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U705 ( .A(KEYINPUT81), .B(n620), .Z(n621) );
  OR2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n659) );
  XOR2_X1 U707 ( .A(n623), .B(n659), .Z(G145) );
  NAND2_X1 U708 ( .A1(G49), .A2(n640), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U711 ( .A1(n644), .A2(n626), .ZN(n627) );
  XNOR2_X1 U712 ( .A(n627), .B(KEYINPUT82), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G87), .A2(n628), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G62), .A2(n644), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G88), .A2(n641), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n638), .A2(G75), .ZN(n633) );
  XOR2_X1 U719 ( .A(KEYINPUT84), .B(n633), .Z(n634) );
  NOR2_X1 U720 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n640), .A2(G50), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(G303) );
  INV_X1 U723 ( .A(G303), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G73), .A2(n638), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n639), .B(KEYINPUT2), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G48), .A2(n640), .ZN(n643) );
  NAND2_X1 U727 ( .A1(G86), .A2(n641), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U729 ( .A1(G61), .A2(n644), .ZN(n645) );
  XNOR2_X1 U730 ( .A(KEYINPUT83), .B(n645), .ZN(n646) );
  NOR2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U732 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(G288), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n650), .B(G290), .ZN(n651) );
  XNOR2_X1 U735 ( .A(n651), .B(n659), .ZN(n653) );
  INV_X1 U736 ( .A(G299), .ZN(n977) );
  XNOR2_X1 U737 ( .A(n977), .B(G166), .ZN(n652) );
  XNOR2_X1 U738 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U739 ( .A(n654), .B(n982), .ZN(n655) );
  XNOR2_X1 U740 ( .A(n655), .B(G305), .ZN(n897) );
  XNOR2_X1 U741 ( .A(KEYINPUT85), .B(n656), .ZN(n657) );
  XNOR2_X1 U742 ( .A(n897), .B(n657), .ZN(n658) );
  NAND2_X1 U743 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n664), .ZN(n666) );
  XNOR2_X1 U749 ( .A(KEYINPUT86), .B(KEYINPUT21), .ZN(n665) );
  XNOR2_X1 U750 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U751 ( .A1(G2072), .A2(n667), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U755 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U756 ( .A1(G96), .A2(n670), .ZN(n832) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n832), .ZN(n671) );
  XNOR2_X1 U758 ( .A(n671), .B(KEYINPUT87), .ZN(n676) );
  NOR2_X1 U759 ( .A1(G235), .A2(G236), .ZN(n672) );
  NAND2_X1 U760 ( .A1(G108), .A2(n672), .ZN(n673) );
  NOR2_X1 U761 ( .A1(G237), .A2(n673), .ZN(n834) );
  NOR2_X1 U762 ( .A1(n674), .A2(n834), .ZN(n675) );
  NOR2_X1 U763 ( .A1(n676), .A2(n675), .ZN(G319) );
  INV_X1 U764 ( .A(G319), .ZN(n678) );
  NAND2_X1 U765 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U766 ( .A1(n678), .A2(n677), .ZN(n831) );
  NAND2_X1 U767 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U768 ( .A1(n879), .A2(G114), .ZN(n679) );
  XNOR2_X1 U769 ( .A(n679), .B(KEYINPUT88), .ZN(n681) );
  NAND2_X1 U770 ( .A1(G102), .A2(n877), .ZN(n680) );
  NAND2_X1 U771 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U772 ( .A1(G126), .A2(n880), .ZN(n683) );
  NAND2_X1 U773 ( .A1(G138), .A2(n885), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U775 ( .A1(n685), .A2(n684), .ZN(G164) );
  NOR2_X1 U776 ( .A1(G1971), .A2(G303), .ZN(n745) );
  XNOR2_X1 U777 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n709) );
  NAND2_X1 U778 ( .A1(G40), .A2(G160), .ZN(n686) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n774) );
  AND2_X1 U780 ( .A1(n725), .A2(G1341), .ZN(n687) );
  INV_X1 U781 ( .A(G1996), .ZN(n924) );
  NOR2_X1 U782 ( .A1(n725), .A2(n924), .ZN(n688) );
  XNOR2_X1 U783 ( .A(n688), .B(KEYINPUT26), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n696), .A2(n988), .ZN(n694) );
  NOR2_X1 U785 ( .A1(G2067), .A2(n725), .ZN(n692) );
  INV_X1 U786 ( .A(n725), .ZN(n710) );
  NOR2_X1 U787 ( .A1(n710), .A2(G1348), .ZN(n691) );
  NOR2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U790 ( .A(n695), .B(KEYINPUT96), .ZN(n698) );
  OR2_X1 U791 ( .A1(n696), .A2(n988), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n710), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U794 ( .A(n699), .B(KEYINPUT27), .ZN(n701) );
  INV_X1 U795 ( .A(G1956), .ZN(n1003) );
  NOR2_X1 U796 ( .A1(n1003), .A2(n710), .ZN(n700) );
  NOR2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n977), .A2(n704), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U800 ( .A1(n977), .A2(n704), .ZN(n705) );
  XOR2_X1 U801 ( .A(n705), .B(KEYINPUT28), .Z(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U803 ( .A(n709), .B(n708), .ZN(n714) );
  INV_X1 U804 ( .A(G1961), .ZN(n1001) );
  NAND2_X1 U805 ( .A1(n725), .A2(n1001), .ZN(n712) );
  XNOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .ZN(n928) );
  NAND2_X1 U807 ( .A1(n710), .A2(n928), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n718), .A2(G171), .ZN(n713) );
  NAND2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n723) );
  NAND2_X1 U811 ( .A1(G8), .A2(n725), .ZN(n767) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n767), .ZN(n738) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n725), .ZN(n735) );
  NOR2_X1 U814 ( .A1(n738), .A2(n735), .ZN(n715) );
  NAND2_X1 U815 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U817 ( .A1(G168), .A2(n717), .ZN(n720) );
  NOR2_X1 U818 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U819 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n721), .Z(n722) );
  NAND2_X1 U821 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U822 ( .A(KEYINPUT98), .B(n724), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n736), .A2(G286), .ZN(n732) );
  INV_X1 U824 ( .A(G8), .ZN(n730) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n767), .ZN(n727) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n725), .ZN(n726) );
  NOR2_X1 U827 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U828 ( .A1(n728), .A2(G303), .ZN(n729) );
  OR2_X1 U829 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U830 ( .A1(G8), .A2(n735), .ZN(n740) );
  INV_X1 U831 ( .A(n736), .ZN(n737) );
  NOR2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n763) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n743) );
  XNOR2_X1 U836 ( .A(KEYINPUT99), .B(n743), .ZN(n989) );
  NAND2_X1 U837 ( .A1(n763), .A2(n989), .ZN(n744) );
  NOR2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n753) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n986) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n755) );
  OR2_X1 U841 ( .A1(n767), .A2(n989), .ZN(n746) );
  NOR2_X1 U842 ( .A1(n755), .A2(n746), .ZN(n747) );
  XOR2_X1 U843 ( .A(n747), .B(KEYINPUT100), .Z(n754) );
  AND2_X1 U844 ( .A1(n986), .A2(n754), .ZN(n749) );
  XNOR2_X1 U845 ( .A(G1981), .B(G305), .ZN(n975) );
  INV_X1 U846 ( .A(n975), .ZN(n748) );
  AND2_X1 U847 ( .A1(n749), .A2(n748), .ZN(n751) );
  OR2_X1 U848 ( .A1(n753), .A2(n752), .ZN(n759) );
  INV_X1 U849 ( .A(n754), .ZN(n756) );
  OR2_X1 U850 ( .A1(n756), .A2(n755), .ZN(n757) );
  OR2_X1 U851 ( .A1(n975), .A2(n757), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U853 ( .A(KEYINPUT101), .B(n760), .ZN(n771) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n761) );
  NAND2_X1 U855 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  AND2_X1 U857 ( .A1(n767), .A2(n764), .ZN(n769) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XOR2_X1 U859 ( .A(n765), .B(KEYINPUT24), .Z(n766) );
  NOR2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n770) );
  AND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n777) );
  INV_X1 U863 ( .A(n772), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n821) );
  XNOR2_X1 U865 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U866 ( .A1(n821), .A2(n979), .ZN(n775) );
  XOR2_X1 U867 ( .A(KEYINPUT90), .B(n775), .Z(n776) );
  XOR2_X1 U868 ( .A(n821), .B(KEYINPUT95), .Z(n797) );
  NAND2_X1 U869 ( .A1(n877), .A2(G105), .ZN(n779) );
  XNOR2_X1 U870 ( .A(KEYINPUT94), .B(KEYINPUT38), .ZN(n778) );
  XNOR2_X1 U871 ( .A(n779), .B(n778), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G117), .A2(n879), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G141), .A2(n885), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G129), .A2(n880), .ZN(n782) );
  XNOR2_X1 U876 ( .A(KEYINPUT93), .B(n782), .ZN(n783) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n891) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n891), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G95), .A2(n877), .ZN(n787) );
  XNOR2_X1 U881 ( .A(n787), .B(KEYINPUT92), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G119), .A2(n880), .ZN(n789) );
  NAND2_X1 U883 ( .A1(G131), .A2(n885), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U885 ( .A1(G107), .A2(n879), .ZN(n790) );
  XNOR2_X1 U886 ( .A(KEYINPUT91), .B(n790), .ZN(n791) );
  NOR2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n890) );
  NAND2_X1 U889 ( .A1(G1991), .A2(n890), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n952) );
  NAND2_X1 U891 ( .A1(n797), .A2(n952), .ZN(n810) );
  NAND2_X1 U892 ( .A1(G104), .A2(n877), .ZN(n799) );
  NAND2_X1 U893 ( .A1(G140), .A2(n885), .ZN(n798) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U895 ( .A(KEYINPUT34), .B(n800), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G116), .A2(n879), .ZN(n802) );
  NAND2_X1 U897 ( .A1(G128), .A2(n880), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U899 ( .A(KEYINPUT35), .B(n803), .Z(n804) );
  NOR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U901 ( .A(KEYINPUT36), .B(n806), .Z(n874) );
  XOR2_X1 U902 ( .A(G2067), .B(KEYINPUT37), .Z(n820) );
  AND2_X1 U903 ( .A1(n874), .A2(n820), .ZN(n948) );
  NAND2_X1 U904 ( .A1(n948), .A2(n821), .ZN(n809) );
  AND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n807) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n825) );
  INV_X1 U907 ( .A(n809), .ZN(n819) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n891), .ZN(n958) );
  INV_X1 U909 ( .A(n810), .ZN(n813) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n890), .ZN(n946) );
  NOR2_X1 U912 ( .A1(n811), .A2(n946), .ZN(n812) );
  NOR2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U914 ( .A1(n958), .A2(n814), .ZN(n816) );
  XNOR2_X1 U915 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n815) );
  XNOR2_X1 U916 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U917 ( .A1(n821), .A2(n817), .ZN(n818) );
  OR2_X1 U918 ( .A1(n819), .A2(n818), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n874), .A2(n820), .ZN(n955) );
  NAND2_X1 U920 ( .A1(n955), .A2(n821), .ZN(n822) );
  AND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U924 ( .A(G223), .ZN(n827) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n827), .ZN(G217) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n828) );
  XOR2_X1 U927 ( .A(KEYINPUT104), .B(n828), .Z(n829) );
  NAND2_X1 U928 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U930 ( .A1(n831), .A2(n830), .ZN(G188) );
  XNOR2_X1 U931 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(n832), .ZN(n833) );
  NAND2_X1 U935 ( .A1(n834), .A2(n833), .ZN(G261) );
  INV_X1 U936 ( .A(G261), .ZN(G325) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n836) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n838) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U942 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U943 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT106), .B(G1991), .Z(n844) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1996), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U949 ( .A(n845), .B(KEYINPUT41), .Z(n847) );
  XNOR2_X1 U950 ( .A(G1971), .B(G1976), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U952 ( .A(G1986), .B(G1981), .Z(n849) );
  XNOR2_X1 U953 ( .A(G1956), .B(G1961), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U955 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U956 ( .A(KEYINPUT105), .B(G2474), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G112), .A2(n879), .ZN(n855) );
  NAND2_X1 U959 ( .A1(G100), .A2(n877), .ZN(n854) );
  NAND2_X1 U960 ( .A1(n855), .A2(n854), .ZN(n861) );
  NAND2_X1 U961 ( .A1(n880), .A2(G124), .ZN(n856) );
  XNOR2_X1 U962 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U963 ( .A1(G136), .A2(n885), .ZN(n857) );
  NAND2_X1 U964 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U965 ( .A(KEYINPUT107), .B(n859), .Z(n860) );
  NOR2_X1 U966 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n872) );
  NAND2_X1 U968 ( .A1(G118), .A2(n879), .ZN(n863) );
  NAND2_X1 U969 ( .A1(G130), .A2(n880), .ZN(n862) );
  NAND2_X1 U970 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G106), .A2(n877), .ZN(n865) );
  NAND2_X1 U972 ( .A1(G142), .A2(n885), .ZN(n864) );
  NAND2_X1 U973 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n866), .Z(n867) );
  XNOR2_X1 U975 ( .A(KEYINPUT108), .B(n867), .ZN(n868) );
  NOR2_X1 U976 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U977 ( .A(G164), .B(n870), .ZN(n871) );
  XNOR2_X1 U978 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U979 ( .A(n873), .B(n947), .Z(n876) );
  XNOR2_X1 U980 ( .A(n874), .B(G162), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n895) );
  NAND2_X1 U982 ( .A1(n877), .A2(G103), .ZN(n878) );
  XNOR2_X1 U983 ( .A(KEYINPUT109), .B(n878), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G115), .A2(n879), .ZN(n882) );
  NAND2_X1 U985 ( .A1(G127), .A2(n880), .ZN(n881) );
  NAND2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n883), .B(KEYINPUT47), .ZN(n884) );
  XNOR2_X1 U988 ( .A(n884), .B(KEYINPUT110), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n885), .A2(G139), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n888) );
  NOR2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n962) );
  XNOR2_X1 U992 ( .A(n962), .B(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(G160), .B(n893), .Z(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U996 ( .A1(G37), .A2(n896), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n899) );
  XNOR2_X1 U998 ( .A(n988), .B(n897), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(G286), .B(G171), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U1003 ( .A(KEYINPUT103), .B(G2427), .Z(n904) );
  XNOR2_X1 U1004 ( .A(G2435), .B(G2438), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n904), .B(n903), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G2443), .B(G2430), .Z(n906) );
  XNOR2_X1 U1007 ( .A(G2454), .B(G2446), .ZN(n905) );
  XNOR2_X1 U1008 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1009 ( .A(n907), .B(G2451), .Z(n909) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1011 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(n912), .A2(G14), .ZN(n918) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1022 ( .A(G2090), .B(G35), .Z(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT54), .B(G34), .ZN(n919) );
  XNOR2_X1 U1024 ( .A(n919), .B(KEYINPUT119), .ZN(n920) );
  XNOR2_X1 U1025 ( .A(G2084), .B(n920), .ZN(n921) );
  NAND2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n938) );
  XOR2_X1 U1027 ( .A(G1991), .B(G25), .Z(n923) );
  NAND2_X1 U1028 ( .A1(n923), .A2(G28), .ZN(n927) );
  XOR2_X1 U1029 ( .A(KEYINPUT118), .B(n924), .Z(n925) );
  XNOR2_X1 U1030 ( .A(G32), .B(n925), .ZN(n926) );
  NOR2_X1 U1031 ( .A1(n927), .A2(n926), .ZN(n935) );
  XOR2_X1 U1032 ( .A(n928), .B(G27), .Z(n933) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1034 ( .A(G2072), .B(G33), .ZN(n929) );
  NOR2_X1 U1035 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1036 ( .A(KEYINPUT117), .B(n931), .ZN(n932) );
  NOR2_X1 U1037 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1039 ( .A(n936), .B(KEYINPUT53), .Z(n937) );
  NOR2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1041 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n969) );
  XOR2_X1 U1042 ( .A(n939), .B(n969), .Z(n940) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n940), .ZN(n942) );
  INV_X1 U1044 ( .A(G29), .ZN(n941) );
  NAND2_X1 U1045 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1046 ( .A1(n943), .A2(G11), .ZN(n944) );
  XNOR2_X1 U1047 ( .A(n944), .B(KEYINPUT121), .ZN(n973) );
  XOR2_X1 U1048 ( .A(G2084), .B(G160), .Z(n945) );
  NOR2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1053 ( .A(KEYINPUT114), .B(n953), .Z(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G162), .ZN(n956) );
  XNOR2_X1 U1056 ( .A(n956), .B(KEYINPUT115), .ZN(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1058 ( .A(KEYINPUT51), .B(n959), .Z(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n967) );
  XOR2_X1 U1060 ( .A(G2072), .B(n962), .Z(n964) );
  XOR2_X1 U1061 ( .A(G164), .B(G2078), .Z(n963) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1063 ( .A(KEYINPUT50), .B(n965), .Z(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT52), .B(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n971), .A2(G29), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n1030) );
  XNOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XOR2_X1 U1070 ( .A(G1966), .B(G168), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1072 ( .A(KEYINPUT57), .B(n976), .Z(n998) );
  XNOR2_X1 U1073 ( .A(n977), .B(G1956), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G303), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n985) );
  XOR2_X1 U1077 ( .A(G1341), .B(n982), .Z(n983) );
  XNOR2_X1 U1078 ( .A(KEYINPUT123), .B(n983), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(n988), .B(G1348), .ZN(n993) );
  XOR2_X1 U1082 ( .A(G171), .B(G1961), .Z(n991) );
  XOR2_X1 U1083 ( .A(n989), .B(KEYINPUT122), .Z(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT124), .B(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1027) );
  INV_X1 U1090 ( .A(G16), .ZN(n1025) );
  XNOR2_X1 U1091 ( .A(G5), .B(n1001), .ZN(n1015) );
  XNOR2_X1 U1092 ( .A(KEYINPUT59), .B(G1348), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(G4), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(G1341), .B(G19), .Z(n1005) );
  XNOR2_X1 U1095 ( .A(n1003), .B(G20), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G6), .B(G1981), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n1010) );
  XNOR2_X1 U1101 ( .A(n1011), .B(n1010), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G23), .B(G1976), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(G1986), .B(G24), .Z(n1018) );
  NAND2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(n1028), .B(KEYINPUT126), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(n1031), .B(KEYINPUT127), .Z(n1032) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1032), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

