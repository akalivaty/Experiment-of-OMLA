//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT22), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n197));
  INV_X1    g011(.A(G110), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n192), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT24), .B(G110), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(new_n195), .A3(new_n198), .A4(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G140), .ZN(new_n211));
  XNOR2_X1  g025(.A(G125), .B(G140), .ZN(new_n212));
  MUX2_X1   g026(.A(new_n211), .B(new_n212), .S(KEYINPUT16), .Z(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n212), .B(KEYINPUT77), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n214), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n201), .A2(KEYINPUT76), .A3(new_n204), .A4(new_n206), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n209), .A2(new_n216), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n196), .A2(new_n200), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G110), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n213), .A2(new_n214), .ZN(new_n223));
  OAI221_X1 g037(.A(new_n222), .B1(new_n202), .B2(new_n203), .C1(new_n223), .C2(new_n215), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n190), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n220), .A2(new_n224), .A3(new_n190), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(G234), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G902), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT78), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n220), .A2(new_n224), .A3(new_n190), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT78), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n235), .B2(new_n229), .ZN(new_n240));
  NOR4_X1   g054(.A1(new_n234), .A2(new_n225), .A3(KEYINPUT25), .A4(G902), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n238), .B1(new_n242), .B2(new_n230), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT11), .B1(new_n246), .B2(G137), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n249), .B2(G134), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n246), .A2(KEYINPUT64), .A3(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n251), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n251), .B2(new_n255), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n245), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n251), .A2(new_n255), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G131), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n251), .A2(new_n255), .A3(new_n256), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(KEYINPUT67), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n214), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n267), .B2(new_n269), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n259), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT1), .B1(new_n265), .B2(G146), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n264), .A2(KEYINPUT65), .A3(KEYINPUT1), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(G128), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n267), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n279));
  AND4_X1   g093(.A1(new_n279), .A2(new_n264), .A3(new_n266), .A4(G128), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n283));
  XOR2_X1   g097(.A(G134), .B(G137), .Z(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G131), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n262), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  OR2_X1    g101(.A1(KEYINPUT2), .A2(G113), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n199), .A2(G116), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G119), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT2), .A2(G113), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n288), .A2(new_n289), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n292), .ZN(new_n296));
  NOR2_X1   g110(.A1(KEYINPUT2), .A2(G113), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G116), .B(G119), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT66), .ZN(new_n300));
  INV_X1    g114(.A(new_n299), .ZN(new_n301));
  INV_X1    g115(.A(new_n298), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n295), .A2(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n280), .B1(new_n277), .B2(new_n267), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n262), .A2(new_n285), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT68), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n272), .A2(new_n287), .A3(new_n303), .A4(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G237), .ZN(new_n311));
  AOI21_X1  g125(.A(G953), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G210), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n312), .B2(G210), .ZN(new_n316));
  OR3_X1    g130(.A1(new_n315), .A2(KEYINPUT26), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT26), .B1(new_n315), .B2(new_n316), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n317), .A2(G101), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(G101), .B1(new_n317), .B2(new_n318), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n264), .A2(new_n266), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n191), .B1(new_n273), .B2(new_n274), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(new_n276), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n262), .B(new_n285), .C1(new_n324), .C2(new_n280), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n271), .B1(new_n257), .B2(new_n258), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n272), .A2(new_n287), .A3(new_n306), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(KEYINPUT30), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n307), .B(new_n321), .C1(new_n330), .C2(new_n303), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT31), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n333));
  INV_X1    g147(.A(new_n321), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n272), .A2(KEYINPUT73), .A3(new_n325), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT73), .B1(new_n272), .B2(new_n325), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT28), .B1(new_n338), .B2(new_n303), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n325), .A2(new_n326), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n302), .A2(new_n301), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n293), .A2(new_n294), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT66), .B1(new_n298), .B2(new_n299), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n342), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  AOI211_X1 g162(.A(KEYINPUT72), .B(new_n303), .C1(new_n325), .C2(new_n326), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n341), .B1(new_n350), .B2(new_n307), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n334), .B1(new_n339), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n307), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n329), .A2(KEYINPUT30), .ZN(new_n354));
  INV_X1    g168(.A(new_n328), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n353), .B1(new_n356), .B2(new_n347), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT31), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n321), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n331), .A2(new_n360), .A3(KEYINPUT31), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n333), .A2(new_n352), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(G472), .A2(G902), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n362), .A2(KEYINPUT32), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT32), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT74), .B1(new_n357), .B2(new_n321), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n368));
  INV_X1    g182(.A(new_n348), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n343), .A2(new_n342), .A3(new_n347), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n307), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n340), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n272), .A2(new_n325), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n303), .A3(new_n335), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT28), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(new_n378), .A3(new_n321), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n307), .B1(new_n330), .B2(new_n303), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n334), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n367), .A2(new_n368), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n329), .A2(new_n347), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT28), .B1(new_n384), .B2(new_n353), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n385), .A2(new_n378), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n334), .A2(new_n368), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G472), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n244), .B1(new_n366), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G469), .ZN(new_n392));
  XNOR2_X1  g206(.A(G110), .B(G140), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n187), .A2(G227), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n393), .B(new_n394), .Z(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(new_n396), .B2(G107), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G104), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  INV_X1    g217(.A(G101), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n397), .A2(new_n400), .A3(new_n404), .A4(new_n401), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n407), .A3(G101), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n271), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n273), .A2(G128), .B1(new_n264), .B2(new_n266), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n280), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n399), .A2(G104), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n396), .A2(G107), .ZN(new_n414));
  OAI21_X1  g228(.A(G101), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n405), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n410), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n409), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n410), .B1(new_n278), .B2(new_n281), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n405), .A2(new_n415), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n420), .B(KEYINPUT10), .C1(new_n324), .C2(new_n280), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n259), .A2(new_n263), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT83), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n409), .A2(new_n417), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT79), .B1(new_n419), .B2(new_n420), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n422), .A2(new_n423), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n259), .A2(new_n263), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n421), .A2(new_n424), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n259), .B2(new_n263), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n259), .A2(new_n263), .A3(new_n437), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n436), .B(new_n428), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n395), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n304), .A2(new_n416), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n420), .B1(new_n280), .B2(new_n411), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n442), .B1(new_n445), .B2(new_n426), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n261), .A2(new_n262), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n443), .B2(new_n444), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(new_n440), .A3(new_n395), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n392), .B(new_n229), .C1(new_n441), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n439), .A2(new_n438), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n443), .A2(new_n444), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT12), .B1(new_n433), .B2(new_n456), .ZN(new_n457));
  OAI22_X1  g271(.A1(new_n431), .A2(new_n455), .B1(new_n457), .B2(new_n450), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT82), .ZN(new_n459));
  INV_X1    g273(.A(new_n395), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n452), .A2(new_n440), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n435), .A2(new_n395), .A3(new_n440), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(G469), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(G469), .A2(G902), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n454), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G221), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT9), .B(G234), .Z(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(new_n229), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G475), .A2(G902), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT20), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(new_n396), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n212), .A2(new_n214), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n217), .B2(new_n214), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n310), .A2(G237), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n483));
  OAI211_X1 g297(.A(G214), .B(new_n187), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n265), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n312), .A2(G143), .A3(G214), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(KEYINPUT18), .A2(G131), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n484), .A2(new_n265), .ZN(new_n490));
  AOI21_X1  g304(.A(G143), .B1(new_n312), .B2(G214), .ZN(new_n491));
  OAI211_X1 g305(.A(KEYINPUT18), .B(G131), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT92), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n256), .B1(new_n485), .B2(new_n486), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT92), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT18), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n481), .B(new_n489), .C1(new_n493), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n487), .A2(G131), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n485), .A2(new_n256), .A3(new_n486), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT19), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n212), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n217), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n214), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n504), .A3(new_n216), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n479), .B1(new_n497), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n481), .ZN(new_n508));
  INV_X1    g322(.A(new_n489), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n492), .A2(KEYINPUT92), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n495), .B1(new_n494), .B2(KEYINPUT18), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n223), .A2(new_n215), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n494), .A2(KEYINPUT17), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n514), .C1(new_n500), .C2(KEYINPUT17), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n478), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n476), .B1(new_n507), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n512), .A2(new_n478), .A3(new_n515), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n478), .B1(new_n512), .B2(new_n505), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT93), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n507), .A2(new_n522), .A3(new_n516), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n474), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT13), .B1(new_n191), .B2(G143), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n246), .ZN(new_n530));
  XNOR2_X1  g344(.A(G128), .B(G143), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G122), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G116), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(G122), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(G116), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n536), .A2(new_n399), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n399), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n536), .B1(KEYINPUT14), .B2(new_n399), .ZN(new_n540));
  INV_X1    g354(.A(new_n538), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT14), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n535), .B2(G116), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n531), .B(G134), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n469), .A2(G217), .A3(new_n187), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n547), .B(KEYINPUT95), .Z(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n549), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n229), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n528), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  INV_X1    g370(.A(new_n552), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(new_n550), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT96), .A3(new_n229), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n555), .B1(new_n560), .B2(new_n528), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n478), .B1(new_n512), .B2(new_n515), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n519), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n229), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G475), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n526), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n472), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G952), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n187), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(G234), .B2(G237), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT21), .B(G898), .ZN(new_n573));
  AOI211_X1 g387(.A(new_n229), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(G214), .B1(G237), .B2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n347), .A2(new_n408), .A3(new_n406), .ZN(new_n578));
  XOR2_X1   g392(.A(G110), .B(G122), .Z(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n295), .A2(new_n300), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n289), .A2(new_n291), .A3(KEYINPUT5), .ZN(new_n582));
  OR3_X1    g396(.A1(new_n290), .A2(KEYINPUT5), .A3(G119), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(G113), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT84), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT84), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n582), .A2(new_n583), .A3(new_n586), .A4(G113), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n581), .A2(new_n585), .A3(new_n420), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n578), .A2(new_n580), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n210), .B1(new_n324), .B2(new_n280), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n271), .A2(G125), .ZN(new_n591));
  INV_X1    g405(.A(G224), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G953), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT7), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n581), .A2(new_n585), .A3(new_n587), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT86), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n598), .A2(new_n599), .A3(new_n416), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n598), .B2(new_n416), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n581), .A2(new_n420), .A3(new_n584), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n579), .B(KEYINPUT8), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n597), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT87), .B1(new_n607), .B2(KEYINPUT7), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(KEYINPUT87), .A3(KEYINPUT7), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n229), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT88), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n590), .A2(new_n591), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n594), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT85), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n578), .A2(new_n617), .A3(new_n588), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n578), .B2(new_n588), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n579), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT6), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n620), .B2(new_n589), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n589), .A2(new_n596), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n598), .A2(new_n416), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT86), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n598), .A2(new_n599), .A3(new_n416), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n602), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n605), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n607), .A2(KEYINPUT87), .A3(KEYINPUT7), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n608), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(KEYINPUT88), .A3(new_n229), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n614), .A2(new_n624), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT89), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n614), .A2(new_n624), .A3(KEYINPUT89), .A4(new_n635), .ZN(new_n639));
  OAI21_X1  g453(.A(G210), .B1(G237), .B2(G902), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT90), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT91), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n641), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n614), .A2(new_n624), .A3(new_n644), .A4(new_n635), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n575), .B(new_n577), .C1(new_n643), .C2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n391), .A2(new_n567), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G101), .ZN(G3));
  AOI21_X1  g462(.A(KEYINPUT88), .B1(new_n634), .B2(new_n229), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n613), .B(G902), .C1(new_n631), .C2(new_n633), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n644), .B1(new_n651), .B2(new_n624), .ZN(new_n652));
  INV_X1    g466(.A(new_n645), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n576), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n575), .ZN(new_n655));
  AOI21_X1  g469(.A(G478), .B1(new_n558), .B2(new_n229), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT33), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n557), .B2(new_n550), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n551), .A2(KEYINPUT33), .A3(new_n552), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n656), .B1(new_n660), .B2(G478), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n526), .B2(new_n565), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(G472), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n362), .B2(new_n229), .ZN(new_n665));
  INV_X1    g479(.A(new_n363), .ZN(new_n666));
  INV_X1    g480(.A(new_n361), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n360), .B1(new_n331), .B2(KEYINPUT31), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n372), .A2(new_n378), .ZN(new_n670));
  INV_X1    g484(.A(new_n331), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n670), .A2(new_n334), .B1(new_n671), .B2(new_n358), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n666), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT98), .B1(new_n665), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n467), .A2(new_n243), .A3(new_n471), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  AOI21_X1  g490(.A(G902), .B1(new_n669), .B2(new_n672), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n676), .B1(new_n677), .B2(new_n664), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n663), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT34), .B(G104), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  INV_X1    g496(.A(new_n561), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT93), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n522), .B1(new_n507), .B2(new_n516), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI22_X1  g500(.A1(new_n525), .A2(new_n524), .B1(new_n686), .B2(new_n476), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n687), .A2(new_n565), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n655), .A2(new_n683), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n679), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT99), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT35), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n399), .ZN(G9));
  NAND2_X1  g507(.A1(new_n235), .A2(new_n229), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT25), .ZN(new_n695));
  INV_X1    g509(.A(new_n241), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n230), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n220), .A2(new_n224), .ZN(new_n698));
  INV_X1    g512(.A(new_n190), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(KEYINPUT36), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n231), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n674), .A2(new_n678), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT100), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n674), .A2(new_n678), .A3(new_n707), .A4(new_n704), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(new_n567), .A3(new_n646), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT37), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n198), .ZN(G12));
  NAND2_X1  g525(.A1(new_n362), .A2(new_n363), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT32), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n362), .A2(KEYINPUT32), .A3(new_n363), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n390), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n472), .A2(new_n703), .ZN(new_n717));
  INV_X1    g531(.A(G900), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n572), .B1(new_n718), .B2(new_n574), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n565), .A2(new_n683), .A3(new_n687), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n636), .A2(new_n641), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n577), .B1(new_n722), .B2(new_n645), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n716), .A2(new_n717), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  AOI21_X1  g539(.A(KEYINPUT89), .B1(new_n651), .B2(new_n624), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n639), .A2(new_n642), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n645), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT38), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n643), .A2(KEYINPUT38), .A3(new_n645), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n472), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n719), .B(KEYINPUT39), .Z(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n732), .B1(KEYINPUT40), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n473), .B1(new_n684), .B2(new_n685), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n517), .B1(new_n737), .B2(KEYINPUT20), .ZN(new_n738));
  INV_X1    g552(.A(new_n565), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n561), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n735), .B2(KEYINPUT40), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n577), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n384), .A2(new_n353), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n229), .B1(new_n744), .B2(new_n321), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n357), .A2(new_n334), .ZN(new_n746));
  OAI21_X1  g560(.A(G472), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n714), .A2(new_n715), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n736), .A2(new_n743), .A3(new_n703), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G143), .ZN(G45));
  INV_X1    g564(.A(new_n661), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n751), .B(new_n720), .C1(new_n738), .C2(new_n739), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n716), .A2(new_n717), .A3(new_n753), .A4(new_n723), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G146), .ZN(G48));
  OAI21_X1  g569(.A(new_n229), .B1(new_n441), .B2(new_n453), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT101), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(G469), .ZN(new_n758));
  OAI221_X1 g572(.A(new_n229), .B1(KEYINPUT101), .B2(new_n392), .C1(new_n441), .C2(new_n453), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n471), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n716), .A2(new_n243), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n663), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT41), .B(G113), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G15));
  NOR2_X1   g579(.A1(new_n689), .A2(new_n762), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n290), .ZN(G18));
  NOR2_X1   g581(.A1(new_n654), .A2(new_n760), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n704), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n566), .A2(new_n575), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n716), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n199), .ZN(G21));
  INV_X1    g587(.A(new_n575), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n741), .A2(new_n774), .A3(new_n723), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n359), .B(new_n332), .C1(new_n386), .C2(new_n321), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n363), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n665), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n761), .A3(new_n243), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n533), .ZN(G24));
  NOR3_X1   g595(.A1(new_n665), .A2(new_n703), .A3(new_n777), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT102), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n752), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT102), .B1(new_n662), .B2(new_n720), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n768), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G125), .ZN(G27));
  INV_X1    g601(.A(KEYINPUT103), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n465), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT103), .A4(G469), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n454), .A3(new_n466), .A4(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n791), .A2(KEYINPUT104), .A3(new_n471), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT104), .B1(new_n791), .B2(new_n471), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n752), .A2(new_n783), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n662), .A2(KEYINPUT102), .A3(new_n720), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n643), .A2(new_n576), .A3(new_n645), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n794), .A2(new_n391), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT42), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n792), .A2(new_n793), .A3(new_n798), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT42), .A3(new_n391), .A4(new_n797), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  INV_X1    g620(.A(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n716), .A2(new_n243), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n721), .A2(KEYINPUT105), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n721), .A2(KEYINPUT105), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G134), .ZN(G36));
  NOR2_X1   g627(.A1(new_n665), .A2(KEYINPUT98), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n712), .B1(new_n677), .B2(new_n664), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(KEYINPUT98), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n704), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n740), .A2(new_n751), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT106), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT43), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT107), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n821), .B(KEYINPUT43), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT107), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n818), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n798), .B1(new_n828), .B2(KEYINPUT44), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n463), .A2(new_n464), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT45), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(G469), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(KEYINPUT46), .A3(new_n466), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT46), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n834), .B(G469), .C1(new_n831), .C2(G902), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n454), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(new_n471), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n734), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT108), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n825), .A2(new_n827), .ZN(new_n840));
  INV_X1    g654(.A(new_n818), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT44), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n828), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n829), .B(new_n838), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(G137), .ZN(G39));
  INV_X1    g661(.A(KEYINPUT47), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n837), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n836), .A2(new_n471), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT47), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n716), .A2(new_n243), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n798), .A2(new_n752), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT109), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n854), .A2(KEYINPUT109), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n851), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT110), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(G140), .ZN(G42));
  NAND3_X1  g673(.A1(new_n732), .A2(new_n577), .A3(new_n761), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT118), .Z(new_n861));
  AND4_X1   g675(.A1(new_n243), .A2(new_n826), .A3(new_n572), .A4(new_n778), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(KEYINPUT50), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n826), .A2(new_n572), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n798), .A2(new_n760), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n782), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n849), .A2(new_n851), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n758), .A2(new_n470), .A3(new_n759), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n798), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n748), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n243), .A2(new_n869), .A3(new_n572), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n526), .A2(new_n565), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n751), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n873), .A2(new_n862), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n867), .A2(new_n870), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n868), .A2(new_n391), .A3(new_n869), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT48), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n571), .B1(new_n875), .B2(new_n662), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n881), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n862), .A2(new_n768), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT112), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n876), .B2(new_n751), .ZN(new_n892));
  AOI211_X1 g706(.A(KEYINPUT112), .B(new_n661), .C1(new_n526), .C2(new_n565), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n728), .A2(new_n774), .A3(new_n576), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n679), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n567), .A2(new_n774), .A3(new_n576), .A4(new_n728), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n808), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT113), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n751), .B1(new_n738), .B2(new_n739), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT112), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n662), .A2(new_n891), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n816), .A2(new_n646), .A3(new_n675), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n647), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n740), .A2(new_n683), .ZN(new_n907));
  OR3_X1    g721(.A1(new_n679), .A2(new_n895), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n899), .A2(new_n709), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n709), .A2(new_n908), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(KEYINPUT114), .A3(new_n899), .A4(new_n906), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n786), .A2(new_n724), .A3(new_n754), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n748), .A2(new_n703), .A3(new_n720), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n723), .A2(new_n876), .A3(new_n683), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n791), .A2(new_n471), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT52), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n654), .B1(new_n366), .B2(new_n390), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n921), .B(new_n717), .C1(new_n721), .C2(new_n753), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n917), .A2(new_n918), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n703), .A3(new_n720), .A4(new_n748), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT52), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n922), .A2(new_n924), .A3(new_n925), .A4(new_n786), .ZN(new_n926));
  OAI22_X1  g740(.A1(new_n689), .A2(new_n762), .B1(new_n769), .B2(new_n771), .ZN(new_n927));
  OAI22_X1  g741(.A1(new_n663), .A2(new_n762), .B1(new_n775), .B2(new_n779), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n805), .A2(new_n920), .A3(new_n926), .A4(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n812), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n797), .A2(new_n782), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n807), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n688), .A2(new_n561), .A3(new_n720), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT115), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n716), .A2(new_n937), .A3(new_n717), .A4(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n934), .B1(new_n939), .B2(new_n799), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n914), .A2(new_n932), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n920), .A2(new_n926), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT116), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT54), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT54), .ZN(new_n948));
  INV_X1    g762(.A(new_n940), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n911), .B2(new_n913), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT117), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT53), .B1(new_n930), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n932), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n950), .B2(new_n932), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n889), .A2(new_n890), .A3(new_n947), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(G952), .B2(G953), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n758), .A2(new_n759), .ZN(new_n959));
  AOI211_X1 g773(.A(new_n577), .B(new_n244), .C1(KEYINPUT49), .C2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n960), .B(new_n874), .C1(KEYINPUT49), .C2(new_n959), .ZN(new_n961));
  INV_X1    g775(.A(new_n732), .ZN(new_n962));
  NOR4_X1   g776(.A1(new_n961), .A2(new_n470), .A3(new_n962), .A4(new_n819), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n958), .A2(new_n964), .ZN(G75));
  NOR3_X1   g779(.A1(new_n954), .A2(new_n955), .A3(new_n229), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT56), .B1(new_n966), .B2(new_n641), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n622), .A2(new_n623), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(new_n616), .Z(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(KEYINPUT119), .Z(new_n972));
  AOI211_X1 g786(.A(KEYINPUT56), .B(new_n972), .C1(new_n966), .C2(new_n642), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n187), .A2(G952), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(G51));
  INV_X1    g789(.A(KEYINPUT120), .ZN(new_n976));
  INV_X1    g790(.A(new_n952), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n941), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(KEYINPUT54), .A3(new_n953), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n956), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(KEYINPUT120), .B(new_n948), .C1(new_n954), .C2(new_n955), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n466), .B(KEYINPUT57), .Z(new_n982));
  NAND3_X1  g796(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n441), .B2(new_n453), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n966), .A2(G469), .A3(new_n831), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n974), .B1(new_n984), .B2(new_n985), .ZN(G54));
  NAND3_X1  g800(.A1(new_n966), .A2(KEYINPUT58), .A3(G475), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n686), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n686), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n989), .A3(new_n974), .ZN(G60));
  NAND2_X1  g804(.A1(new_n658), .A2(new_n659), .ZN(new_n991));
  NAND2_X1  g805(.A1(G478), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT59), .Z(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  AND4_X1   g808(.A1(new_n991), .A2(new_n980), .A3(new_n981), .A4(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n974), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n947), .B2(new_n956), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n991), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n995), .A2(new_n998), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT60), .Z(new_n1001));
  NAND3_X1  g815(.A1(new_n978), .A2(new_n953), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n235), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n1002), .A2(KEYINPUT122), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT122), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n978), .A2(new_n701), .A3(new_n953), .A4(new_n1001), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n996), .A2(KEYINPUT61), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1006), .A2(new_n996), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(KEYINPUT123), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1010), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1006), .A2(new_n996), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT123), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT122), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1012), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1002), .A2(KEYINPUT122), .A3(new_n1003), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1018), .B(new_n1019), .C1(new_n1023), .C2(new_n1008), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1014), .A2(new_n1024), .ZN(G66));
  OAI21_X1  g839(.A(G953), .B1(new_n573), .B2(new_n592), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n914), .A2(new_n929), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1026), .B1(new_n1028), .B2(G953), .ZN(new_n1029));
  INV_X1    g843(.A(G898), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n968), .B1(new_n1030), .B2(G953), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1029), .B(new_n1031), .Z(G69));
  AOI21_X1  g846(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n838), .A2(new_n391), .A3(new_n723), .A4(new_n741), .ZN(new_n1035));
  AND4_X1   g849(.A1(new_n805), .A2(new_n1035), .A3(new_n812), .A4(new_n857), .ZN(new_n1036));
  INV_X1    g850(.A(new_n915), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n846), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1038), .A2(G953), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G900), .A2(G953), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n356), .B(KEYINPUT124), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1041), .B(new_n503), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n749), .A2(new_n1037), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT62), .Z(new_n1045));
  AOI211_X1 g859(.A(new_n735), .B(new_n808), .C1(new_n907), .C2(new_n894), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n799), .ZN(new_n1047));
  AND3_X1   g861(.A1(new_n846), .A2(KEYINPUT126), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(KEYINPUT126), .B1(new_n846), .B2(new_n1047), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n857), .B(new_n1045), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AND2_X1   g864(.A1(new_n1050), .A2(new_n187), .ZN(new_n1051));
  XOR2_X1   g865(.A(new_n1042), .B(KEYINPUT125), .Z(new_n1052));
  OAI211_X1 g866(.A(new_n1034), .B(new_n1043), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1052), .B1(new_n1050), .B2(new_n187), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1043), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1033), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1053), .A2(new_n1056), .ZN(G72));
  NAND2_X1  g871(.A1(G472), .A2(G902), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT63), .Z(new_n1059));
  OAI21_X1  g873(.A(new_n1059), .B1(new_n1038), .B2(new_n1027), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1060), .A2(new_n334), .A3(new_n357), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n367), .A2(new_n331), .A3(new_n382), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1062), .A2(new_n1059), .ZN(new_n1063));
  XNOR2_X1  g877(.A(new_n1063), .B(KEYINPUT127), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1064), .B1(new_n945), .B2(new_n946), .ZN(new_n1065));
  NAND3_X1  g879(.A1(new_n1061), .A2(new_n996), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1059), .B1(new_n1050), .B2(new_n1027), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1066), .B1(new_n1067), .B2(new_n746), .ZN(G57));
endmodule


