

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766;

  XNOR2_X1 U376 ( .A(n609), .B(KEYINPUT6), .ZN(n602) );
  XNOR2_X1 U377 ( .A(n432), .B(n431), .ZN(n609) );
  OR2_X1 U378 ( .A1(n733), .A2(G902), .ZN(n400) );
  XNOR2_X1 U379 ( .A(n375), .B(n354), .ZN(n428) );
  XNOR2_X1 U380 ( .A(n427), .B(G101), .ZN(n354) );
  XNOR2_X1 U381 ( .A(n374), .B(n424), .ZN(n488) );
  XNOR2_X1 U382 ( .A(G143), .B(KEYINPUT81), .ZN(n374) );
  OR2_X4 U383 ( .A1(n692), .A2(n615), .ZN(n382) );
  AND2_X4 U384 ( .A1(n681), .A2(n385), .ZN(n386) );
  XNOR2_X2 U385 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X2 U386 ( .A(n441), .B(G902), .ZN(n675) );
  BUF_X2 U387 ( .A(n617), .Z(n694) );
  BUF_X1 U388 ( .A(n620), .Z(n696) );
  XNOR2_X1 U389 ( .A(n705), .B(KEYINPUT64), .ZN(n355) );
  INV_X2 U390 ( .A(n387), .ZN(n388) );
  AND2_X2 U391 ( .A1(n600), .A2(n599), .ZN(n616) );
  XNOR2_X2 U392 ( .A(n419), .B(n418), .ZN(n421) );
  INV_X1 U393 ( .A(n739), .ZN(n356) );
  INV_X4 U394 ( .A(G953), .ZN(n761) );
  INV_X1 U395 ( .A(KEYINPUT56), .ZN(n357) );
  NOR2_X1 U396 ( .A1(n766), .A2(n765), .ZN(n521) );
  XNOR2_X1 U397 ( .A(n527), .B(KEYINPUT80), .ZN(n722) );
  XNOR2_X1 U398 ( .A(n520), .B(n519), .ZN(n765) );
  NOR2_X1 U399 ( .A1(n542), .A2(n517), .ZN(n518) );
  AND2_X1 U400 ( .A1(n588), .A2(n587), .ZN(n606) );
  AND2_X1 U401 ( .A1(n404), .A2(n380), .ZN(n381) );
  XNOR2_X1 U402 ( .A(n428), .B(n429), .ZN(n687) );
  XNOR2_X1 U403 ( .A(n460), .B(n378), .ZN(n397) );
  XOR2_X1 U404 ( .A(n745), .B(KEYINPUT69), .Z(n378) );
  XNOR2_X1 U405 ( .A(n488), .B(n373), .ZN(n460) );
  XNOR2_X1 U406 ( .A(n457), .B(G110), .ZN(n459) );
  XOR2_X1 U407 ( .A(G140), .B(G104), .Z(n471) );
  XNOR2_X1 U408 ( .A(KEYINPUT4), .B(G101), .ZN(n373) );
  INV_X2 U409 ( .A(KEYINPUT74), .ZN(n457) );
  XNOR2_X1 U410 ( .A(G128), .B(G119), .ZN(n434) );
  XNOR2_X1 U411 ( .A(G107), .B(G104), .ZN(n458) );
  XOR2_X1 U412 ( .A(G137), .B(G140), .Z(n461) );
  BUF_X1 U413 ( .A(KEYINPUT63), .Z(n690) );
  XOR2_X1 U414 ( .A(G113), .B(G119), .Z(n420) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(G51) );
  NAND2_X1 U416 ( .A1(n362), .A2(n356), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(KEYINPUT121), .ZN(G63) );
  NAND2_X1 U418 ( .A1(n364), .A2(n356), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n690), .ZN(G57) );
  NAND2_X1 U420 ( .A1(n366), .A2(n356), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n355), .ZN(G60) );
  NAND2_X1 U422 ( .A1(n368), .A2(n356), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n396), .B(n397), .ZN(n376) );
  XNOR2_X2 U424 ( .A(n746), .B(n503), .ZN(n396) );
  XNOR2_X1 U425 ( .A(n711), .B(n363), .ZN(n362) );
  INV_X1 U426 ( .A(n710), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n684), .B(n365), .ZN(n364) );
  INV_X1 U428 ( .A(n683), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n689), .B(n367), .ZN(n366) );
  INV_X1 U430 ( .A(n688), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n704), .B(n369), .ZN(n368) );
  INV_X1 U432 ( .A(n703), .ZN(n369) );
  XNOR2_X2 U433 ( .A(n371), .B(n370), .ZN(n746) );
  INV_X1 U434 ( .A(n502), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n464), .ZN(n423) );
  XNOR2_X2 U436 ( .A(n421), .B(n372), .ZN(n371) );
  INV_X1 U437 ( .A(n420), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n488), .B(KEYINPUT4), .ZN(n375) );
  NOR2_X1 U439 ( .A1(n535), .A2(n642), .ZN(n610) );
  XNOR2_X1 U440 ( .A(n396), .B(n397), .ZN(n706) );
  XNOR2_X2 U441 ( .A(n392), .B(KEYINPUT22), .ZN(n403) );
  XNOR2_X1 U442 ( .A(n479), .B(n393), .ZN(n755) );
  INV_X1 U443 ( .A(n461), .ZN(n393) );
  XNOR2_X1 U444 ( .A(n478), .B(n395), .ZN(n702) );
  XNOR2_X1 U445 ( .A(n479), .B(n477), .ZN(n395) );
  NAND2_X1 U446 ( .A1(n680), .A2(n759), .ZN(n385) );
  NAND2_X1 U447 ( .A1(n678), .A2(n677), .ZN(n681) );
  AND2_X1 U448 ( .A1(KEYINPUT2), .A2(n628), .ZN(n680) );
  XNOR2_X1 U449 ( .A(n531), .B(n394), .ZN(n533) );
  INV_X1 U450 ( .A(KEYINPUT72), .ZN(n394) );
  NOR2_X1 U451 ( .A1(n722), .A2(n530), .ZN(n531) );
  NOR2_X1 U452 ( .A1(n724), .A2(n727), .ZN(n637) );
  INV_X1 U453 ( .A(G128), .ZN(n424) );
  NAND2_X1 U454 ( .A1(n507), .A2(n675), .ZN(n415) );
  XNOR2_X1 U455 ( .A(G131), .B(G134), .ZN(n753) );
  XNOR2_X1 U456 ( .A(G116), .B(G134), .ZN(n486) );
  XOR2_X1 U457 ( .A(G122), .B(G107), .Z(n487) );
  XNOR2_X1 U458 ( .A(G113), .B(G122), .ZN(n472) );
  XOR2_X1 U459 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n473) );
  XNOR2_X1 U460 ( .A(KEYINPUT18), .B(KEYINPUT77), .ZN(n497) );
  XNOR2_X1 U461 ( .A(KEYINPUT94), .B(KEYINPUT17), .ZN(n498) );
  OR2_X1 U462 ( .A1(n632), .A2(KEYINPUT90), .ZN(n409) );
  OR2_X1 U463 ( .A1(n706), .A2(n405), .ZN(n410) );
  OR2_X1 U464 ( .A1(n414), .A2(n406), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n501), .B(G122), .ZN(n502) );
  XOR2_X1 U466 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n501) );
  INV_X1 U467 ( .A(KEYINPUT28), .ZN(n389) );
  XOR2_X1 U468 ( .A(KEYINPUT62), .B(n687), .Z(n688) );
  XNOR2_X1 U469 ( .A(n755), .B(KEYINPUT23), .ZN(n440) );
  XOR2_X1 U470 ( .A(KEYINPUT120), .B(n682), .Z(n683) );
  XOR2_X1 U471 ( .A(KEYINPUT59), .B(n702), .Z(n703) );
  XNOR2_X1 U472 ( .A(n686), .B(KEYINPUT93), .ZN(n739) );
  XNOR2_X1 U473 ( .A(KEYINPUT104), .B(n529), .ZN(n718) );
  OR2_X1 U474 ( .A1(n635), .A2(n575), .ZN(n379) );
  AND2_X1 U475 ( .A1(n632), .A2(KEYINPUT90), .ZN(n380) );
  XOR2_X1 U476 ( .A(n574), .B(KEYINPUT0), .Z(n383) );
  XOR2_X1 U477 ( .A(KEYINPUT87), .B(KEYINPUT45), .Z(n384) );
  XNOR2_X1 U478 ( .A(n709), .B(n708), .ZN(n710) );
  BUF_X1 U479 ( .A(n679), .Z(n628) );
  INV_X1 U480 ( .A(n386), .ZN(n387) );
  NOR2_X1 U481 ( .A1(n381), .A2(n408), .ZN(n398) );
  XNOR2_X1 U482 ( .A(n390), .B(n389), .ZN(n469) );
  NOR2_X1 U483 ( .A1(n537), .A2(n609), .ZN(n390) );
  NOR2_X1 U484 ( .A1(n391), .A2(n696), .ZN(n624) );
  NAND2_X1 U485 ( .A1(n618), .A2(n619), .ZN(n391) );
  INV_X1 U486 ( .A(n667), .ZN(n401) );
  XNOR2_X2 U487 ( .A(n402), .B(n591), .ZN(n667) );
  NOR2_X2 U488 ( .A1(n607), .A2(n379), .ZN(n392) );
  NAND2_X1 U489 ( .A1(n413), .A2(n415), .ZN(n404) );
  NAND2_X1 U490 ( .A1(n410), .A2(n409), .ZN(n408) );
  XNOR2_X2 U491 ( .A(n416), .B(n383), .ZN(n607) );
  NOR2_X2 U492 ( .A1(n573), .A2(n572), .ZN(n416) );
  NAND2_X1 U493 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U494 ( .A(n627), .B(n384), .ZN(n679) );
  XNOR2_X2 U495 ( .A(n608), .B(KEYINPUT31), .ZN(n726) );
  OR2_X2 U496 ( .A1(n726), .A2(n713), .ZN(n613) );
  XNOR2_X2 U497 ( .A(n538), .B(KEYINPUT19), .ZN(n573) );
  NAND2_X2 U498 ( .A1(n398), .A2(n399), .ZN(n538) );
  XNOR2_X1 U499 ( .A(n397), .B(n466), .ZN(n733) );
  NAND2_X1 U500 ( .A1(n407), .A2(n411), .ZN(n399) );
  XNOR2_X2 U501 ( .A(n535), .B(n534), .ZN(n588) );
  XNOR2_X2 U502 ( .A(n400), .B(n467), .ZN(n535) );
  NAND2_X1 U503 ( .A1(n401), .A2(n592), .ZN(n595) );
  NAND2_X1 U504 ( .A1(n606), .A2(n602), .ZN(n402) );
  NAND2_X1 U505 ( .A1(n403), .A2(n583), .ZN(n584) );
  AND2_X2 U506 ( .A1(n403), .A2(n641), .ZN(n604) );
  INV_X1 U507 ( .A(n404), .ZN(n411) );
  OR2_X1 U508 ( .A1(n706), .A2(n414), .ZN(n412) );
  INV_X1 U509 ( .A(n380), .ZN(n406) );
  NAND2_X1 U510 ( .A1(n411), .A2(n412), .ZN(n522) );
  AND2_X1 U511 ( .A1(n412), .A2(n523), .ZN(n407) );
  NAND2_X1 U512 ( .A1(n376), .A2(n507), .ZN(n413) );
  OR2_X1 U513 ( .A1(n507), .A2(n675), .ZN(n414) );
  NOR2_X1 U514 ( .A1(n616), .A2(n382), .ZN(n626) );
  NOR2_X1 U515 ( .A1(n566), .A2(n718), .ZN(n417) );
  AND2_X1 U516 ( .A1(n695), .A2(KEYINPUT44), .ZN(n619) );
  INV_X1 U517 ( .A(KEYINPUT48), .ZN(n555) );
  XNOR2_X1 U518 ( .A(n555), .B(KEYINPUT65), .ZN(n556) );
  XNOR2_X1 U519 ( .A(n557), .B(n556), .ZN(n563) );
  INV_X1 U520 ( .A(KEYINPUT117), .ZN(n670) );
  XNOR2_X1 U521 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n519) );
  XNOR2_X1 U522 ( .A(n672), .B(n671), .ZN(G75) );
  INV_X1 U523 ( .A(KEYINPUT88), .ZN(n565) );
  XNOR2_X2 U524 ( .A(G116), .B(KEYINPUT67), .ZN(n419) );
  XNOR2_X2 U525 ( .A(KEYINPUT68), .B(KEYINPUT3), .ZN(n418) );
  XNOR2_X1 U526 ( .A(G146), .B(n753), .ZN(n464) );
  NOR2_X1 U527 ( .A1(G953), .A2(G237), .ZN(n476) );
  NAND2_X1 U528 ( .A1(n476), .A2(G210), .ZN(n422) );
  XNOR2_X1 U529 ( .A(n423), .B(n422), .ZN(n429) );
  XOR2_X1 U530 ( .A(KEYINPUT101), .B(KEYINPUT5), .Z(n426) );
  XNOR2_X1 U531 ( .A(G137), .B(KEYINPUT100), .ZN(n425) );
  XNOR2_X1 U532 ( .A(n426), .B(n425), .ZN(n427) );
  INV_X1 U533 ( .A(G902), .ZN(n505) );
  NAND2_X1 U534 ( .A1(n687), .A2(n505), .ZN(n432) );
  INV_X1 U535 ( .A(KEYINPUT102), .ZN(n430) );
  XNOR2_X1 U536 ( .A(n430), .B(G472), .ZN(n431) );
  XNOR2_X2 U537 ( .A(G146), .B(G125), .ZN(n495) );
  XNOR2_X1 U538 ( .A(n495), .B(KEYINPUT10), .ZN(n479) );
  NAND2_X1 U539 ( .A1(G234), .A2(n761), .ZN(n433) );
  XOR2_X1 U540 ( .A(KEYINPUT8), .B(n433), .Z(n483) );
  NAND2_X1 U541 ( .A1(n483), .A2(G221), .ZN(n438) );
  XOR2_X1 U542 ( .A(KEYINPUT75), .B(G110), .Z(n435) );
  XNOR2_X1 U543 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U544 ( .A(n436), .B(KEYINPUT24), .Z(n437) );
  XNOR2_X1 U545 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U546 ( .A(n440), .B(n439), .ZN(n698) );
  NAND2_X1 U547 ( .A1(n698), .A2(n505), .ZN(n448) );
  XOR2_X1 U548 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n444) );
  INV_X1 U549 ( .A(KEYINPUT15), .ZN(n441) );
  INV_X1 U550 ( .A(n675), .ZN(n442) );
  NAND2_X1 U551 ( .A1(G234), .A2(n442), .ZN(n443) );
  XNOR2_X1 U552 ( .A(n444), .B(n443), .ZN(n453) );
  NAND2_X1 U553 ( .A1(n453), .A2(G217), .ZN(n446) );
  XOR2_X1 U554 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n445) );
  XNOR2_X1 U555 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X2 U556 ( .A(n448), .B(n447), .ZN(n580) );
  NOR2_X1 U557 ( .A1(G900), .A2(n761), .ZN(n449) );
  NAND2_X1 U558 ( .A1(n449), .A2(G902), .ZN(n450) );
  NAND2_X1 U559 ( .A1(n761), .A2(G952), .ZN(n569) );
  NAND2_X1 U560 ( .A1(n450), .A2(n569), .ZN(n452) );
  NAND2_X1 U561 ( .A1(G237), .A2(G234), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n451), .B(KEYINPUT14), .ZN(n631) );
  NAND2_X1 U563 ( .A1(n452), .A2(n631), .ZN(n514) );
  NOR2_X1 U564 ( .A1(n580), .A2(n514), .ZN(n456) );
  NAND2_X1 U565 ( .A1(n453), .A2(G221), .ZN(n455) );
  XNOR2_X1 U566 ( .A(KEYINPUT99), .B(KEYINPUT21), .ZN(n454) );
  XNOR2_X1 U567 ( .A(n455), .B(n454), .ZN(n645) );
  NAND2_X1 U568 ( .A1(n456), .A2(n645), .ZN(n537) );
  XNOR2_X1 U569 ( .A(n459), .B(n458), .ZN(n745) );
  XOR2_X1 U570 ( .A(n461), .B(KEYINPUT76), .Z(n463) );
  NAND2_X1 U571 ( .A1(G227), .A2(n761), .ZN(n462) );
  XNOR2_X1 U572 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U573 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U574 ( .A(KEYINPUT66), .B(G469), .Z(n467) );
  XOR2_X1 U575 ( .A(n535), .B(KEYINPUT111), .Z(n468) );
  NOR2_X1 U576 ( .A1(n469), .A2(n468), .ZN(n525) );
  INV_X1 U577 ( .A(n525), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G143), .B(G131), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n471), .B(n470), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U581 ( .A(n475), .B(n474), .Z(n478) );
  NAND2_X1 U582 ( .A1(G214), .A2(n476), .ZN(n477) );
  NOR2_X1 U583 ( .A1(G902), .A2(n702), .ZN(n481) );
  XNOR2_X1 U584 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U586 ( .A(n482), .B(G475), .ZN(n544) );
  XOR2_X1 U587 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n485) );
  NAND2_X1 U588 ( .A1(G217), .A2(n483), .ZN(n484) );
  XNOR2_X1 U589 ( .A(n485), .B(n484), .ZN(n492) );
  XNOR2_X1 U590 ( .A(n487), .B(n486), .ZN(n490) );
  INV_X1 U591 ( .A(n488), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n492), .B(n491), .ZN(n682) );
  NAND2_X1 U594 ( .A1(n682), .A2(n505), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n493), .B(G478), .ZN(n528) );
  INV_X1 U596 ( .A(n528), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n635) );
  NAND2_X1 U598 ( .A1(n761), .A2(G224), .ZN(n494) );
  XNOR2_X1 U599 ( .A(n494), .B(KEYINPUT78), .ZN(n496) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U601 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U602 ( .A(n500), .B(n499), .ZN(n503) );
  INV_X1 U603 ( .A(G237), .ZN(n504) );
  NAND2_X1 U604 ( .A1(n505), .A2(n504), .ZN(n509) );
  NAND2_X1 U605 ( .A1(n509), .A2(G210), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n506), .B(KEYINPUT95), .ZN(n507) );
  XOR2_X1 U607 ( .A(KEYINPUT38), .B(KEYINPUT73), .Z(n508) );
  XNOR2_X1 U608 ( .A(n522), .B(n508), .ZN(n516) );
  INV_X1 U609 ( .A(n516), .ZN(n633) );
  NAND2_X1 U610 ( .A1(n509), .A2(G214), .ZN(n632) );
  NAND2_X1 U611 ( .A1(n633), .A2(n632), .ZN(n636) );
  NOR2_X1 U612 ( .A1(n635), .A2(n636), .ZN(n510) );
  XNOR2_X1 U613 ( .A(KEYINPUT41), .B(n510), .ZN(n666) );
  NOR2_X1 U614 ( .A1(n511), .A2(n666), .ZN(n512) );
  XNOR2_X1 U615 ( .A(n512), .B(KEYINPUT42), .ZN(n766) );
  OR2_X1 U616 ( .A1(n544), .A2(n528), .ZN(n721) );
  INV_X1 U617 ( .A(n609), .ZN(n648) );
  NAND2_X1 U618 ( .A1(n648), .A2(n632), .ZN(n513) );
  XNOR2_X1 U619 ( .A(n513), .B(KEYINPUT30), .ZN(n542) );
  INV_X1 U620 ( .A(n514), .ZN(n515) );
  NAND2_X1 U621 ( .A1(n580), .A2(n645), .ZN(n642) );
  NAND2_X1 U622 ( .A1(n515), .A2(n610), .ZN(n541) );
  OR2_X1 U623 ( .A1(n541), .A2(n516), .ZN(n517) );
  XNOR2_X1 U624 ( .A(n518), .B(KEYINPUT39), .ZN(n566) );
  NOR2_X1 U625 ( .A1(n721), .A2(n566), .ZN(n520) );
  XNOR2_X1 U626 ( .A(n521), .B(KEYINPUT46), .ZN(n554) );
  INV_X1 U627 ( .A(KEYINPUT90), .ZN(n523) );
  BUF_X1 U628 ( .A(n573), .Z(n524) );
  INV_X1 U629 ( .A(n524), .ZN(n526) );
  NAND2_X1 U630 ( .A1(n526), .A2(n525), .ZN(n527) );
  INV_X1 U631 ( .A(n721), .ZN(n724) );
  NAND2_X1 U632 ( .A1(n528), .A2(n544), .ZN(n529) );
  INV_X1 U633 ( .A(n718), .ZN(n727) );
  OR2_X1 U634 ( .A1(KEYINPUT47), .A2(n637), .ZN(n530) );
  NAND2_X1 U635 ( .A1(n722), .A2(KEYINPUT47), .ZN(n532) );
  AND2_X1 U636 ( .A1(n533), .A2(n532), .ZN(n552) );
  INV_X1 U637 ( .A(KEYINPUT1), .ZN(n534) );
  INV_X1 U638 ( .A(n588), .ZN(n641) );
  NAND2_X1 U639 ( .A1(n724), .A2(n602), .ZN(n536) );
  NOR2_X1 U640 ( .A1(n537), .A2(n536), .ZN(n558) );
  NAND2_X1 U641 ( .A1(n558), .A2(n538), .ZN(n539) );
  XNOR2_X1 U642 ( .A(n539), .B(KEYINPUT36), .ZN(n540) );
  NOR2_X1 U643 ( .A1(n641), .A2(n540), .ZN(n729) );
  OR2_X1 U644 ( .A1(n542), .A2(n541), .ZN(n546) );
  NOR2_X1 U645 ( .A1(n544), .A2(n543), .ZN(n596) );
  INV_X1 U646 ( .A(n596), .ZN(n545) );
  NOR2_X1 U647 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U648 ( .A1(n547), .A2(n522), .ZN(n691) );
  NAND2_X1 U649 ( .A1(KEYINPUT47), .A2(n637), .ZN(n548) );
  NAND2_X1 U650 ( .A1(n691), .A2(n548), .ZN(n549) );
  XNOR2_X1 U651 ( .A(KEYINPUT82), .B(n549), .ZN(n550) );
  NOR2_X1 U652 ( .A1(n729), .A2(n550), .ZN(n551) );
  AND2_X1 U653 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U654 ( .A1(n554), .A2(n553), .ZN(n557) );
  XNOR2_X1 U655 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n561) );
  NAND2_X1 U656 ( .A1(n558), .A2(n632), .ZN(n559) );
  NOR2_X1 U657 ( .A1(n588), .A2(n559), .ZN(n560) );
  XNOR2_X1 U658 ( .A(n561), .B(n560), .ZN(n562) );
  NOR2_X1 U659 ( .A1(n562), .A2(n522), .ZN(n731) );
  NOR2_X1 U660 ( .A1(n563), .A2(n731), .ZN(n564) );
  XNOR2_X1 U661 ( .A(n565), .B(n564), .ZN(n567) );
  NOR2_X2 U662 ( .A1(n567), .A2(n417), .ZN(n759) );
  NOR2_X1 U663 ( .A1(G898), .A2(n761), .ZN(n568) );
  XNOR2_X1 U664 ( .A(KEYINPUT96), .B(n568), .ZN(n750) );
  NAND2_X1 U665 ( .A1(n750), .A2(G902), .ZN(n570) );
  NAND2_X1 U666 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U667 ( .A1(n571), .A2(n631), .ZN(n572) );
  INV_X1 U668 ( .A(KEYINPUT91), .ZN(n574) );
  INV_X1 U669 ( .A(n645), .ZN(n575) );
  INV_X1 U670 ( .A(n580), .ZN(n576) );
  AND2_X1 U671 ( .A1(n609), .A2(n576), .ZN(n577) );
  NAND2_X1 U672 ( .A1(n604), .A2(n577), .ZN(n579) );
  INV_X1 U673 ( .A(KEYINPUT108), .ZN(n578) );
  XNOR2_X2 U674 ( .A(n579), .B(n578), .ZN(n620) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT79), .ZN(n582) );
  XNOR2_X1 U676 ( .A(n580), .B(KEYINPUT106), .ZN(n644) );
  INV_X1 U677 ( .A(n644), .ZN(n601) );
  AND2_X1 U678 ( .A1(n588), .A2(n601), .ZN(n581) );
  AND2_X1 U679 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X2 U680 ( .A(n584), .B(KEYINPUT32), .ZN(n695) );
  INV_X1 U681 ( .A(KEYINPUT44), .ZN(n621) );
  NAND2_X1 U682 ( .A1(n695), .A2(n621), .ZN(n585) );
  OR2_X2 U683 ( .A1(n620), .A2(n585), .ZN(n586) );
  INV_X1 U684 ( .A(KEYINPUT89), .ZN(n622) );
  NAND2_X1 U685 ( .A1(n586), .A2(n622), .ZN(n600) );
  INV_X1 U686 ( .A(n607), .ZN(n592) );
  INV_X1 U687 ( .A(n642), .ZN(n587) );
  XOR2_X1 U688 ( .A(KEYINPUT109), .B(KEYINPUT33), .Z(n590) );
  INV_X1 U689 ( .A(KEYINPUT92), .ZN(n589) );
  XNOR2_X1 U690 ( .A(n590), .B(n589), .ZN(n591) );
  INV_X1 U691 ( .A(KEYINPUT70), .ZN(n593) );
  XNOR2_X1 U692 ( .A(n593), .B(KEYINPUT34), .ZN(n594) );
  XNOR2_X1 U693 ( .A(n595), .B(n594), .ZN(n597) );
  NAND2_X1 U694 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X2 U695 ( .A(n598), .B(KEYINPUT35), .ZN(n617) );
  INV_X1 U696 ( .A(n694), .ZN(n599) );
  NOR2_X1 U697 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U698 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U699 ( .A(n605), .B(KEYINPUT107), .ZN(n692) );
  NAND2_X1 U700 ( .A1(n606), .A2(n648), .ZN(n651) );
  OR2_X1 U701 ( .A1(n607), .A2(n651), .ZN(n608) );
  AND2_X1 U702 ( .A1(n610), .A2(n609), .ZN(n611) );
  AND2_X1 U703 ( .A1(n592), .A2(n611), .ZN(n713) );
  INV_X1 U704 ( .A(n637), .ZN(n612) );
  NAND2_X1 U705 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U706 ( .A(n614), .B(KEYINPUT105), .ZN(n615) );
  NAND2_X1 U707 ( .A1(n617), .A2(n622), .ZN(n618) );
  AND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n623) );
  OR2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n759), .A2(n628), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n629), .A2(KEYINPUT84), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT2), .ZN(n665) );
  INV_X1 U713 ( .A(n631), .ZN(n660) );
  NOR2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n639) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U718 ( .A1(n667), .A2(n640), .ZN(n657) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT50), .ZN(n650) );
  NOR2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U722 ( .A(KEYINPUT49), .B(n646), .Z(n647) );
  NOR2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n655), .A2(n666), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(KEYINPUT52), .ZN(n659) );
  NOR2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n661), .A2(G952), .ZN(n662) );
  XOR2_X1 U733 ( .A(KEYINPUT116), .B(n662), .Z(n663) );
  NOR2_X1 U734 ( .A1(G953), .A2(n663), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n670), .B(KEYINPUT53), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n679), .A2(n675), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n673), .B(KEYINPUT85), .ZN(n674) );
  NAND2_X1 U741 ( .A1(n674), .A2(n759), .ZN(n678) );
  XNOR2_X1 U742 ( .A(n675), .B(KEYINPUT86), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n676), .A2(KEYINPUT2), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n386), .A2(G478), .ZN(n684) );
  INV_X1 U745 ( .A(G952), .ZN(n685) );
  NAND2_X1 U746 ( .A1(n685), .A2(G953), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n386), .A2(G472), .ZN(n689) );
  XNOR2_X1 U748 ( .A(n691), .B(G143), .ZN(G45) );
  XOR2_X1 U749 ( .A(G101), .B(n692), .Z(G3) );
  XNOR2_X1 U750 ( .A(G122), .B(KEYINPUT127), .ZN(n693) );
  XNOR2_X1 U751 ( .A(n694), .B(n693), .ZN(G24) );
  XNOR2_X1 U752 ( .A(n695), .B(G119), .ZN(G21) );
  XOR2_X1 U753 ( .A(n696), .B(G110), .Z(G12) );
  NAND2_X1 U754 ( .A1(n388), .A2(G217), .ZN(n700) );
  XNOR2_X1 U755 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U758 ( .A1(n701), .A2(n739), .ZN(G66) );
  NAND2_X1 U759 ( .A1(n386), .A2(G475), .ZN(n704) );
  XNOR2_X1 U760 ( .A(KEYINPUT119), .B(KEYINPUT60), .ZN(n705) );
  NAND2_X1 U761 ( .A1(n386), .A2(G210), .ZN(n711) );
  BUF_X1 U762 ( .A(n376), .Z(n709) );
  XNOR2_X1 U763 ( .A(KEYINPUT83), .B(KEYINPUT54), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n707), .B(KEYINPUT55), .ZN(n708) );
  NAND2_X1 U765 ( .A1(n713), .A2(n724), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(G104), .ZN(G6) );
  XOR2_X1 U767 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n715) );
  NAND2_X1 U768 ( .A1(n713), .A2(n727), .ZN(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(n717) );
  XOR2_X1 U770 ( .A(G107), .B(KEYINPUT26), .Z(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(G9) );
  XNOR2_X1 U772 ( .A(G128), .B(KEYINPUT29), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n718), .A2(n722), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(G30) );
  NOR2_X1 U775 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U776 ( .A(G146), .B(n723), .Z(G48) );
  NAND2_X1 U777 ( .A1(n726), .A2(n724), .ZN(n725) );
  XNOR2_X1 U778 ( .A(n725), .B(G113), .ZN(G15) );
  NAND2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(G116), .ZN(G18) );
  XNOR2_X1 U781 ( .A(G125), .B(n729), .ZN(n730) );
  XNOR2_X1 U782 ( .A(n730), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U783 ( .A(G134), .B(n417), .Z(G36) );
  XOR2_X1 U784 ( .A(G140), .B(n731), .Z(n732) );
  XNOR2_X1 U785 ( .A(KEYINPUT114), .B(n732), .ZN(G42) );
  NAND2_X1 U786 ( .A1(n388), .A2(G469), .ZN(n737) );
  XOR2_X1 U787 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n735) );
  XNOR2_X1 U788 ( .A(n733), .B(KEYINPUT118), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(G54) );
  NAND2_X1 U791 ( .A1(n628), .A2(n761), .ZN(n744) );
  NAND2_X1 U792 ( .A1(G224), .A2(G953), .ZN(n740) );
  XNOR2_X1 U793 ( .A(n740), .B(KEYINPUT61), .ZN(n741) );
  XNOR2_X1 U794 ( .A(KEYINPUT124), .B(n741), .ZN(n742) );
  NAND2_X1 U795 ( .A1(n742), .A2(G898), .ZN(n743) );
  NAND2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n752) );
  XNOR2_X1 U797 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n747), .B(KEYINPUT125), .ZN(n748) );
  XNOR2_X1 U799 ( .A(n748), .B(G101), .ZN(n749) );
  NOR2_X1 U800 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(G69) );
  XNOR2_X1 U802 ( .A(n375), .B(n753), .ZN(n754) );
  XNOR2_X1 U803 ( .A(n755), .B(n754), .ZN(n760) );
  XOR2_X1 U804 ( .A(G227), .B(n760), .Z(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n757), .A2(G953), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n758), .B(KEYINPUT126), .ZN(n764) );
  XNOR2_X1 U808 ( .A(n760), .B(n759), .ZN(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U811 ( .A(n765), .B(G131), .Z(G33) );
  XOR2_X1 U812 ( .A(G137), .B(n766), .Z(G39) );
endmodule

