//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT66), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n193), .A3(new_n196), .A4(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(new_n202), .B2(new_n204), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR3_X1   g023(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n206), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n200), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n201), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G128), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n202), .A3(new_n204), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n191), .A2(new_n193), .A3(new_n223), .A4(new_n194), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n192), .A2(G134), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n194), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n222), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n213), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(KEYINPUT67), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n232), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT28), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n219), .A2(new_n221), .B1(G131), .B2(new_n226), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n224), .A2(new_n242), .B1(new_n200), .B2(new_n212), .ZN(new_n243));
  INV_X1    g057(.A(new_n237), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT28), .B1(new_n245), .B2(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(G237), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G210), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT27), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n188), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n241), .A2(new_n246), .A3(KEYINPUT70), .A4(new_n252), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT29), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n243), .B2(KEYINPUT64), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n229), .A2(new_n259), .A3(KEYINPUT30), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n244), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n253), .B1(new_n261), .B2(new_n238), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n247), .A2(new_n253), .ZN(new_n264));
  AOI21_X1  g078(.A(G902), .B1(new_n264), .B2(KEYINPUT29), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n187), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT30), .B1(new_n229), .B2(new_n259), .ZN(new_n267));
  AOI211_X1 g081(.A(KEYINPUT64), .B(new_n257), .C1(new_n213), .C2(new_n228), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n237), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n252), .A3(new_n239), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n252), .A4(new_n239), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(KEYINPUT31), .A3(new_n273), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n261), .A2(new_n253), .A3(new_n238), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n275), .A2(new_n276), .B1(new_n247), .B2(new_n253), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n187), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT32), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n274), .A2(new_n277), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(KEYINPUT69), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT32), .B1(new_n278), .B2(new_n187), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n266), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G475), .ZN(new_n290));
  INV_X1    g104(.A(G237), .ZN(new_n291));
  INV_X1    g105(.A(G953), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(G214), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n203), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n248), .A2(G143), .A3(G214), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n223), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT83), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n295), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G131), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n294), .A2(new_n301), .A3(new_n223), .A4(new_n295), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n297), .A2(new_n299), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT16), .ZN(new_n304));
  INV_X1    g118(.A(G125), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n307));
  OAI21_X1  g121(.A(G140), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT71), .B(G125), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n312), .A2(KEYINPUT16), .A3(G140), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n201), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n310), .B1(new_n312), .B2(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(new_n312), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n304), .A3(new_n309), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(G146), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n298), .A2(KEYINPUT17), .A3(G131), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n303), .A2(new_n314), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT18), .A2(G131), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n298), .B(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(G125), .B(G140), .Z(new_n324));
  OR2_X1    g138(.A1(new_n324), .A2(G146), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n315), .B2(new_n201), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G113), .B(G122), .ZN(new_n328));
  INV_X1    g142(.A(G104), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT85), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n321), .A2(new_n327), .A3(KEYINPUT86), .A4(new_n331), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n321), .A2(new_n327), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(new_n330), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n290), .B1(new_n338), .B2(new_n283), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n297), .A2(new_n302), .A3(new_n299), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT19), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n342));
  OAI22_X1  g156(.A1(new_n315), .A2(new_n341), .B1(new_n324), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n340), .B(new_n319), .C1(G146), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n330), .B1(new_n344), .B2(new_n327), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  NOR2_X1   g162(.A1(G475), .A2(G902), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n347), .A2(KEYINPUT87), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n334), .B2(new_n335), .ZN(new_n351));
  INV_X1    g165(.A(new_n349), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT87), .B1(new_n355), .B2(new_n348), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n339), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G116), .B(G122), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT88), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT89), .B1(new_n214), .B2(G143), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n203), .A3(G128), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(G128), .B2(new_n203), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(G134), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n362), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT13), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n367), .A2(new_n372), .B1(new_n214), .B2(G143), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT90), .B1(new_n367), .B2(new_n372), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n364), .A2(new_n366), .A3(new_n375), .A4(KEYINPUT13), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G134), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n377), .B2(G134), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n363), .B(new_n371), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n368), .B(new_n190), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n359), .A2(new_n360), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n359), .A2(KEYINPUT92), .A3(new_n360), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G116), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(G122), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n360), .B1(new_n391), .B2(KEYINPUT14), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n359), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n383), .B1(new_n384), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n389), .A2(new_n395), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n368), .B(G134), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT93), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT9), .B(G234), .ZN(new_n402));
  INV_X1    g216(.A(G217), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n402), .A2(new_n403), .A3(G953), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n382), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n382), .B2(new_n401), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n283), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G478), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT15), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n382), .A2(new_n401), .ZN(new_n412));
  INV_X1    g226(.A(new_n404), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(G902), .B1(new_n414), .B2(new_n405), .ZN(new_n415));
  INV_X1    g229(.A(new_n410), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G952), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G953), .ZN(new_n420));
  NAND2_X1  g234(.A1(G234), .A2(G237), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n421), .A2(G902), .A3(G953), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(G898), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n358), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G221), .B1(new_n402), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n221), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n220), .A2(new_n202), .A3(new_n204), .A4(KEYINPUT76), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n219), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT3), .B1(new_n329), .B2(G107), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT3), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n360), .A3(G104), .ZN(new_n437));
  INV_X1    g251(.A(G101), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n329), .A2(G107), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n435), .A2(new_n437), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n329), .A2(G107), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n360), .A2(G104), .ZN(new_n442));
  OAI21_X1  g256(.A(G101), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n434), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT10), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n200), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G101), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT4), .A3(new_n440), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n452), .A3(G101), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n212), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n446), .B1(new_n219), .B2(new_n221), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n444), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n447), .A2(new_n448), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n445), .A2(new_n446), .B1(new_n444), .B2(new_n455), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT77), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n448), .A4(new_n454), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n292), .A2(G227), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT75), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G140), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n440), .A2(new_n443), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n220), .A2(new_n204), .B1(new_n202), .B2(G128), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n431), .B2(new_n221), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n470), .B2(new_n433), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n444), .A2(new_n222), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n200), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(KEYINPUT12), .B(new_n200), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n462), .A2(new_n467), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n459), .A2(new_n454), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n200), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n467), .B1(new_n462), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n430), .B(new_n283), .C1(new_n478), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n466), .B1(new_n458), .B2(new_n461), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n480), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n458), .A2(new_n461), .B1(new_n476), .B2(new_n475), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n485), .B(G469), .C1(new_n467), .C2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n430), .A2(new_n283), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n429), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n211), .A2(new_n207), .ZN(new_n492));
  INV_X1    g306(.A(new_n206), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n317), .ZN(new_n494));
  INV_X1    g308(.A(new_n221), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n312), .B1(new_n495), .B2(new_n469), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G224), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(G953), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT79), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(KEYINPUT7), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n231), .A2(new_n232), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n232), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G119), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G116), .ZN(new_n507));
  OAI21_X1  g321(.A(G113), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n468), .B(new_n502), .C1(new_n505), .C2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G110), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT8), .ZN(new_n511));
  INV_X1    g325(.A(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n232), .A2(KEYINPUT5), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n512), .A2(new_n513), .B1(new_n231), .B2(new_n232), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n509), .B(new_n511), .C1(new_n514), .C2(new_n468), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n500), .A2(KEYINPUT7), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n494), .A2(new_n496), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT80), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT80), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n494), .A2(new_n496), .A3(new_n519), .A4(new_n516), .ZN(new_n520));
  AND4_X1   g334(.A1(new_n501), .A2(new_n515), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n237), .A2(new_n451), .A3(new_n453), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n444), .B(new_n502), .C1(new_n508), .C2(new_n505), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n510), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n523), .ZN(new_n526));
  INV_X1    g340(.A(new_n510), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n524), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT6), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n497), .B(new_n500), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G210), .B1(G237), .B2(G902), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n535), .B(KEYINPUT81), .Z(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n536), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n525), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G214), .B1(G237), .B2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT82), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(KEYINPUT82), .A3(new_n541), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n491), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n428), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT74), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(KEYINPUT25), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n506), .A2(G128), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n506), .A2(G128), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT24), .B(G110), .Z(new_n554));
  NAND3_X1  g368(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(new_n552), .C1(new_n550), .C2(KEYINPUT23), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n553), .A2(new_n554), .B1(G110), .B2(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n319), .A2(new_n325), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n554), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(G110), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n314), .B2(new_n319), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT72), .B1(new_n558), .B2(new_n562), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT22), .B(G137), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n292), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(KEYINPUT73), .Z(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n569), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n549), .B1(new_n573), .B2(G902), .ZN(new_n574));
  INV_X1    g388(.A(new_n549), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n571), .A2(new_n283), .A3(new_n572), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n403), .B1(G234), .B2(new_n283), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(G902), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n571), .A2(new_n572), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n289), .A2(new_n547), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n438), .ZN(G3));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n491), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n525), .A2(new_n533), .A3(new_n586), .A4(new_n538), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n541), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n534), .B2(new_n536), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(new_n539), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n278), .A2(new_n187), .ZN(new_n591));
  AOI211_X1 g405(.A(G472), .B(G902), .C1(new_n274), .C2(new_n277), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n585), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n339), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n350), .A2(new_n353), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(new_n356), .ZN(new_n597));
  INV_X1    g411(.A(new_n425), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n409), .A2(new_n283), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n415), .B2(new_n409), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT33), .B1(new_n406), .B2(new_n407), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n414), .A2(new_n405), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(G478), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n594), .A2(new_n597), .A3(new_n598), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT95), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n610));
  INV_X1    g424(.A(new_n353), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n351), .A2(KEYINPUT20), .A3(new_n352), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n353), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n339), .B1(new_n411), .B2(new_n417), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n598), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n594), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  INV_X1    g436(.A(new_n580), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n565), .A2(new_n566), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n570), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n579), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n428), .A2(new_n593), .A3(new_n546), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT97), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT37), .B(G110), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  NOR2_X1   g445(.A1(new_n289), .A2(new_n491), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n627), .A2(new_n590), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n422), .B1(new_n423), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n616), .A2(new_n617), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  NOR2_X1   g454(.A1(new_n286), .A2(new_n287), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n592), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n272), .A2(new_n273), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n253), .B1(new_n245), .B2(new_n238), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT99), .Z(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  OAI22_X1  g460(.A1(new_n641), .A2(new_n642), .B1(new_n187), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n597), .A2(new_n418), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n540), .B(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n541), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n627), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n647), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n656));
  INV_X1    g470(.A(new_n429), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n462), .A2(new_n477), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n658), .A2(new_n466), .B1(new_n484), .B2(new_n480), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n488), .B1(new_n659), .B2(G469), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n657), .B1(new_n660), .B2(new_n482), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n635), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n655), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n203), .ZN(G45));
  NAND3_X1  g480(.A1(new_n597), .A2(new_n605), .A3(new_n636), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n633), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n632), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT101), .B(G146), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G48));
  INV_X1    g485(.A(new_n266), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n641), .B2(new_n642), .ZN(new_n673));
  INV_X1    g487(.A(new_n582), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n478), .A2(new_n481), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n590), .A2(new_n429), .A3(new_n482), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n597), .A2(new_n605), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n677), .A2(new_n678), .A3(new_n425), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n673), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  NOR2_X1   g496(.A1(new_n618), .A2(new_n582), .ZN(new_n683));
  INV_X1    g497(.A(new_n677), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n673), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NOR2_X1   g500(.A1(new_n626), .A2(new_n623), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n578), .B2(new_n577), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n427), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n673), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT102), .B(G119), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G21));
  NAND2_X1  g506(.A1(new_n282), .A2(new_n283), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G472), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(KEYINPUT103), .A3(new_n279), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n278), .A2(KEYINPUT103), .A3(new_n187), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n597), .A2(new_n418), .A3(new_n598), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n677), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n700), .A3(new_n674), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  AOI21_X1  g516(.A(new_n688), .B1(new_n695), .B2(new_n697), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n667), .A2(new_n677), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n703), .A2(KEYINPUT104), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n661), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n537), .A2(new_n541), .A3(new_n539), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n661), .B2(new_n711), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n673), .A2(new_n674), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n597), .A2(new_n605), .A3(new_n636), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n714), .B1(new_n491), .B2(KEYINPUT105), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n712), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n672), .B1(new_n592), .B2(KEYINPUT32), .ZN(new_n723));
  INV_X1    g537(.A(new_n284), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n674), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT42), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n223), .ZN(G33));
  INV_X1    g542(.A(new_n637), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n673), .A2(new_n674), .A3(new_n729), .A4(new_n717), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  AOI21_X1  g545(.A(KEYINPUT43), .B1(new_n358), .B2(new_n605), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n597), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n595), .B(KEYINPUT108), .C1(new_n596), .C2(new_n356), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n605), .A2(KEYINPUT43), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT109), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n737), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n734), .A4(new_n735), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n732), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n593), .A3(new_n688), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(KEYINPUT44), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT110), .Z(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n484), .A2(new_n480), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n486), .A2(new_n467), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n658), .A2(new_n466), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT45), .A3(new_n485), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n753), .A3(G469), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT106), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n751), .A2(new_n753), .A3(new_n756), .A4(G469), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n747), .B(new_n488), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n746), .B1(new_n758), .B2(new_n483), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n752), .A2(new_n485), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n430), .B1(new_n760), .B2(new_n748), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n756), .B1(new_n761), .B2(new_n753), .ZN(new_n762));
  INV_X1    g576(.A(new_n757), .ZN(new_n763));
  OAI211_X1 g577(.A(KEYINPUT46), .B(new_n489), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(KEYINPUT107), .A3(new_n482), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n763), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n747), .B1(new_n766), .B2(new_n488), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n759), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n429), .A3(new_n662), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n714), .B(new_n769), .C1(KEYINPUT44), .C2(new_n743), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n745), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(KEYINPUT111), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n765), .A2(new_n767), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT107), .B1(new_n764), .B2(new_n482), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n429), .B(new_n775), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n768), .B2(new_n429), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n673), .A2(new_n674), .A3(new_n667), .A4(new_n714), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  AND2_X1   g599(.A1(new_n676), .A2(new_n482), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n429), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n715), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n674), .A2(new_n422), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n597), .A2(new_n605), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n647), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n422), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n742), .A2(new_n793), .A3(new_n789), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n792), .B1(new_n794), .B2(new_n703), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n742), .A2(new_n793), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n582), .B1(new_n695), .B2(new_n697), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n788), .A2(new_n652), .A3(new_n651), .ZN(new_n798));
  NOR2_X1   g612(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n738), .A2(new_n741), .ZN(new_n801));
  INV_X1    g615(.A(new_n732), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n422), .A3(new_n797), .A4(new_n798), .ZN(new_n804));
  XOR2_X1   g618(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n795), .A2(new_n800), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n786), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n429), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n429), .B1(new_n776), .B2(new_n777), .ZN(new_n810));
  INV_X1    g624(.A(new_n780), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n809), .B1(new_n812), .B2(new_n778), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n796), .A2(new_n797), .A3(new_n715), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT115), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n779), .A2(new_n781), .B1(new_n429), .B2(new_n808), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  INV_X1    g631(.A(new_n814), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n807), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n795), .A2(new_n806), .A3(new_n800), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n795), .A2(new_n806), .A3(new_n825), .A4(new_n800), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n821), .B1(new_n816), .B2(new_n818), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n796), .A2(new_n684), .A3(new_n797), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n647), .A2(new_n789), .A3(new_n790), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n829), .B(new_n420), .C1(new_n678), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n725), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n794), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT48), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT48), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n822), .A2(new_n828), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n719), .A2(new_n730), .A3(new_n726), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n680), .A2(new_n685), .A3(new_n690), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n418), .A2(new_n339), .A3(new_n635), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n616), .A2(new_n627), .A3(new_n715), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n673), .A2(new_n661), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT103), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n591), .A2(new_n592), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n627), .B1(new_n846), .B2(new_n696), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n844), .B1(new_n847), .B2(new_n722), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n703), .A2(KEYINPUT112), .A3(new_n717), .A4(new_n720), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n843), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n617), .B1(new_n356), .B2(new_n596), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n678), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n425), .B1(new_n544), .B2(new_n545), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n585), .A3(new_n853), .A4(new_n593), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n701), .A2(new_n628), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n583), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n839), .A2(new_n840), .A3(new_n850), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n673), .B(new_n661), .C1(new_n638), .C2(new_n668), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n649), .A2(new_n590), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n627), .A2(new_n491), .A3(new_n635), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n647), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n708), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT104), .B1(new_n703), .B2(new_n704), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n858), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n709), .A2(KEYINPUT52), .A3(new_n858), .A4(new_n861), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT53), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n839), .A2(new_n840), .A3(new_n850), .A4(new_n856), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n866), .A2(new_n867), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n873), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n870), .B2(new_n871), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n877), .A2(KEYINPUT114), .B1(new_n868), .B2(KEYINPUT53), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n868), .B2(new_n876), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n822), .A2(new_n883), .A3(new_n828), .A4(new_n836), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n838), .A2(new_n875), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n882), .A2(new_n875), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n887), .A2(new_n888), .A3(new_n838), .A4(new_n884), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n419), .A2(new_n292), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n786), .B(KEYINPUT49), .Z(new_n892));
  NOR2_X1   g706(.A1(new_n657), .A2(new_n652), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n674), .A2(new_n605), .A3(new_n651), .A4(new_n893), .ZN(new_n894));
  OR4_X1    g708(.A1(new_n647), .A2(new_n892), .A3(new_n736), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(G75));
  XOR2_X1   g710(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n897));
  NAND3_X1  g711(.A1(new_n872), .A2(KEYINPUT114), .A3(new_n873), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT53), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n877), .A2(KEYINPUT114), .ZN(new_n901));
  OAI211_X1 g715(.A(G902), .B(new_n536), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n529), .A2(new_n531), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n532), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n902), .B2(new_n903), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n897), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n903), .ZN(new_n909));
  INV_X1    g723(.A(new_n905), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n897), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n292), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n908), .A2(new_n914), .A3(new_n916), .ZN(G51));
  XNOR2_X1  g731(.A(new_n488), .B(KEYINPUT57), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n879), .B1(new_n878), .B2(new_n881), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n882), .B1(new_n919), .B2(KEYINPUT121), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n921), .B(new_n879), .C1(new_n878), .C2(new_n881), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n675), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n900), .A2(new_n901), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n283), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n766), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n915), .B1(new_n925), .B2(new_n928), .ZN(G54));
  NAND3_X1  g743(.A1(new_n927), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n351), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n916), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n351), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G60));
  XNOR2_X1  g748(.A(new_n599), .B(KEYINPUT59), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n882), .B2(new_n875), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n601), .A2(new_n603), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT122), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n916), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n920), .A2(new_n922), .ZN(new_n940));
  INV_X1    g754(.A(new_n935), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n573), .B1(new_n926), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n945), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n626), .B(KEYINPUT123), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n947), .B(new_n948), .C1(new_n900), .C2(new_n901), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(new_n916), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n424), .B2(new_n498), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n840), .A2(new_n856), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n904), .B1(G898), .B2(new_n292), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  NAND2_X1  g772(.A1(new_n709), .A2(new_n858), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n665), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT62), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n663), .A2(new_n714), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n673), .A2(new_n674), .A3(new_n852), .A4(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n961), .A2(new_n771), .A3(new_n784), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n292), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n267), .A2(new_n268), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(new_n343), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n292), .A2(G900), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n839), .B(KEYINPUT125), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n832), .A2(new_n859), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n769), .A2(new_n972), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n959), .B(new_n973), .C1(new_n782), .C2(new_n783), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n771), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n975), .B2(new_n292), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n968), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n292), .B1(G227), .B2(G900), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n978), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n968), .B(new_n980), .C1(new_n967), .C2(new_n976), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(G72));
  XNOR2_X1  g796(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n964), .B2(new_n954), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n261), .A2(new_n238), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n252), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n643), .A2(new_n262), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n985), .B(new_n990), .C1(new_n869), .C2(new_n874), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n985), .B1(new_n975), .B2(new_n954), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n988), .A2(new_n252), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n916), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n995), .A2(KEYINPUT127), .A3(new_n916), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(G57));
endmodule


