//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G227gat), .ZN(new_n204));
  INV_X1    g003(.A(G233gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(G120gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT67), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G127gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(G120gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(new_n208), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n214), .B(new_n218), .C1(new_n223), .C2(new_n209), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(KEYINPUT24), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  OR3_X1    g030(.A1(new_n231), .A2(G169gat), .A3(G176gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n229), .A2(KEYINPUT24), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n230), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT64), .B(G176gat), .ZN(new_n240));
  INV_X1    g039(.A(G169gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(KEYINPUT23), .A3(new_n241), .ZN(new_n242));
  AND4_X1   g041(.A1(new_n239), .A2(new_n242), .A3(new_n236), .A4(new_n234), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n230), .A2(new_n233), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n238), .A2(KEYINPUT25), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT27), .B(G183gat), .Z(new_n246));
  OAI21_X1  g045(.A(KEYINPUT28), .B1(new_n246), .B2(G190gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n248), .A2(new_n226), .A3(KEYINPUT27), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT27), .B1(new_n248), .B2(new_n226), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n227), .A4(new_n251), .ZN(new_n252));
  OR3_X1    g051(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n236), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n247), .A2(new_n252), .A3(new_n229), .A4(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n225), .B1(new_n245), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n242), .A2(new_n239), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(new_n236), .A3(new_n234), .A4(new_n244), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT25), .B1(new_n235), .B2(new_n237), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n221), .A2(new_n224), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n206), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n225), .A3(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n262), .ZN(new_n266));
  INV_X1    g065(.A(new_n206), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n268), .A3(KEYINPUT32), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT32), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n265), .A2(new_n266), .A3(new_n270), .A4(new_n267), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n203), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n264), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n274), .A2(KEYINPUT33), .ZN(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G71gat), .ZN(new_n277));
  INV_X1    g076(.A(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n269), .A2(new_n203), .A3(new_n271), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n273), .A2(new_n275), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n279), .ZN(new_n282));
  INV_X1    g081(.A(new_n280), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n272), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT36), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G1gat), .B(G29gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT78), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G85gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G155gat), .B(G162gat), .Z(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(KEYINPUT2), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(G155gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G162gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n299), .B1(new_n303), .B2(KEYINPUT2), .ZN(new_n304));
  INV_X1    g103(.A(G148gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT72), .B1(new_n305), .B2(G141gat), .ZN(new_n306));
  OR3_X1    g105(.A1(new_n305), .A2(KEYINPUT72), .A3(G141gat), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT73), .B(G148gat), .Z(new_n308));
  INV_X1    g107(.A(G141gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n306), .B(new_n307), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(KEYINPUT75), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT75), .B1(new_n304), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n301), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n304), .A2(new_n310), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n311), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n301), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(new_n321), .A3(new_n262), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT5), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT4), .B1(new_n314), .B2(new_n262), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n319), .A2(new_n225), .A3(new_n330), .A4(new_n301), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n332), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT80), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n328), .A3(new_n339), .ZN(new_n340));
  AOI211_X1 g139(.A(new_n323), .B(new_n327), .C1(new_n336), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n328), .A2(new_n331), .A3(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT76), .B(KEYINPUT4), .C1(new_n314), .C2(new_n262), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n343), .A2(new_n324), .A3(new_n344), .A4(new_n322), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n314), .A2(new_n262), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n225), .B1(new_n319), .B2(new_n301), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n325), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(KEYINPUT5), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n298), .B1(new_n341), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n334), .A2(new_n335), .A3(new_n329), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n328), .B1(new_n338), .B2(new_n339), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n322), .B(new_n326), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(new_n297), .A3(new_n349), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n297), .B1(new_n355), .B2(new_n349), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT6), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT84), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT84), .B1(new_n358), .B2(KEYINPUT6), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n261), .A2(G226gat), .A3(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n261), .A2(new_n365), .B1(G226gat), .B2(G233gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G197gat), .B(G204gat), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  INV_X1    g167(.A(G218gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(KEYINPUT22), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G211gat), .B(G218gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  OR3_X1    g172(.A1(new_n364), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n364), .B2(new_n366), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT37), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  INV_X1    g178(.A(G36gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT71), .B(G8gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  AND2_X1   g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT38), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n374), .A2(new_n375), .ZN(new_n388));
  INV_X1    g187(.A(new_n383), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n378), .A2(new_n383), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(KEYINPUT38), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n361), .A2(new_n363), .A3(new_n387), .A4(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  INV_X1    g194(.A(G50gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT83), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n320), .B1(new_n373), .B2(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n314), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n403), .A2(new_n404), .B1(G228gat), .B2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n373), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n321), .B2(new_n365), .ZN(new_n407));
  INV_X1    g206(.A(new_n403), .ZN(new_n408));
  OR3_X1    g207(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n401), .B(new_n412), .C1(new_n414), .C2(new_n400), .ZN(new_n415));
  INV_X1    g214(.A(new_n412), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT83), .B(new_n400), .C1(new_n416), .C2(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n376), .B2(new_n383), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n390), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n388), .A2(new_n420), .A3(new_n389), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OR3_X1    g223(.A1(new_n346), .A2(new_n347), .A3(new_n325), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n323), .B1(new_n336), .B2(new_n340), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT39), .B(new_n425), .C1(new_n426), .C2(new_n324), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n322), .B1(new_n353), .B2(new_n354), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT39), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n325), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n430), .A3(new_n297), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT40), .ZN(new_n432));
  AOI211_X1 g231(.A(new_n358), .B(new_n424), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT40), .A4(new_n297), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n419), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n291), .B1(new_n394), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n360), .ZN(new_n437));
  INV_X1    g236(.A(new_n424), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n419), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n285), .B1(new_n415), .B2(new_n417), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n360), .A2(new_n424), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n445), .B1(new_n357), .B2(new_n359), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n440), .B(new_n444), .C1(new_n446), .C2(new_n362), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n436), .A2(new_n439), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449));
  NAND2_X1  g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n449), .B1(new_n450), .B2(KEYINPUT94), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT94), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(G85gat), .A3(G92gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT7), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n457), .A2(KEYINPUT8), .ZN(new_n458));
  NOR2_X1   g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT95), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(KEYINPUT8), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT95), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n462), .C1(G85gat), .C2(G92gat), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n456), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n450), .A2(KEYINPUT93), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G99gat), .B(G106gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(new_n467), .A3(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G57gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(G64gat), .ZN(new_n473));
  INV_X1    g272(.A(G64gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(G57gat), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT90), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G71gat), .A2(G78gat), .ZN(new_n477));
  OR2_X1    g276(.A1(G71gat), .A2(G78gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT9), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(G57gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(G64gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT91), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n476), .A2(new_n487), .A3(new_n480), .A4(new_n484), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n478), .A2(new_n477), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n481), .A2(new_n482), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(KEYINPUT9), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT92), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n495));
  AOI211_X1 g294(.A(new_n495), .B(new_n492), .C1(new_n486), .C2(new_n488), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n471), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n464), .A2(new_n467), .A3(new_n465), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n467), .B1(new_n464), .B2(new_n465), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n489), .A2(new_n493), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G230gat), .A2(G233gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT100), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT101), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n505), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT99), .B(KEYINPUT10), .Z(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n497), .B2(new_n502), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n500), .B(KEYINPUT10), .C1(new_n494), .C2(new_n496), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n507), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n508), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G176gat), .B(G204gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n519), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n508), .A2(new_n521), .A3(new_n514), .A4(new_n515), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n396), .A2(G43gat), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT15), .B1(new_n396), .B2(G43gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n396), .A2(G43gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT88), .B(G43gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(G50gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n380), .A3(KEYINPUT14), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT87), .B(G36gat), .Z(new_n536));
  OAI211_X1 g335(.A(new_n533), .B(new_n535), .C1(new_n536), .C2(new_n534), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n524), .B2(new_n525), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT16), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(G1gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G1gat), .B2(new_n543), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n546), .B(G8gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n547), .ZN(new_n549));
  INV_X1    g348(.A(new_n540), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT89), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n548), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n555), .A2(KEYINPUT18), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n547), .A2(new_n540), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n553), .B(KEYINPUT13), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(KEYINPUT18), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G169gat), .B(G197gat), .Z(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT12), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n556), .A2(new_n570), .A3(new_n561), .A4(new_n560), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n448), .A2(new_n523), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n542), .A2(new_n471), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n550), .A2(new_n500), .ZN(new_n576));
  NAND3_X1  g375(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT96), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT97), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n586), .A3(new_n583), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(KEYINPUT97), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n501), .A2(new_n495), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n489), .A2(KEYINPUT92), .A3(new_n493), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(G183gat), .B1(new_n600), .B2(new_n549), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT21), .B1(new_n494), .B2(new_n496), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n226), .A3(new_n547), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT21), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n601), .B2(new_n603), .ZN(new_n608));
  INV_X1    g407(.A(G231gat), .ZN(new_n609));
  OAI22_X1  g408(.A1(new_n607), .A2(new_n608), .B1(new_n609), .B2(new_n205), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n601), .A2(new_n603), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n604), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n612), .A2(new_n606), .A3(G231gat), .A4(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G211gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n610), .B2(new_n613), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n596), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n595), .A3(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n594), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT98), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n594), .A2(new_n622), .A3(new_n620), .A4(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n574), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n437), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g430(.A(G8gat), .B1(new_n628), .B2(new_n424), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT42), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G8gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n629), .A2(new_n438), .A3(new_n635), .ZN(new_n636));
  MUX2_X1   g435(.A(KEYINPUT42), .B(new_n633), .S(new_n636), .Z(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n628), .B2(new_n285), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT103), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n291), .B(KEYINPUT104), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n628), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(G1326gat));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n418), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT43), .B(G22gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  NOR2_X1   g445(.A1(new_n448), .A2(new_n594), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n622), .A2(new_n620), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n649), .A2(new_n523), .A3(new_n573), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n534), .A3(new_n437), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT45), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT44), .B1(new_n448), .B2(new_n594), .ZN(new_n655));
  INV_X1    g454(.A(new_n291), .ZN(new_n656));
  NOR4_X1   g455(.A1(new_n446), .A2(new_n362), .A3(new_n386), .A4(new_n392), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n424), .B1(new_n431), .B2(new_n432), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n351), .A3(new_n434), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n418), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n439), .B(new_n656), .C1(new_n657), .C2(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n442), .A2(new_n447), .A3(KEYINPUT106), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT106), .B1(new_n442), .B2(new_n447), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  INV_X1    g464(.A(new_n594), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n655), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n650), .B(KEYINPUT105), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n360), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n671), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT107), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n652), .A2(new_n536), .A3(new_n438), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(KEYINPUT107), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n536), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n670), .B2(new_n424), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n651), .A2(new_n678), .A3(new_n424), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(KEYINPUT107), .A3(new_n673), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT108), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n677), .A2(new_n684), .A3(new_n679), .A4(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1329gat));
  INV_X1    g485(.A(new_n285), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n652), .A2(new_n528), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n670), .A2(new_n641), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(new_n528), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n670), .A2(new_n656), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n693), .B2(new_n528), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n691), .B2(new_n694), .ZN(G1330gat));
  OAI21_X1  g494(.A(G50gat), .B1(new_n670), .B2(new_n418), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT48), .B1(new_n696), .B2(KEYINPUT110), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n418), .B1(new_n651), .B2(KEYINPUT109), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n698), .B(new_n396), .C1(KEYINPUT109), .C2(new_n651), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n696), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n697), .B(new_n700), .ZN(G1331gat));
  NAND4_X1  g500(.A1(new_n664), .A2(new_n627), .A3(new_n523), .A4(new_n573), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n360), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(new_n472), .ZN(G1332gat));
  NAND2_X1  g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n702), .A2(new_n706), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n438), .B(new_n705), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT112), .ZN(new_n711));
  INV_X1    g510(.A(new_n702), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n707), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n438), .A4(new_n705), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n711), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n711), .B2(new_n716), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(G1333gat));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n641), .B1(new_n713), .B2(new_n707), .ZN(new_n722));
  INV_X1    g521(.A(G71gat), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n712), .A2(new_n723), .A3(new_n687), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n721), .B(new_n725), .C1(new_n722), .C2(new_n723), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n419), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n649), .A2(new_n572), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n668), .A2(new_n523), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n360), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n735));
  INV_X1    g534(.A(new_n663), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n442), .A2(new_n447), .A3(KEYINPUT106), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n594), .B1(new_n738), .B2(new_n661), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(new_n732), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n735), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AND4_X1   g542(.A1(new_n666), .A2(new_n664), .A3(new_n732), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n523), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n360), .A2(new_n746), .A3(G85gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT114), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n734), .B1(new_n745), .B2(new_n748), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n733), .B2(new_n424), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n746), .A2(G92gat), .A3(new_n424), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT115), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n745), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n733), .B2(new_n641), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n523), .B1(new_n740), .B2(new_n744), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n687), .A2(new_n278), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(G1338gat));
  NAND4_X1  g557(.A1(new_n668), .A2(new_n419), .A3(new_n523), .A4(new_n732), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G106gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n418), .A2(G106gat), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n523), .B(new_n761), .C1(new_n740), .C2(new_n744), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n763));
  AND3_X1   g562(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n760), .B2(new_n762), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT117), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(G1339gat));
  AOI21_X1  g570(.A(new_n554), .B1(new_n548), .B2(new_n551), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n558), .A2(new_n559), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n567), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT119), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(KEYINPUT119), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n571), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n746), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n505), .B(new_n512), .C1(new_n503), .C2(new_n510), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(KEYINPUT54), .A3(new_n514), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n781), .B(new_n509), .C1(new_n511), .C2(new_n513), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n782), .A2(new_n783), .A3(new_n519), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n782), .B2(new_n519), .ZN(new_n785));
  OAI211_X1 g584(.A(KEYINPUT55), .B(new_n780), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n572), .A2(new_n522), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n666), .B1(new_n778), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n522), .A3(new_n786), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n594), .A2(new_n792), .A3(new_n777), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n648), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n624), .A2(new_n626), .A3(new_n746), .A4(new_n573), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n419), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT120), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n360), .A2(new_n438), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n687), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n573), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n794), .A2(new_n795), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n440), .ZN(new_n802));
  INV_X1    g601(.A(new_n798), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n208), .A3(new_n572), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n805), .ZN(G1340gat));
  OAI21_X1  g605(.A(G120gat), .B1(new_n799), .B2(new_n746), .ZN(new_n807));
  INV_X1    g606(.A(new_n222), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n808), .A3(new_n523), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1341gat));
  NOR3_X1   g609(.A1(new_n799), .A2(new_n216), .A3(new_n648), .ZN(new_n811));
  AOI21_X1  g610(.A(G127gat), .B1(new_n804), .B2(new_n649), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(G1342gat));
  OAI21_X1  g612(.A(G134gat), .B1(new_n799), .B2(new_n594), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n802), .A2(G134gat), .A3(new_n594), .A4(new_n803), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT56), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1343gat));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n792), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n789), .A2(KEYINPUT121), .A3(new_n522), .A4(new_n786), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n572), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n778), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(KEYINPUT122), .A3(new_n778), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n594), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n793), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n649), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n795), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n419), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT57), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n418), .B1(new_n794), .B2(new_n795), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n803), .A2(new_n291), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n831), .A2(new_n572), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G141gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT123), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n832), .A2(new_n641), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n803), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n309), .A3(new_n572), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n842), .A3(KEYINPUT58), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n837), .B(new_n841), .C1(KEYINPUT123), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1344gat));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n418), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n795), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n828), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(new_n523), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n847), .B1(new_n853), .B2(new_n835), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n746), .A2(new_n308), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n854), .A2(G148gat), .B1(new_n840), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n831), .A2(new_n834), .A3(new_n835), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n523), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n308), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n859), .B2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g659(.A(new_n302), .B1(new_n840), .B2(new_n649), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n649), .A2(new_n302), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n857), .B2(new_n862), .ZN(G1346gat));
  AOI21_X1  g662(.A(G162gat), .B1(new_n840), .B2(new_n666), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n666), .A2(G162gat), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n857), .B2(new_n865), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n437), .A2(new_n424), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT125), .Z(new_n868));
  NAND3_X1  g667(.A1(new_n797), .A2(new_n687), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869), .B2(new_n573), .ZN(new_n870));
  INV_X1    g669(.A(new_n867), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n802), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n241), .A3(new_n572), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(G1348gat));
  NOR3_X1   g673(.A1(new_n869), .A2(new_n240), .A3(new_n746), .ZN(new_n875));
  AOI21_X1  g674(.A(G176gat), .B1(new_n872), .B2(new_n523), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(G1349gat));
  OAI21_X1  g676(.A(G183gat), .B1(new_n869), .B2(new_n648), .ZN(new_n878));
  INV_X1    g677(.A(new_n246), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n872), .A2(new_n649), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n872), .A2(new_n227), .A3(new_n666), .ZN(new_n883));
  OAI21_X1  g682(.A(G190gat), .B1(new_n869), .B2(new_n594), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(KEYINPUT61), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n886), .B(G190gat), .C1(new_n869), .C2(new_n594), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n883), .B1(new_n885), .B2(new_n888), .ZN(G1351gat));
  AND2_X1   g688(.A1(new_n868), .A2(new_n641), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n851), .A2(new_n852), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G197gat), .B1(new_n891), .B2(new_n573), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n839), .A2(new_n871), .ZN(new_n893));
  INV_X1    g692(.A(G197gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n572), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1352gat));
  INV_X1    g695(.A(G204gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n897), .A3(new_n523), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT62), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n853), .B2(new_n890), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n899), .A2(new_n900), .ZN(G1353gat));
  NAND4_X1  g700(.A1(new_n851), .A2(new_n649), .A3(new_n852), .A4(new_n890), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G211gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT63), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n893), .A2(new_n368), .A3(new_n649), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT126), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n893), .A2(new_n907), .A3(new_n368), .A4(new_n649), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n902), .A2(new_n910), .A3(G211gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT127), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n904), .A2(new_n909), .A3(new_n914), .A4(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n891), .B2(new_n594), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n369), .A3(new_n666), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1355gat));
endmodule


