//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  INV_X1    g001(.A(G101), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT3), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT74), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(KEYINPUT74), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n189), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n188), .B1(new_n195), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT4), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G116), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT2), .B(G113), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n208), .ZN(new_n210));
  XNOR2_X1  g024(.A(G116), .B(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n201), .A2(new_n202), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n193), .A2(KEYINPUT3), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n194), .B1(new_n192), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n191), .A2(G107), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n199), .B2(new_n197), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT75), .B(G101), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n195), .A2(new_n219), .A3(new_n200), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n188), .B1(new_n216), .B2(new_n199), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n215), .A2(new_n217), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(new_n219), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n207), .A2(new_n208), .ZN(new_n225));
  INV_X1    g039(.A(G113), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n227));
  INV_X1    g041(.A(new_n204), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n211), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n225), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n213), .A2(new_n221), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G110), .B(G122), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT81), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT6), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n233), .B2(new_n234), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n218), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n212), .A2(new_n209), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n202), .B(G101), .C1(new_n215), .C2(new_n217), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n231), .B(G113), .C1(new_n204), .C2(new_n230), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n212), .ZN(new_n243));
  INV_X1    g057(.A(new_n222), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n220), .A2(new_n244), .ZN(new_n245));
  OAI22_X1  g059(.A1(new_n238), .A2(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT81), .ZN(new_n247));
  INV_X1    g061(.A(new_n234), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n235), .A2(new_n237), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT0), .B(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n255), .A2(new_n262), .A3(G128), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n252), .B(new_n254), .C1(KEYINPUT1), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n268), .B(new_n270), .Z(new_n271));
  NAND3_X1  g085(.A1(new_n246), .A2(new_n236), .A3(new_n248), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT82), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n246), .A2(new_n274), .A3(new_n236), .A4(new_n248), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n250), .A2(new_n271), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n234), .B(KEYINPUT8), .Z(new_n278));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n229), .B1(new_n279), .B2(new_n207), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n224), .A2(new_n212), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n243), .A2(new_n245), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n270), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n268), .A2(new_n285), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n284), .B(new_n270), .C1(new_n261), .C2(new_n267), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n233), .A2(new_n234), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n276), .A2(new_n277), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n277), .B1(new_n276), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(KEYINPUT83), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n294), .B(new_n277), .C1(new_n276), .C2(new_n290), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G214), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n187), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT84), .B(new_n297), .C1(new_n293), .C2(new_n295), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G131), .ZN(new_n302));
  INV_X1    g116(.A(G137), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT11), .B1(new_n303), .B2(G134), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(G134), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(KEYINPUT64), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT64), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G137), .ZN(new_n309));
  AND2_X1   g123(.A1(KEYINPUT11), .A2(G134), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n302), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT64), .B(G137), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n314), .A2(new_n310), .B1(new_n304), .B2(new_n305), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT65), .B(G131), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n312), .A2(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT66), .B1(new_n315), .B2(new_n302), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n317), .A2(new_n318), .B1(new_n257), .B2(new_n259), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n263), .A2(new_n266), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n316), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n305), .B1(new_n314), .B2(G134), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n319), .A2(new_n324), .A3(new_n239), .ZN(new_n325));
  INV_X1    g139(.A(new_n239), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n306), .A2(new_n311), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n313), .A3(G131), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n321), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n312), .A2(new_n313), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n260), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT28), .B1(new_n325), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT68), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n325), .B2(KEYINPUT28), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n326), .A3(new_n332), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(KEYINPUT68), .A3(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n334), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(G237), .A2(G953), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G210), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT27), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G101), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(KEYINPUT69), .A3(KEYINPUT29), .A4(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n334), .A2(new_n336), .A3(new_n345), .A4(new_n339), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G902), .ZN(new_n351));
  INV_X1    g165(.A(new_n345), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT30), .B1(new_n319), .B2(new_n324), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n331), .A2(new_n354), .A3(new_n332), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n326), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(new_n325), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n348), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n346), .A2(new_n350), .A3(new_n351), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G472), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT30), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n354), .B1(new_n331), .B2(new_n332), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n239), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n345), .A4(new_n337), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT67), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n353), .A2(new_n355), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n325), .B1(new_n369), .B2(new_n239), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT67), .A3(new_n365), .A4(new_n345), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n334), .A2(new_n336), .A3(new_n339), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n345), .A3(new_n337), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n352), .A2(new_n373), .B1(new_n374), .B2(KEYINPUT31), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G472), .ZN(new_n377));
  AND4_X1   g191(.A1(new_n361), .A2(new_n376), .A3(new_n377), .A4(new_n351), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n372), .B2(new_n375), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n361), .B1(new_n379), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n360), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n191), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n341), .A2(G143), .A3(G214), .ZN(new_n385));
  AOI21_X1  g199(.A(G143), .B1(new_n341), .B2(G214), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n384), .B1(new_n387), .B2(new_n316), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n316), .ZN(new_n389));
  INV_X1    g203(.A(new_n316), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n390), .B(KEYINPUT85), .C1(new_n385), .C2(new_n386), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G140), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n264), .A2(G140), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT16), .ZN(new_n396));
  OR3_X1    g210(.A1(new_n264), .A2(KEYINPUT16), .A3(G140), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G146), .ZN(new_n398));
  XNOR2_X1  g212(.A(G125), .B(G140), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT19), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n251), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n387), .B1(new_n403), .B2(new_n302), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT18), .B(G131), .C1(new_n385), .C2(new_n386), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n399), .B(new_n251), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n383), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n407), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n397), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n251), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n398), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n388), .A2(new_n391), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(KEYINPUT17), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n388), .A2(new_n389), .A3(new_n415), .A4(new_n391), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n409), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n383), .B(KEYINPUT86), .Z(new_n418));
  AOI21_X1  g232(.A(new_n408), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(new_n416), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n424), .A2(new_n407), .A3(new_n418), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n423), .B(new_n420), .C1(new_n425), .C2(new_n408), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n253), .A2(G128), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n265), .A2(G143), .ZN(new_n429));
  INV_X1    g243(.A(G134), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n205), .A2(G122), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G107), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n189), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n432), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n265), .A2(G143), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n428), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n439), .B1(new_n430), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n205), .A3(G122), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT14), .B1(new_n433), .B2(G116), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n433), .A2(G116), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n449), .A2(new_n450), .A3(G107), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n449), .B2(G107), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n430), .B1(new_n428), .B2(new_n429), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT87), .B1(new_n432), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n253), .A2(G128), .ZN(new_n456));
  OAI21_X1  g270(.A(G134), .B1(new_n440), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n431), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n438), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n444), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT9), .B(G234), .ZN(new_n462));
  INV_X1    g276(.A(G217), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n462), .A2(new_n463), .A3(G953), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n444), .B(new_n464), .C1(new_n453), .C2(new_n460), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n351), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n469), .A2(new_n471), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(G234), .A2(G237), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(G952), .A3(new_n269), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT21), .B(G898), .Z(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(G902), .A3(G953), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n479), .B(KEYINPUT89), .Z(new_n480));
  NOR2_X1   g294(.A1(new_n417), .A2(new_n383), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n351), .B1(new_n425), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G475), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n427), .A2(new_n474), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n422), .A2(new_n426), .B1(new_n482), .B2(G475), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(KEYINPUT90), .A3(new_n480), .A4(new_n474), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G221), .B1(new_n462), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G469), .ZN(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G140), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n269), .A2(G227), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n493), .B(new_n494), .Z(new_n495));
  NAND2_X1  g309(.A1(new_n240), .A2(new_n260), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT10), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n220), .A2(new_n266), .A3(new_n263), .A4(new_n244), .ZN(new_n498));
  OAI22_X1  g312(.A1(new_n238), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n498), .B2(new_n497), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n317), .A2(new_n318), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT78), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n498), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT10), .ZN(new_n509));
  INV_X1    g323(.A(new_n496), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n221), .ZN(new_n511));
  INV_X1    g325(.A(new_n501), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n509), .B(new_n511), .C1(new_n512), .C2(new_n502), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT78), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n499), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n517), .B(new_n506), .C1(new_n512), .C2(new_n502), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n495), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n495), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT12), .B1(new_n505), .B2(KEYINPUT77), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n220), .A2(new_n244), .B1(new_n266), .B2(new_n263), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n505), .B1(new_n508), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI221_X1 g338(.A(new_n505), .B1(KEYINPUT77), .B2(KEYINPUT12), .C1(new_n508), .C2(new_n522), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT79), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(KEYINPUT79), .A3(new_n525), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n520), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n492), .B(new_n351), .C1(new_n519), .C2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n495), .B1(new_n518), .B2(new_n526), .ZN(new_n532));
  INV_X1    g346(.A(new_n495), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n504), .B2(new_n506), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n516), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G469), .B1(new_n535), .B2(G902), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n491), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n489), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n463), .B1(G234), .B2(new_n351), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n265), .A2(G119), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n203), .A2(G128), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT70), .B1(new_n203), .B2(G128), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT23), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n540), .A2(KEYINPUT70), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n548), .A3(new_n541), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n549), .B2(G110), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n412), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G110), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n546), .A2(new_n548), .A3(new_n552), .A4(new_n541), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n542), .A2(new_n543), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n399), .A2(new_n251), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n398), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT22), .B(G137), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n562), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n558), .B1(new_n551), .B2(new_n557), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n551), .A2(new_n557), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n562), .B(new_n563), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n569), .A2(KEYINPUT72), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n351), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT25), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT25), .B(new_n351), .C1(new_n568), .C2(new_n571), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT73), .ZN(new_n577));
  INV_X1    g391(.A(new_n567), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n565), .A3(new_n559), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n566), .A2(new_n567), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT25), .B1(new_n581), .B2(new_n351), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n539), .B(new_n575), .C1(new_n577), .C2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n539), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n301), .A2(new_n381), .A3(new_n538), .A4(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(new_n219), .Z(G3));
  NAND2_X1  g403(.A1(new_n531), .A2(new_n536), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n490), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT91), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n377), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n379), .A2(new_n594), .ZN(new_n595));
  AOI211_X1 g409(.A(G902), .B(new_n593), .C1(new_n372), .C2(new_n375), .ZN(new_n596));
  NOR4_X1   g410(.A1(new_n591), .A2(new_n595), .A3(new_n586), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n276), .A2(new_n290), .ZN(new_n598));
  INV_X1    g412(.A(new_n277), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n298), .B1(new_n600), .B2(new_n291), .ZN(new_n601));
  INV_X1    g415(.A(new_n480), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT93), .B(G478), .Z(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n468), .B2(new_n351), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n459), .A2(new_n438), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n607), .B(new_n455), .C1(new_n451), .C2(new_n452), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n464), .B1(new_n608), .B2(new_n444), .ZN(new_n609));
  INV_X1    g423(.A(new_n467), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n466), .A2(new_n612), .A3(new_n467), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n470), .A2(G902), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n606), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n615), .ZN(new_n617));
  AOI211_X1 g431(.A(KEYINPUT92), .B(new_n617), .C1(new_n611), .C2(new_n613), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n605), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT94), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n466), .A2(new_n612), .A3(new_n467), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n612), .B1(new_n466), .B2(new_n467), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT92), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n614), .A2(new_n606), .A3(new_n615), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n605), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n602), .B(new_n487), .C1(new_n620), .C2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n597), .A2(new_n601), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT95), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT34), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n191), .ZN(G6));
  OR2_X1    g447(.A1(new_n472), .A2(new_n473), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n487), .A2(new_n634), .A3(new_n480), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n487), .A2(new_n634), .A3(KEYINPUT96), .A4(new_n480), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n597), .A2(new_n601), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n570), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT97), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n569), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n584), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n583), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n595), .A2(new_n596), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n301), .A2(new_n538), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT98), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT37), .B(G110), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  AND2_X1   g467(.A1(new_n359), .A2(G472), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n376), .A2(new_n377), .A3(new_n351), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT32), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n379), .A2(new_n361), .A3(new_n377), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n591), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n601), .A2(new_n647), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n487), .A2(new_n634), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n478), .A2(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n476), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XNOR2_X1  g481(.A(new_n663), .B(KEYINPUT39), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n537), .A2(KEYINPUT40), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT40), .B1(new_n537), .B2(new_n668), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n296), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n487), .A2(new_n474), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(new_n298), .A3(new_n647), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n352), .B1(new_n325), .B2(new_n333), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n374), .A2(KEYINPUT100), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n351), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT100), .B1(new_n374), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT101), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n684), .A2(KEYINPUT101), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n685), .B(new_n686), .C1(new_n378), .C2(new_n380), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n672), .A2(new_n679), .A3(KEYINPUT102), .A4(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n675), .A3(new_n678), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n670), .A2(new_n671), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n253), .ZN(G45));
  INV_X1    g508(.A(new_n487), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n627), .B1(new_n626), .B2(new_n605), .ZN(new_n696));
  AOI211_X1 g510(.A(KEYINPUT94), .B(new_n604), .C1(new_n624), .C2(new_n625), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n695), .B(new_n663), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n660), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n659), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NOR3_X1   g515(.A1(new_n504), .A2(KEYINPUT78), .A3(new_n506), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n514), .B1(new_n513), .B2(new_n505), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n518), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n528), .A2(new_n529), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n704), .A2(new_n533), .B1(new_n705), .B2(new_n534), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n490), .A3(new_n531), .ZN(new_n708));
  INV_X1    g522(.A(new_n601), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n381), .A2(new_n710), .A3(new_n629), .A4(new_n587), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT103), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  AND3_X1   g528(.A1(new_n637), .A2(new_n587), .A3(new_n638), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n381), .A2(new_n715), .A3(new_n710), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AOI21_X1  g531(.A(new_n648), .B1(new_n486), .B2(new_n488), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n381), .A2(new_n710), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  NAND3_X1  g534(.A1(new_n601), .A2(new_n676), .A3(new_n480), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n708), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n379), .A2(new_n723), .A3(new_n377), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n723), .B1(new_n379), .B2(new_n377), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n655), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n587), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  AND4_X1   g542(.A1(new_n723), .A2(new_n376), .A3(new_n377), .A4(new_n351), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n655), .B2(new_n725), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n487), .B(new_n664), .C1(new_n620), .C2(new_n628), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n647), .A3(new_n731), .A4(new_n710), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n658), .B2(new_n586), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n600), .A2(new_n294), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n292), .A2(KEYINPUT83), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n297), .A3(new_n737), .A4(new_n291), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n293), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(KEYINPUT105), .A3(new_n297), .A4(new_n737), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n537), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n620), .A2(new_n628), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n695), .A4(new_n663), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n381), .A2(KEYINPUT106), .A3(new_n587), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n735), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n381), .A2(new_n587), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n749), .A2(new_n698), .A3(new_n743), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n748), .B1(new_n750), .B2(KEYINPUT42), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  AND3_X1   g566(.A1(new_n740), .A2(new_n537), .A3(new_n742), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n661), .A2(new_n664), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n381), .A3(new_n587), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT107), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n658), .A2(new_n586), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n754), .A4(new_n753), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NAND2_X1  g575(.A1(new_n740), .A2(new_n742), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n520), .B1(new_n507), .B2(new_n515), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT45), .B1(new_n764), .B2(new_n532), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n516), .A2(new_n534), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  INV_X1    g581(.A(new_n532), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(G469), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(G469), .C1(new_n770), .C2(G902), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n531), .A3(new_n775), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n490), .A2(new_n763), .A3(new_n668), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n779), .B(new_n647), .C1(new_n595), .C2(new_n596), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n487), .B1(new_n696), .B2(new_n697), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT43), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n744), .A2(new_n783), .A3(new_n487), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n780), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n647), .B1(new_n595), .B2(new_n596), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n778), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n744), .B2(new_n487), .ZN(new_n789));
  AOI211_X1 g603(.A(KEYINPUT43), .B(new_n695), .C1(new_n620), .C2(new_n628), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n778), .A2(new_n791), .A3(new_n787), .A4(new_n780), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n777), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  NOR4_X1   g608(.A1(new_n381), .A2(new_n762), .A3(new_n587), .A4(new_n698), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n776), .A2(KEYINPUT47), .A3(new_n490), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT47), .B1(new_n776), .B2(new_n490), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(new_n635), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n736), .A2(new_n737), .A3(new_n291), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT84), .B1(new_n801), .B2(new_n297), .ZN(new_n802));
  INV_X1    g616(.A(new_n300), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT109), .B(new_n800), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n597), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT109), .B1(new_n301), .B2(new_n800), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n595), .A2(new_n596), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n537), .A2(new_n587), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n301), .A2(new_n808), .A3(new_n809), .A4(new_n629), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n588), .A2(new_n810), .A3(new_n650), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n711), .A2(new_n716), .A3(new_n719), .A4(new_n727), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n381), .A2(new_n537), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n487), .A2(new_n647), .A3(new_n474), .A4(new_n663), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n740), .A3(new_n742), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n726), .A2(new_n731), .A3(new_n647), .A4(new_n724), .ZN(new_n817));
  OAI22_X1  g631(.A1(new_n814), .A2(new_n816), .B1(new_n817), .B2(new_n743), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n812), .A2(new_n819), .A3(new_n760), .A4(new_n751), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n709), .A2(new_n677), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n583), .A2(new_n646), .A3(new_n663), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT111), .B1(new_n537), .B2(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(KEYINPUT111), .A2(new_n590), .A3(new_n822), .A4(new_n490), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n687), .B(new_n821), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n381), .B(new_n537), .C1(new_n699), .C2(new_n665), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n732), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n825), .A2(new_n732), .A3(new_n826), .A4(KEYINPUT52), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n820), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n833), .B2(KEYINPUT110), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n832), .B(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n476), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n791), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n708), .A3(new_n762), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n735), .A2(new_n747), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT48), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT48), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n587), .A2(new_n838), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n687), .A2(new_n762), .A3(new_n708), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n695), .A3(new_n744), .ZN(new_n847));
  INV_X1    g661(.A(G952), .ZN(new_n848));
  INV_X1    g662(.A(new_n730), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n839), .A2(new_n586), .A3(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n848), .B(G953), .C1(new_n850), .C2(new_n710), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n843), .A2(new_n844), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n675), .A2(new_n297), .A3(new_n708), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n849), .A2(new_n648), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n744), .A2(new_n695), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n840), .A2(new_n857), .B1(new_n846), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n850), .A2(new_n763), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n707), .A2(new_n531), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n490), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n796), .A2(new_n797), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n867), .B2(new_n861), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n852), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT114), .B1(new_n856), .B2(new_n859), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n867), .B(KEYINPUT112), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n861), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT53), .B1(new_n820), .B2(new_n831), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n805), .A2(new_n806), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n711), .A2(new_n716), .A3(new_n719), .A4(new_n727), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n588), .A2(new_n810), .A3(new_n650), .ZN(new_n877));
  INV_X1    g691(.A(new_n818), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n757), .A2(new_n731), .A3(new_n753), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT42), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n883), .A2(new_n748), .B1(new_n756), .B2(new_n759), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n879), .A2(new_n880), .A3(new_n833), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n836), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n837), .A2(new_n873), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n848), .A2(new_n269), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT115), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n587), .A2(new_n297), .A3(new_n490), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n675), .A2(new_n781), .A3(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n864), .B(KEYINPUT49), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n889), .A2(new_n891), .B1(new_n687), .B2(new_n895), .ZN(G75));
  NAND3_X1  g710(.A1(new_n250), .A2(new_n273), .A3(new_n275), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT116), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n271), .B(KEYINPUT55), .Z(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  INV_X1    g715(.A(new_n886), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(G210), .A3(G902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n903), .B2(KEYINPUT117), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(KEYINPUT117), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n848), .A2(G953), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT118), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n900), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n905), .A2(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n902), .A2(G902), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n771), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n706), .B(KEYINPUT119), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n874), .A2(new_n885), .A3(KEYINPUT54), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n887), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n772), .B(KEYINPUT57), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n920), .B2(KEYINPUT120), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n887), .B2(new_n916), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n915), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n908), .B1(new_n921), .B2(new_n924), .ZN(G54));
  INV_X1    g739(.A(new_n419), .ZN(new_n926));
  NAND2_X1  g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n913), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n913), .B2(new_n927), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n908), .B1(new_n928), .B2(new_n929), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT59), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n614), .B(KEYINPUT121), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n917), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n907), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n932), .B1(new_n837), .B2(new_n888), .ZN(new_n936));
  INV_X1    g750(.A(new_n933), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND4_X1  g754(.A1(new_n874), .A2(new_n885), .A3(new_n645), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n907), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n874), .A2(new_n885), .A3(new_n940), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n581), .B(KEYINPUT122), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT61), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n945), .B(new_n947), .Z(G66));
  NAND3_X1  g762(.A1(new_n477), .A2(G224), .A3(G953), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n807), .A2(new_n813), .A3(new_n811), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n951), .B2(G953), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n898), .B1(G898), .B2(new_n269), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n269), .A2(G900), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n793), .A2(new_n751), .A3(new_n760), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n776), .A2(new_n490), .A3(new_n668), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n821), .A3(new_n735), .A4(new_n747), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n732), .A2(new_n826), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n798), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT126), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n798), .A2(new_n961), .A3(new_n963), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n966), .A2(new_n884), .A3(new_n967), .A4(new_n793), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n956), .B(new_n958), .C1(new_n969), .C2(G953), .ZN(new_n970));
  AOI21_X1  g784(.A(G953), .B1(new_n965), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT127), .B1(new_n971), .B2(new_n957), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n369), .B(new_n400), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n537), .A2(new_n668), .ZN(new_n976));
  INV_X1    g790(.A(new_n661), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n744), .B2(new_n695), .ZN(new_n978));
  OR4_X1    g792(.A1(new_n749), .A2(new_n976), .A3(new_n762), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n793), .A2(new_n798), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n693), .B2(new_n962), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n963), .A2(new_n688), .A3(KEYINPUT62), .A4(new_n692), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n973), .B1(new_n984), .B2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n975), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n975), .B2(new_n986), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n993), .B(new_n835), .C1(new_n357), .C2(new_n374), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n969), .B2(new_n950), .ZN(new_n995));
  INV_X1    g809(.A(new_n370), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n345), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n984), .B2(new_n950), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n345), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n907), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n994), .A2(new_n997), .A3(new_n1000), .ZN(G57));
endmodule


