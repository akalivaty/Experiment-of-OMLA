

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U322 ( .A(n461), .B(n460), .ZN(n520) );
  XNOR2_X1 U323 ( .A(n340), .B(n339), .ZN(n341) );
  AND2_X1 U324 ( .A1(G227GAT), .A2(G233GAT), .ZN(n290) );
  OR2_X1 U325 ( .A1(n452), .A2(n451), .ZN(n453) );
  XOR2_X1 U326 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XNOR2_X1 U327 ( .A(KEYINPUT48), .B(KEYINPUT106), .ZN(n460) );
  OR2_X1 U328 ( .A1(n433), .A2(n432), .ZN(n434) );
  XNOR2_X1 U329 ( .A(n372), .B(n290), .ZN(n340) );
  XNOR2_X1 U330 ( .A(n438), .B(n437), .ZN(n439) );
  NOR2_X1 U331 ( .A1(n525), .A2(n381), .ZN(n363) );
  XNOR2_X1 U332 ( .A(n440), .B(n439), .ZN(n445) );
  XNOR2_X1 U333 ( .A(n344), .B(n343), .ZN(n514) );
  XNOR2_X1 U334 ( .A(KEYINPUT38), .B(n446), .ZN(n494) );
  XNOR2_X1 U335 ( .A(n468), .B(G169GAT), .ZN(n469) );
  XNOR2_X1 U336 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n447) );
  XNOR2_X1 U337 ( .A(n470), .B(n469), .ZN(G1348GAT) );
  XNOR2_X1 U338 ( .A(n448), .B(n447), .ZN(G1328GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n292) );
  XNOR2_X1 U340 ( .A(KEYINPUT6), .B(KEYINPUT89), .ZN(n291) );
  XNOR2_X1 U341 ( .A(n292), .B(n291), .ZN(n310) );
  XOR2_X1 U342 ( .A(G120GAT), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U343 ( .A(G29GAT), .B(G162GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U345 ( .A(G57GAT), .B(G1GAT), .Z(n296) );
  XNOR2_X1 U346 ( .A(G148GAT), .B(G155GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U348 ( .A(n298), .B(n297), .Z(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT0), .B(G134GAT), .Z(n300) );
  XNOR2_X1 U350 ( .A(G127GAT), .B(G113GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U352 ( .A(KEYINPUT80), .B(n301), .Z(n344) );
  XOR2_X1 U353 ( .A(G141GAT), .B(KEYINPUT2), .Z(n303) );
  XNOR2_X1 U354 ( .A(KEYINPUT88), .B(KEYINPUT3), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n350) );
  XOR2_X1 U356 ( .A(n350), .B(KEYINPUT5), .Z(n305) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n344), .B(n306), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n508) );
  XOR2_X1 U362 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n312) );
  NAND2_X1 U363 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U365 ( .A(G155GAT), .B(G22GAT), .Z(n349) );
  XOR2_X1 U366 ( .A(n313), .B(n349), .Z(n321) );
  XOR2_X1 U367 ( .A(KEYINPUT77), .B(G8GAT), .Z(n315) );
  XNOR2_X1 U368 ( .A(G211GAT), .B(G64GAT), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U370 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n317) );
  XNOR2_X1 U371 ( .A(KEYINPUT76), .B(KEYINPUT12), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G71GAT), .Z(n323) );
  XOR2_X1 U376 ( .A(G57GAT), .B(KEYINPUT13), .Z(n430) );
  XOR2_X1 U377 ( .A(G1GAT), .B(G15GAT), .Z(n415) );
  XNOR2_X1 U378 ( .A(n430), .B(n415), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(n325), .B(n324), .Z(n327) );
  XNOR2_X1 U381 ( .A(G127GAT), .B(G183GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n575) );
  XNOR2_X1 U383 ( .A(KEYINPUT91), .B(KEYINPUT26), .ZN(n364) );
  XOR2_X1 U384 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n329) );
  XNOR2_X1 U385 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U387 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n331) );
  XNOR2_X1 U388 ( .A(G190GAT), .B(G169GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n342) );
  XOR2_X1 U391 ( .A(KEYINPUT18), .B(KEYINPUT82), .Z(n335) );
  XNOR2_X1 U392 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U394 ( .A(G183GAT), .B(n336), .Z(n372) );
  XOR2_X1 U395 ( .A(G176GAT), .B(n428), .Z(n338) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(G99GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  INV_X1 U399 ( .A(n514), .ZN(n525) );
  INV_X1 U400 ( .A(G78GAT), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT69), .B(G204GAT), .Z(n346) );
  XNOR2_X1 U402 ( .A(G148GAT), .B(G106GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n429) );
  XOR2_X1 U405 ( .A(n429), .B(n349), .Z(n352) );
  XOR2_X1 U406 ( .A(G162GAT), .B(G50GAT), .Z(n391) );
  XNOR2_X1 U407 ( .A(n350), .B(n391), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U409 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n354) );
  NAND2_X1 U410 ( .A1(G228GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U412 ( .A(n356), .B(n355), .Z(n362) );
  XNOR2_X1 U413 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n357), .B(KEYINPUT87), .ZN(n358) );
  XOR2_X1 U415 ( .A(n358), .B(KEYINPUT21), .Z(n360) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(G211GAT), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n365), .B(KEYINPUT24), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n381) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n565) );
  XOR2_X1 U421 ( .A(G8GAT), .B(G169GAT), .Z(n413) );
  XOR2_X1 U422 ( .A(n413), .B(G204GAT), .Z(n367) );
  XNOR2_X1 U423 ( .A(G92GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U425 ( .A(G64GAT), .B(G176GAT), .Z(n436) );
  XOR2_X1 U426 ( .A(n436), .B(KEYINPUT75), .Z(n369) );
  NAND2_X1 U427 ( .A1(G226GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U429 ( .A(n371), .B(n370), .Z(n374) );
  XOR2_X1 U430 ( .A(G190GAT), .B(G36GAT), .Z(n392) );
  XNOR2_X1 U431 ( .A(n392), .B(n372), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n511) );
  XNOR2_X1 U433 ( .A(n511), .B(KEYINPUT27), .ZN(n382) );
  NOR2_X1 U434 ( .A1(n565), .A2(n382), .ZN(n375) );
  XOR2_X1 U435 ( .A(KEYINPUT92), .B(n375), .Z(n379) );
  INV_X1 U436 ( .A(n381), .ZN(n464) );
  NOR2_X1 U437 ( .A1(n511), .A2(n514), .ZN(n376) );
  NOR2_X1 U438 ( .A1(n464), .A2(n376), .ZN(n377) );
  XNOR2_X1 U439 ( .A(KEYINPUT25), .B(n377), .ZN(n378) );
  NAND2_X1 U440 ( .A1(n379), .A2(n378), .ZN(n380) );
  NAND2_X1 U441 ( .A1(n380), .A2(n508), .ZN(n386) );
  XOR2_X1 U442 ( .A(n381), .B(KEYINPUT28), .Z(n523) );
  OR2_X1 U443 ( .A1(n508), .A2(n382), .ZN(n521) );
  NOR2_X1 U444 ( .A1(n523), .A2(n521), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n383), .B(KEYINPUT90), .ZN(n384) );
  NAND2_X1 U446 ( .A1(n384), .A2(n514), .ZN(n385) );
  NAND2_X1 U447 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n387), .B(KEYINPUT93), .ZN(n475) );
  NOR2_X1 U449 ( .A1(n575), .A2(n475), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n388), .B(KEYINPUT98), .ZN(n409) );
  XOR2_X1 U451 ( .A(G92GAT), .B(G99GAT), .Z(n390) );
  XNOR2_X1 U452 ( .A(G85GAT), .B(KEYINPUT70), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n431) );
  XNOR2_X1 U454 ( .A(n391), .B(n431), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n399) );
  XOR2_X1 U456 ( .A(G43GAT), .B(KEYINPUT7), .Z(n395) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n416) );
  XOR2_X1 U459 ( .A(n416), .B(KEYINPUT73), .Z(n397) );
  NAND2_X1 U460 ( .A1(G232GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U462 ( .A(n399), .B(n398), .Z(n407) );
  XOR2_X1 U463 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n401) );
  XNOR2_X1 U464 ( .A(G134GAT), .B(G218GAT), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U466 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n403) );
  XNOR2_X1 U467 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n552) );
  XNOR2_X1 U471 ( .A(n552), .B(KEYINPUT97), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n408), .B(KEYINPUT36), .ZN(n579) );
  NAND2_X1 U473 ( .A1(n409), .A2(n579), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n410), .B(KEYINPUT37), .ZN(n507) );
  XOR2_X1 U475 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n412) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(G22GAT), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U478 ( .A(n414), .B(n413), .Z(n418) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U481 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n420) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U484 ( .A(n422), .B(n421), .Z(n427) );
  XOR2_X1 U485 ( .A(G197GAT), .B(G36GAT), .Z(n424) );
  XNOR2_X1 U486 ( .A(G113GAT), .B(G50GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n425), .B(KEYINPUT29), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n526) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U491 ( .A(n431), .B(n430), .Z(n432) );
  NAND2_X1 U492 ( .A1(n433), .A2(n432), .ZN(n435) );
  NAND2_X1 U493 ( .A1(n435), .A2(n434), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n436), .B(KEYINPUT68), .ZN(n438) );
  INV_X1 U495 ( .A(KEYINPUT32), .ZN(n437) );
  XOR2_X1 U496 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n442) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U499 ( .A(KEYINPUT33), .B(n443), .Z(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n572) );
  NOR2_X1 U501 ( .A1(n526), .A2(n572), .ZN(n479) );
  NAND2_X1 U502 ( .A1(n507), .A2(n479), .ZN(n446) );
  NOR2_X1 U503 ( .A1(n508), .A2(n494), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT105), .B(KEYINPUT46), .Z(n450) );
  XNOR2_X1 U505 ( .A(n572), .B(KEYINPUT41), .ZN(n541) );
  NOR2_X1 U506 ( .A1(n541), .A2(n526), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n452) );
  INV_X1 U508 ( .A(n575), .ZN(n562) );
  NAND2_X1 U509 ( .A1(n562), .A2(n552), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n453), .B(KEYINPUT47), .ZN(n459) );
  XOR2_X1 U511 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n455) );
  NAND2_X1 U512 ( .A1(n575), .A2(n579), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n456), .A2(n526), .ZN(n457) );
  NOR2_X1 U515 ( .A1(n572), .A2(n457), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n511), .A2(n520), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT54), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n463), .A2(n508), .ZN(n566) );
  NOR2_X1 U520 ( .A1(n464), .A2(n566), .ZN(n466) );
  INV_X1 U521 ( .A(KEYINPUT55), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n467), .A2(n525), .ZN(n561) );
  NOR2_X1 U524 ( .A1(n526), .A2(n561), .ZN(n470) );
  XNOR2_X1 U525 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n468) );
  INV_X1 U526 ( .A(G190GAT), .ZN(n474) );
  NOR2_X1 U527 ( .A1(n561), .A2(n552), .ZN(n472) );
  XNOR2_X1 U528 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n474), .B(n473), .ZN(G1351GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n477) );
  NAND2_X1 U532 ( .A1(n575), .A2(n552), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n477), .B(n476), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n475), .A2(n478), .ZN(n498) );
  NAND2_X1 U535 ( .A1(n479), .A2(n498), .ZN(n488) );
  NOR2_X1 U536 ( .A1(n508), .A2(n488), .ZN(n481) );
  XNOR2_X1 U537 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n482), .Z(G1324GAT) );
  NOR2_X1 U540 ( .A1(n511), .A2(n488), .ZN(n484) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n514), .A2(n488), .ZN(n486) );
  XNOR2_X1 U544 ( .A(KEYINPUT96), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  INV_X1 U547 ( .A(n523), .ZN(n517) );
  NOR2_X1 U548 ( .A1(n517), .A2(n488), .ZN(n489) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n489), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n511), .A2(n494), .ZN(n490) );
  XOR2_X1 U551 ( .A(G36GAT), .B(n490), .Z(G1329GAT) );
  NOR2_X1 U552 ( .A1(n494), .A2(n514), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT99), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NOR2_X1 U556 ( .A1(n494), .A2(n517), .ZN(n495) );
  XOR2_X1 U557 ( .A(G50GAT), .B(n495), .Z(G1331GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n497) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(KEYINPUT101), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n500) );
  INV_X1 U561 ( .A(n526), .ZN(n567) );
  XNOR2_X1 U562 ( .A(n541), .B(KEYINPUT100), .ZN(n555) );
  NOR2_X1 U563 ( .A1(n567), .A2(n555), .ZN(n506) );
  NAND2_X1 U564 ( .A1(n506), .A2(n498), .ZN(n503) );
  NOR2_X1 U565 ( .A1(n508), .A2(n503), .ZN(n499) );
  XOR2_X1 U566 ( .A(n500), .B(n499), .Z(G1332GAT) );
  NOR2_X1 U567 ( .A1(n511), .A2(n503), .ZN(n501) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n501), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n514), .A2(n503), .ZN(n502) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n502), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n507), .A2(n506), .ZN(n516) );
  NOR2_X1 U575 ( .A1(n508), .A2(n516), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT103), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n511), .A2(n516), .ZN(n512) );
  XOR2_X1 U579 ( .A(KEYINPUT104), .B(n512), .Z(n513) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n516), .ZN(n515) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT107), .ZN(n539) );
  NOR2_X1 U588 ( .A1(n523), .A2(n539), .ZN(n524) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n535) );
  NOR2_X1 U590 ( .A1(n526), .A2(n535), .ZN(n528) );
  XNOR2_X1 U591 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  NOR2_X1 U594 ( .A1(n555), .A2(n535), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U597 ( .A1(n562), .A2(n535), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT110), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  NOR2_X1 U601 ( .A1(n552), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT111), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n538), .Z(G1343GAT) );
  NOR2_X1 U605 ( .A1(n565), .A2(n539), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n547), .A2(n567), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  INV_X1 U608 ( .A(n547), .ZN(n551) );
  NOR2_X1 U609 ( .A1(n541), .A2(n551), .ZN(n543) );
  XNOR2_X1 U610 ( .A(KEYINPUT113), .B(KEYINPUT53), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U612 ( .A(n544), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT112), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n549) );
  NAND2_X1 U616 ( .A1(n547), .A2(n575), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT116), .B(n553), .Z(n554) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U622 ( .A1(n561), .A2(n555), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n557) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(KEYINPUT119), .B(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n580) );
  AND2_X1 U632 ( .A1(n567), .A2(n580), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n580), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT124), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1355GAT) );
endmodule

