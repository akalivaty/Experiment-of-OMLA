//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT82), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT81), .A2(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT81), .A2(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n190), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n191), .B2(new_n192), .ZN(new_n199));
  NOR2_X1   g013(.A1(G125), .A2(G140), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT16), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n193), .A2(KEYINPUT82), .A3(new_n195), .A4(new_n196), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n201), .A3(G146), .A4(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT83), .B(G110), .ZN(new_n212));
  AOI22_X1  g026(.A1(KEYINPUT79), .A2(new_n210), .B1(new_n207), .B2(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(KEYINPUT79), .B2(new_n210), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n213), .B(KEYINPUT80), .C1(KEYINPUT79), .C2(new_n210), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI211_X1 g032(.A(new_n211), .B(new_n212), .C1(new_n218), .C2(new_n209), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT24), .B(G110), .Z(new_n220));
  XNOR2_X1  g034(.A(G119), .B(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n203), .B(new_n206), .C1(new_n219), .C2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n198), .A2(new_n201), .A3(new_n202), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n205), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n203), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(new_n221), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n211), .B1(new_n218), .B2(new_n209), .ZN(new_n228));
  INV_X1    g042(.A(G110), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(G953), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(G221), .A3(G234), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n232), .B(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n230), .A3(new_n235), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n239), .B2(new_n188), .ZN(new_n240));
  AND4_X1   g054(.A1(KEYINPUT25), .A2(new_n237), .A3(new_n188), .A4(new_n238), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n189), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n189), .A2(G902), .ZN(new_n243));
  XOR2_X1   g057(.A(new_n243), .B(KEYINPUT84), .Z(new_n244));
  INV_X1    g058(.A(new_n239), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n256), .A3(G131), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n249), .A2(new_n251), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n250), .A2(G134), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT65), .A2(G131), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT65), .A2(G131), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT66), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n249), .A2(new_n251), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT65), .A2(G131), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n252), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n255), .B(new_n257), .C1(new_n263), .C2(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(KEYINPUT64), .A2(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT64), .A2(G143), .ZN(new_n274));
  AOI21_X1  g088(.A(G146), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n205), .A2(G143), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G143), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G146), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT64), .B(G143), .Z(new_n285));
  AOI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(G146), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n278), .A2(new_n282), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n258), .A2(new_n262), .A3(KEYINPUT66), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n270), .B1(new_n264), .B2(new_n269), .ZN(new_n289));
  OR3_X1    g103(.A1(new_n250), .A2(KEYINPUT68), .A3(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n290), .B(new_n291), .C1(new_n248), .C2(G137), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n288), .A2(new_n289), .B1(new_n292), .B2(G131), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n294));
  OAI21_X1  g108(.A(G128), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n275), .B2(new_n276), .ZN(new_n296));
  INV_X1    g110(.A(new_n284), .ZN(new_n297));
  INV_X1    g111(.A(G128), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n273), .A2(new_n274), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n299), .C1(new_n300), .C2(new_n205), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n272), .A2(new_n287), .B1(new_n293), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n207), .A2(G116), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G119), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G119), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G113), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G113), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT69), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT69), .B1(new_n313), .B2(new_n315), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n308), .B(new_n311), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g133(.A(new_n317), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT69), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n304), .A2(new_n306), .A3(new_n310), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n310), .B1(new_n304), .B2(new_n306), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n313), .A2(new_n315), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n309), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT28), .B1(new_n303), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n272), .A2(new_n287), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n288), .A2(new_n289), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n292), .A2(G131), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n302), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n330), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n303), .A2(new_n331), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n332), .B1(new_n340), .B2(KEYINPUT28), .ZN(new_n341));
  OR2_X1    g155(.A1(KEYINPUT74), .A2(G237), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT74), .A2(G237), .ZN(new_n343));
  AOI21_X1  g157(.A(G953), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G210), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT75), .B(KEYINPUT27), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n345), .B(new_n346), .Z(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G101), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n341), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT30), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n293), .B2(new_n302), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n354), .A2(new_n333), .A3(KEYINPUT72), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT72), .B1(new_n354), .B2(new_n333), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n330), .B1(new_n303), .B2(KEYINPUT30), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT73), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT72), .ZN(new_n360));
  INV_X1    g174(.A(new_n282), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n297), .B1(new_n300), .B2(new_n205), .ZN(new_n362));
  OAI22_X1  g176(.A1(new_n277), .A2(new_n361), .B1(new_n362), .B2(new_n279), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n253), .A2(new_n256), .A3(G131), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n289), .B2(new_n288), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n363), .B1(new_n365), .B2(new_n255), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n336), .A2(KEYINPUT30), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n354), .A2(new_n333), .A3(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT73), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n331), .B1(new_n337), .B2(new_n353), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n359), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n350), .A2(new_n339), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT31), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT31), .ZN(new_n378));
  AOI211_X1 g192(.A(new_n378), .B(new_n375), .C1(new_n359), .C2(new_n373), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n352), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n371), .B1(new_n370), .B2(new_n372), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n376), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n378), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(KEYINPUT31), .A3(new_n376), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n352), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G472), .A2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT32), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n337), .A2(new_n330), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n303), .A2(new_n331), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT28), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n332), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n350), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n339), .B1(new_n382), .B2(new_n383), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(new_n349), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT77), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n341), .B2(new_n404), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n350), .A2(KEYINPUT29), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n188), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G472), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT78), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n411), .B(G472), .C1(new_n403), .C2(new_n408), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n390), .A2(new_n394), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n388), .B1(new_n387), .B2(new_n352), .ZN(new_n414));
  AOI211_X1 g228(.A(KEYINPUT76), .B(new_n351), .C1(new_n385), .C2(new_n386), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n391), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n393), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n246), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT99), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n285), .A2(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n298), .A2(G143), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n420), .A2(new_n248), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n248), .B1(new_n420), .B2(new_n421), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G116), .B(G122), .ZN(new_n425));
  INV_X1    g239(.A(G107), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT98), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(KEYINPUT98), .A3(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n305), .A2(KEYINPUT14), .A3(G122), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(G107), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n419), .B1(new_n424), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n420), .A2(new_n421), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G134), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n420), .A2(new_n248), .A3(new_n421), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n441), .A2(KEYINPUT99), .A3(new_n431), .A4(new_n435), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n420), .A2(KEYINPUT13), .A3(new_n421), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n444), .B(G134), .C1(KEYINPUT13), .C2(new_n420), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n425), .B(new_n426), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT9), .B(G234), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n448), .A2(new_n187), .A3(G953), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n443), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n443), .B2(new_n447), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n188), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G478), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT100), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n443), .A2(new_n447), .ZN(new_n460));
  INV_X1    g274(.A(new_n449), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n443), .A2(new_n447), .A3(new_n449), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n458), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n188), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n468));
  AND2_X1   g282(.A1(G143), .A2(G214), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n344), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(KEYINPUT74), .A2(G237), .ZN(new_n471));
  NOR2_X1   g285(.A1(KEYINPUT74), .A2(G237), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n233), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT93), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n344), .A2(G214), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n470), .A2(new_n474), .B1(new_n475), .B2(new_n285), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT18), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n266), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n199), .A2(new_n200), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G146), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n476), .A2(new_n479), .B1(new_n206), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n470), .A2(new_n474), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n285), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n478), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G113), .B(G122), .ZN(new_n488));
  INV_X1    g302(.A(G104), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n480), .A2(KEYINPUT19), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n204), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n203), .B1(new_n496), .B2(G146), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n260), .A2(new_n261), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n476), .A2(new_n498), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(G475), .A2(G902), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n485), .A2(KEYINPUT17), .A3(new_n499), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n225), .A3(new_n203), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT95), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n509), .A3(new_n501), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT95), .A4(new_n509), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n511), .A2(new_n512), .B1(new_n486), .B2(new_n482), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n504), .B(new_n505), .C1(new_n513), .C2(new_n491), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT20), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n508), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n506), .A2(new_n225), .A3(new_n203), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n512), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n487), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n503), .B1(new_n519), .B2(new_n490), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n505), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n491), .A2(KEYINPUT96), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n518), .B2(new_n487), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n518), .A2(new_n524), .A3(new_n487), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n188), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n515), .A2(new_n522), .B1(G475), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT97), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n188), .ZN(new_n531));
  OAI21_X1  g345(.A(G475), .B1(new_n531), .B2(new_n525), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n521), .B1(new_n520), .B2(new_n505), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n491), .B1(new_n518), .B2(new_n487), .ZN(new_n534));
  INV_X1    g348(.A(new_n505), .ZN(new_n535));
  NOR4_X1   g349(.A1(new_n534), .A2(new_n503), .A3(KEYINPUT20), .A4(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n467), .B1(new_n530), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT3), .B1(new_n489), .B2(G107), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT3), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n426), .A3(G104), .ZN(new_n544));
  INV_X1    g358(.A(G101), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n489), .A2(G107), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n489), .A2(G107), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n426), .A2(G104), .ZN(new_n549));
  OAI21_X1  g363(.A(G101), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n302), .A2(KEYINPUT10), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G128), .B1(new_n275), .B2(new_n294), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n362), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n301), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n552), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT10), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G101), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT86), .B1(new_n562), .B2(KEYINPUT4), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT86), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT4), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n561), .A2(new_n564), .A3(new_n565), .A4(G101), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n547), .A2(KEYINPUT4), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n563), .A2(new_n566), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n287), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n272), .A2(KEYINPUT87), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n272), .A2(KEYINPUT87), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n560), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n558), .A2(new_n559), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n569), .A3(new_n553), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n272), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n233), .A2(G227), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT85), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G140), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT91), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n572), .A2(new_n580), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT89), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT88), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n296), .A2(new_n551), .A3(new_n586), .A4(new_n301), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT88), .B1(new_n302), .B2(new_n552), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n551), .B1(new_n556), .B2(new_n301), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n272), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n588), .A2(new_n589), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n272), .A2(new_n587), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n593), .A2(KEYINPUT89), .A3(KEYINPUT12), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n591), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n584), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT91), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n576), .A2(new_n599), .A3(new_n581), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n583), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G469), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n188), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n188), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n584), .A2(new_n575), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT90), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n597), .A2(new_n607), .A3(new_n572), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n581), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n597), .B2(new_n572), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n603), .B(new_n605), .C1(new_n611), .C2(new_n602), .ZN(new_n612));
  OAI21_X1  g426(.A(G221), .B1(new_n448), .B2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G952), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(G953), .ZN(new_n616));
  NAND2_X1  g430(.A1(G234), .A2(G237), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(G902), .A3(G953), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT21), .B(G898), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G214), .B1(G237), .B2(G902), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT6), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT5), .B1(new_n323), .B2(new_n324), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n304), .A2(KEYINPUT5), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n312), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n627), .A2(new_n629), .B1(new_n309), .B2(new_n328), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n330), .A2(new_n568), .B1(new_n552), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(G110), .B(G122), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n626), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n330), .A2(new_n568), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n630), .A2(new_n552), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n632), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n302), .A2(new_n194), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n363), .B2(new_n194), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n233), .A2(G224), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n641), .B(new_n642), .Z(new_n643));
  NAND3_X1  g457(.A1(new_n636), .A2(new_n626), .A3(new_n637), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT92), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT92), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n639), .A2(new_n647), .A3(new_n643), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(G210), .B1(G237), .B2(G902), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT7), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n641), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n641), .A2(new_n653), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n630), .A2(new_n551), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n632), .B(KEYINPUT8), .Z(new_n658));
  INV_X1    g472(.A(new_n629), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n309), .A2(KEYINPUT5), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n329), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n658), .B1(new_n661), .B2(new_n552), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n656), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n631), .A2(new_n632), .ZN(new_n664));
  AOI21_X1  g478(.A(G902), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n649), .A2(new_n650), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n650), .B1(new_n649), .B2(new_n665), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n624), .B(new_n625), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n541), .A2(new_n614), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n418), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT101), .B(G101), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G3));
  INV_X1    g487(.A(G472), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n390), .B2(new_n188), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n392), .B1(new_n381), .B2(new_n389), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n649), .A2(new_n665), .ZN(new_n678));
  INV_X1    g492(.A(new_n650), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(KEYINPUT102), .A3(new_n666), .ZN(new_n681));
  INV_X1    g495(.A(new_n625), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n668), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n452), .A2(G478), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n453), .A2(new_n188), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR3_X1    g502(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT33), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n464), .A2(KEYINPUT33), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(G478), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n530), .A2(new_n539), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n685), .A2(new_n694), .A3(new_n623), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n614), .A2(new_n246), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n677), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT34), .B(G104), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G6));
  OAI211_X1 g513(.A(new_n467), .B(new_n532), .C1(new_n533), .C2(new_n536), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n681), .A2(new_n684), .A3(new_n624), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n677), .A3(new_n696), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT35), .B(G107), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G9));
  INV_X1    g520(.A(new_n613), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n603), .A2(new_n605), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n611), .A2(new_n602), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n669), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n231), .B(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n244), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n242), .A2(new_n715), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n540), .A2(new_n710), .A3(new_n711), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n677), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT37), .B(G110), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G12));
  OAI21_X1  g534(.A(new_n394), .B1(new_n414), .B2(new_n415), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n410), .A2(new_n412), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n721), .B(new_n722), .C1(new_n676), .C2(KEYINPUT32), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n681), .A2(new_n684), .A3(new_n716), .ZN(new_n724));
  INV_X1    g538(.A(G900), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n619), .B1(new_n621), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT104), .B1(new_n700), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  INV_X1    g542(.A(new_n726), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n529), .A2(new_n728), .A3(new_n467), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n724), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n723), .A2(new_n732), .A3(new_n710), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n723), .A2(new_n732), .A3(new_n735), .A4(new_n710), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G128), .ZN(G30));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n726), .B(KEYINPUT39), .ZN(new_n740));
  OR3_X1    g554(.A1(new_n614), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n739), .B1(new_n614), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT40), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT40), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(new_n745), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n402), .A2(new_n350), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n188), .C1(new_n340), .C2(new_n350), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(G472), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n417), .A2(new_n721), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n716), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n667), .A2(new_n668), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT38), .ZN(new_n755));
  INV_X1    g569(.A(new_n467), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n530), .A2(new_n539), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n682), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n747), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n285), .ZN(G45));
  NAND4_X1  g575(.A1(new_n530), .A2(new_n539), .A3(new_n693), .A4(new_n729), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT107), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n724), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n723), .A2(new_n710), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n205), .ZN(G48));
  INV_X1    g582(.A(new_n246), .ZN(new_n769));
  INV_X1    g583(.A(new_n603), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n602), .B1(new_n601), .B2(new_n188), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n770), .A2(new_n771), .A3(new_n707), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n695), .A2(new_n723), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT108), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT41), .B(G113), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G15));
  NAND3_X1  g590(.A1(new_n703), .A2(new_n418), .A3(new_n772), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G116), .ZN(G18));
  NAND2_X1  g592(.A1(new_n601), .A2(new_n188), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(G469), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n613), .A3(new_n603), .A4(new_n624), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n723), .A2(new_n540), .A3(new_n765), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G119), .ZN(G21));
  NAND2_X1  g598(.A1(new_n406), .A2(new_n349), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n392), .B1(new_n387), .B2(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n675), .A2(new_n246), .A3(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n685), .A2(new_n781), .A3(new_n757), .A4(new_n756), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G122), .ZN(G24));
  INV_X1    g604(.A(new_n685), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n772), .ZN(new_n792));
  INV_X1    g606(.A(new_n786), .ZN(new_n793));
  AOI21_X1  g607(.A(G902), .B1(new_n381), .B2(new_n389), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n716), .B(new_n793), .C1(new_n794), .C2(new_n674), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n763), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G125), .ZN(G27));
  NAND2_X1  g612(.A1(new_n754), .A2(new_n625), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n710), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n614), .A2(KEYINPUT109), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(KEYINPUT42), .A3(new_n763), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT110), .B(new_n721), .C1(new_n676), .C2(KEYINPUT32), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n722), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT110), .B1(new_n417), .B2(new_n721), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n769), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(KEYINPUT111), .B(new_n769), .C1(new_n806), .C2(new_n807), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n804), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n801), .A2(new_n802), .ZN(new_n813));
  INV_X1    g627(.A(new_n799), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n723), .A2(new_n769), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT42), .B1(new_n817), .B2(new_n763), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n266), .ZN(G33));
  XNOR2_X1  g634(.A(new_n731), .B(KEYINPUT112), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n803), .A2(new_n418), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT113), .B(G134), .Z(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(G36));
  INV_X1    g638(.A(new_n677), .ZN(new_n825));
  NOR2_X1   g639(.A1(KEYINPUT115), .A2(KEYINPUT43), .ZN(new_n826));
  AND2_X1   g640(.A1(KEYINPUT115), .A2(KEYINPUT43), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n757), .B(new_n693), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n757), .A2(new_n693), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n830), .B2(new_n827), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n825), .A2(new_n716), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT44), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n814), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n611), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n602), .B1(new_n611), .B2(new_n838), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n604), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT46), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(new_n841), .B2(KEYINPUT46), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n770), .B1(new_n841), .B2(KEYINPUT46), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n613), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n740), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n837), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G137), .ZN(G39));
  NAND2_X1  g664(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n846), .B2(new_n613), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n846), .A2(new_n613), .A3(new_n851), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n723), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n763), .A2(new_n859), .A3(new_n246), .A4(new_n814), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(new_n196), .ZN(G42));
  NOR2_X1   g676(.A1(new_n770), .A2(new_n771), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(KEYINPUT49), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(KEYINPUT49), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n769), .A2(new_n613), .A3(new_n625), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n751), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n755), .A4(new_n830), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n723), .A2(new_n710), .A3(new_n765), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n763), .B1(new_n871), .B2(new_n796), .ZN(new_n872));
  INV_X1    g686(.A(new_n757), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n791), .A2(new_n467), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n614), .A3(new_n726), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n753), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n737), .A3(new_n876), .A4(KEYINPUT52), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n737), .A3(new_n876), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n878), .A3(new_n881), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n675), .A2(new_n786), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n763), .A2(new_n813), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n614), .B1(new_n413), .B2(new_n417), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n529), .A2(new_n756), .A3(new_n729), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n799), .A2(new_n752), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n822), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n757), .A2(new_n693), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n540), .A3(new_n669), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n677), .A3(new_n696), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n789), .A2(new_n896), .A3(new_n783), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n671), .A2(new_n718), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n893), .A2(new_n899), .A3(new_n774), .A4(new_n777), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n819), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n885), .A2(KEYINPUT53), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n782), .A2(new_n540), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n417), .B2(new_n413), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n905), .A2(new_n765), .B1(new_n787), .B2(new_n788), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n418), .A2(new_n670), .B1(new_n717), .B2(new_n677), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n777), .A4(new_n896), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT108), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n773), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n911), .B(new_n893), .C1(new_n818), .C2(new_n812), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n882), .A2(new_n877), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT118), .B1(new_n915), .B2(KEYINPUT54), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n831), .A2(new_n787), .A3(new_n619), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n864), .A2(new_n613), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n799), .B(new_n917), .C1(new_n858), .C2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n799), .A2(new_n864), .A3(new_n707), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n769), .A2(new_n869), .A3(new_n619), .A4(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n873), .A2(new_n693), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n831), .A2(new_n619), .A3(new_n923), .ZN(new_n926));
  INV_X1    g740(.A(new_n795), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n924), .A2(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n917), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n755), .A2(new_n682), .A3(new_n772), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n929), .A2(KEYINPUT50), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT50), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT119), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(KEYINPUT119), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n922), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n921), .B1(new_n920), .B2(new_n933), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n810), .A2(new_n811), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(KEYINPUT48), .A3(new_n926), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n924), .A2(new_n873), .A3(new_n693), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n940), .B(new_n616), .C1(new_n792), .C2(new_n917), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT48), .B1(new_n938), .B2(new_n926), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n936), .A2(new_n937), .A3(new_n939), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n885), .B2(new_n901), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n912), .A2(new_n913), .A3(new_n903), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT54), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT118), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT54), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n902), .A2(new_n914), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  AND4_X1   g764(.A1(new_n916), .A2(new_n944), .A3(new_n947), .A4(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(G952), .A2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n870), .B1(new_n951), .B2(new_n952), .ZN(G75));
  AOI21_X1  g767(.A(new_n188), .B1(new_n902), .B2(new_n914), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(G210), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n639), .A2(new_n644), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n643), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT55), .Z(new_n958));
  XOR2_X1   g772(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n959));
  AND3_X1   g773(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT56), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n233), .A2(G952), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(G51));
  XNOR2_X1  g778(.A(new_n604), .B(KEYINPUT57), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n902), .A2(new_n914), .A3(new_n949), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n949), .B1(new_n902), .B2(new_n914), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n601), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n954), .A2(new_n839), .A3(new_n840), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(G54));
  AND2_X1   g785(.A1(KEYINPUT58), .A2(G475), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n954), .A2(new_n520), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n520), .B1(new_n954), .B2(new_n972), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n974), .A3(new_n963), .ZN(G60));
  AND2_X1   g789(.A1(new_n689), .A2(new_n690), .ZN(new_n976));
  XNOR2_X1  g790(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(new_n687), .Z(new_n978));
  NOR2_X1   g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n966), .B2(new_n967), .ZN(new_n980));
  INV_X1    g794(.A(new_n963), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n916), .A2(new_n947), .A3(new_n950), .ZN(new_n983));
  INV_X1    g797(.A(new_n978), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n985), .B2(new_n976), .ZN(G63));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n915), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n963), .B1(new_n990), .B2(new_n245), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n902), .B2(new_n914), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n713), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT122), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n991), .B(new_n993), .C1(new_n994), .C2(KEYINPUT61), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n994), .B(new_n981), .C1(new_n992), .C2(new_n239), .ZN(new_n997));
  INV_X1    g811(.A(new_n993), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n981), .B1(new_n992), .B2(new_n239), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n996), .B(new_n997), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n995), .A2(new_n1000), .ZN(G66));
  INV_X1    g815(.A(new_n622), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n233), .B1(new_n1002), .B2(G224), .ZN(new_n1003));
  INV_X1    g817(.A(new_n911), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n233), .ZN(new_n1005));
  INV_X1    g819(.A(G898), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n956), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1005), .B(new_n1007), .ZN(G69));
  OR2_X1    g822(.A1(new_n858), .A2(new_n860), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n541), .B1(new_n757), .B2(new_n693), .ZN(new_n1010));
  OR4_X1    g824(.A1(new_n816), .A2(new_n743), .A3(new_n799), .A4(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n849), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT62), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n747), .A2(new_n759), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n872), .A2(new_n737), .A3(KEYINPUT123), .ZN(new_n1015));
  AOI21_X1  g829(.A(KEYINPUT123), .B1(new_n872), .B2(new_n737), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1013), .B(new_n1014), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT124), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT123), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n735), .B1(new_n888), .B2(new_n732), .ZN(new_n1021));
  AND4_X1   g835(.A1(new_n735), .A2(new_n723), .A3(new_n710), .A4(new_n732), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n792), .A2(new_n795), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n764), .B1(new_n1024), .B2(new_n766), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1020), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n872), .A2(new_n737), .A3(KEYINPUT123), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n760), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(KEYINPUT124), .B1(new_n1028), .B2(new_n1013), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1012), .B1(new_n1019), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT125), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1028), .A2(new_n1031), .A3(new_n1013), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1033));
  AOI21_X1  g847(.A(KEYINPUT125), .B1(new_n1033), .B2(KEYINPUT62), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n233), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n370), .B1(KEYINPUT30), .B2(new_n303), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(new_n496), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT127), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n233), .B1(G227), .B2(G900), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G900), .A2(G953), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT126), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1044), .B1(new_n819), .B2(new_n822), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n861), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1046));
  INV_X1    g860(.A(new_n822), .ZN(new_n1047));
  OAI211_X1 g861(.A(KEYINPUT126), .B(new_n1047), .C1(new_n812), .C2(new_n818), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n874), .B1(new_n810), .B2(new_n811), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n848), .B1(new_n837), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n1038), .B(new_n1043), .C1(new_n1051), .C2(G953), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1042), .A2(new_n1041), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n1042), .A2(new_n1041), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1031), .B1(new_n1028), .B2(new_n1013), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1033), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1028), .A2(KEYINPUT124), .A3(new_n1013), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1058), .A2(new_n1061), .A3(new_n1012), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1038), .B1(new_n1062), .B2(new_n233), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1064));
  INV_X1    g878(.A(new_n1051), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1064), .B1(new_n1065), .B2(new_n233), .ZN(new_n1066));
  OAI211_X1 g880(.A(new_n1054), .B(new_n1055), .C1(new_n1063), .C2(new_n1066), .ZN(new_n1067));
  AND2_X1   g881(.A1(new_n1053), .A2(new_n1067), .ZN(G72));
  OR2_X1    g882(.A1(new_n1062), .A2(new_n1004), .ZN(new_n1069));
  NAND2_X1  g883(.A1(G472), .A2(G902), .ZN(new_n1070));
  XOR2_X1   g884(.A(new_n1070), .B(KEYINPUT63), .Z(new_n1071));
  AOI21_X1  g885(.A(new_n748), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g886(.A(new_n402), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1073), .A2(new_n349), .ZN(new_n1074));
  NAND2_X1  g888(.A1(new_n1065), .A2(new_n911), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n1074), .B1(new_n1075), .B2(new_n1071), .ZN(new_n1076));
  NOR2_X1   g890(.A1(new_n945), .A2(new_n946), .ZN(new_n1077));
  OAI21_X1  g891(.A(new_n384), .B1(new_n1073), .B2(new_n350), .ZN(new_n1078));
  NAND2_X1  g892(.A1(new_n1078), .A2(new_n1071), .ZN(new_n1079));
  OAI21_X1  g893(.A(new_n981), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g894(.A1(new_n1072), .A2(new_n1076), .A3(new_n1080), .ZN(G57));
endmodule


