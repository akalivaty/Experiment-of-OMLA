//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT10), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .A4(G128), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n196), .A2(new_n204), .A3(KEYINPUT1), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(G128), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n196), .A2(new_n198), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n201), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n209));
  XNOR2_X1  g023(.A(G104), .B(G107), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G107), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n217), .A3(new_n211), .A4(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(G104), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n213), .A2(G107), .ZN(new_n221));
  OAI211_X1 g035(.A(KEYINPUT73), .B(G101), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n212), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n194), .B1(new_n208), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT75), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT4), .A3(new_n219), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n196), .A2(new_n198), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n196), .A2(new_n198), .A3(new_n230), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n207), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  XNOR2_X1  g050(.A(G143), .B(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n230), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n226), .A2(new_n240), .A3(G101), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n228), .A2(new_n233), .A3(new_n239), .A4(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n212), .A2(new_n219), .A3(new_n222), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n200), .B1(new_n245), .B2(new_n237), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(KEYINPUT10), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n248), .B(new_n194), .C1(new_n208), .C2(new_n223), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n225), .A2(new_n242), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(G137), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(G137), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT11), .A3(G134), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G131), .ZN(new_n258));
  INV_X1    g072(.A(G131), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n253), .A2(new_n256), .A3(new_n259), .A4(new_n254), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n250), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G140), .ZN(new_n263));
  INV_X1    g077(.A(G227), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n263), .B(new_n265), .Z(new_n266));
  AND2_X1   g080(.A1(new_n247), .A2(new_n242), .ZN(new_n267));
  INV_X1    g081(.A(new_n261), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n225), .A4(new_n249), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n262), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G469), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n208), .A2(new_n223), .ZN(new_n272));
  INV_X1    g086(.A(new_n246), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n223), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n261), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n261), .A2(KEYINPUT76), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT12), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n266), .B1(new_n278), .B2(new_n269), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT77), .B(new_n193), .C1(new_n271), .C2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n275), .B1(KEYINPUT12), .B2(new_n276), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n277), .B(new_n261), .C1(new_n272), .C2(new_n274), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n269), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n266), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n266), .B1(new_n262), .B2(new_n269), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n190), .B(new_n191), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n193), .B1(new_n271), .B2(new_n279), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n189), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G475), .ZN(new_n293));
  INV_X1    g107(.A(G125), .ZN(new_n294));
  OR3_X1    g108(.A1(new_n294), .A2(KEYINPUT16), .A3(G140), .ZN(new_n295));
  XOR2_X1   g109(.A(G125), .B(G140), .Z(new_n296));
  INV_X1    g110(.A(KEYINPUT16), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n195), .ZN(new_n299));
  OAI211_X1 g113(.A(G146), .B(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  INV_X1    g117(.A(G953), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G214), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(new_n197), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT17), .A3(G131), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(G131), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n305), .B(G143), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n259), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n302), .B(new_n307), .C1(KEYINPUT17), .C2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(G113), .B(G122), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(new_n213), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT18), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n309), .B1(new_n315), .B2(new_n259), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n296), .A2(G146), .ZN(new_n317));
  XNOR2_X1  g131(.A(G125), .B(G140), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n195), .ZN(new_n319));
  OAI221_X1 g133(.A(new_n316), .B1(new_n317), .B2(new_n319), .C1(new_n308), .C2(new_n315), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n312), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n311), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n300), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n318), .B(KEYINPUT19), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n195), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT84), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n314), .B1(new_n329), .B2(new_n320), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n293), .B(new_n191), .C1(new_n322), .C2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n321), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n335), .A2(KEYINPUT20), .A3(new_n293), .A4(new_n191), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n314), .B1(new_n312), .B2(new_n320), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n191), .B1(new_n322), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G475), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT86), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT13), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n244), .B2(G143), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n197), .A2(KEYINPUT85), .A3(KEYINPUT13), .A4(G128), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n197), .A2(G128), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n197), .A2(G128), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n346), .A2(new_n347), .B1(new_n348), .B2(new_n342), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n252), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n244), .A2(G143), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n351), .A3(new_n252), .ZN(new_n352));
  INV_X1    g166(.A(G116), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G122), .ZN(new_n354));
  INV_X1    g168(.A(G122), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G116), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n354), .A2(new_n356), .A3(new_n216), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n216), .B1(new_n354), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n352), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n341), .B1(new_n350), .B2(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n348), .A2(new_n351), .A3(new_n252), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(new_n356), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G107), .ZN(new_n363));
  XNOR2_X1  g177(.A(G116), .B(G122), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n216), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n361), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n244), .A2(G143), .ZN(new_n367));
  AOI22_X1  g181(.A1(KEYINPUT13), .A2(new_n367), .B1(new_n351), .B2(KEYINPUT85), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n343), .A2(new_n344), .ZN(new_n369));
  OAI21_X1  g183(.A(G134), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n370), .A3(KEYINPUT86), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT14), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n354), .A2(new_n356), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G107), .B1(new_n354), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n365), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n252), .B1(new_n348), .B2(new_n351), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n361), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n373), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n355), .A2(G116), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n216), .B1(new_n381), .B2(KEYINPUT14), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n354), .A2(new_n356), .A3(new_n374), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n382), .A2(new_n383), .B1(new_n216), .B2(new_n364), .ZN(new_n384));
  OAI21_X1  g198(.A(G134), .B1(new_n367), .B2(new_n346), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n352), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(KEYINPUT87), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n187), .A2(new_n389), .A3(G953), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n372), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n372), .B2(new_n388), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n191), .ZN(new_n395));
  INV_X1    g209(.A(G478), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(KEYINPUT15), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n395), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G952), .ZN(new_n399));
  AOI211_X1 g213(.A(G953), .B(new_n399), .C1(G234), .C2(G237), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n191), .B(new_n304), .C1(G234), .C2(G237), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT21), .B(G898), .Z(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n405), .B(KEYINPUT88), .Z(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n340), .A2(new_n398), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G116), .B(G119), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT5), .ZN(new_n410));
  INV_X1    g224(.A(G113), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n353), .A2(G119), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(KEYINPUT2), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G113), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT66), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(new_n409), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n420), .B1(new_n419), .B2(new_n409), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n415), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT78), .B1(new_n423), .B2(new_n223), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n417), .A2(G113), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n411), .A2(KEYINPUT2), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT65), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G119), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G116), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n353), .A2(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n416), .A2(new_n418), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n421), .B2(new_n422), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n241), .A3(new_n228), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT2), .B(G113), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT66), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n419), .A2(new_n409), .A3(new_n420), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n438), .A2(new_n439), .B1(new_n410), .B2(new_n414), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT78), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n243), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n424), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G122), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT79), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT79), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n443), .A2(new_n449), .A3(new_n444), .A4(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n200), .B(new_n294), .C1(new_n245), .C2(new_n237), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n235), .A2(G125), .A3(new_n238), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n202), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n207), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n294), .A4(new_n200), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G224), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n424), .A2(new_n436), .A3(new_n442), .A4(new_n445), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n463), .A2(KEYINPUT6), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n443), .A2(new_n446), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n451), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G113), .B1(new_n429), .B2(KEYINPUT5), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n410), .B1(new_n468), .B2(KEYINPUT81), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n469), .A2(new_n470), .B1(new_n421), .B2(new_n422), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n243), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n445), .B(KEYINPUT8), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n472), .B(new_n473), .C1(new_n243), .C2(new_n423), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(new_n460), .B2(G953), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n459), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT82), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n459), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  AND4_X1   g293(.A1(new_n463), .A2(new_n474), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n459), .A2(new_n475), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n467), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT83), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n467), .A2(new_n485), .A3(new_n483), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G214), .B1(G237), .B2(G902), .ZN(new_n491));
  AND4_X1   g305(.A1(new_n292), .A2(new_n408), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n494));
  NAND3_X1  g308(.A1(new_n303), .A2(new_n304), .A3(G210), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G101), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT70), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n261), .A2(new_n233), .A3(new_n239), .ZN(new_n500));
  INV_X1    g314(.A(new_n254), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n252), .A2(G137), .ZN(new_n502));
  OAI21_X1  g316(.A(G131), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n246), .A2(new_n260), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n409), .B1(new_n432), .B2(new_n437), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n427), .A2(new_n505), .B1(new_n438), .B2(new_n439), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n246), .A2(new_n260), .A3(new_n503), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n258), .A2(new_n260), .B1(new_n235), .B2(new_n238), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n435), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n507), .B2(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n507), .A2(new_n513), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n499), .B(new_n512), .C1(new_n514), .C2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n504), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n508), .B2(new_n509), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n522), .A3(new_n435), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT68), .ZN(new_n524));
  INV_X1    g338(.A(new_n498), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n520), .A2(new_n522), .A3(new_n526), .A4(new_n435), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n524), .A2(new_n507), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n519), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n493), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n512), .B1(new_n517), .B2(new_n514), .ZN(new_n536));
  INV_X1    g350(.A(new_n499), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n507), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n506), .B1(new_n500), .B2(new_n504), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT28), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n515), .A3(new_n525), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT29), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n524), .A2(new_n507), .A3(new_n527), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n498), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n539), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G472), .B1(new_n547), .B2(G902), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n528), .A2(new_n529), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n528), .A2(new_n529), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n518), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT32), .A3(new_n533), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n535), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n304), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT22), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(G137), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n428), .A2(G128), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n244), .A2(G119), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT24), .B(G110), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OR3_X1    g376(.A1(new_n428), .A2(KEYINPUT23), .A3(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(KEYINPUT23), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n563), .A2(new_n564), .B1(new_n428), .B2(G128), .ZN(new_n565));
  INV_X1    g379(.A(G110), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n301), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n565), .A2(new_n566), .B1(new_n560), .B2(new_n561), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n570), .A2(new_n325), .A3(new_n317), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n557), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n568), .A3(new_n556), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n574), .A3(new_n191), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT25), .ZN(new_n576));
  NAND2_X1  g390(.A1(G217), .A2(G902), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n389), .B2(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT72), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n572), .A2(new_n574), .A3(new_n580), .A4(new_n191), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n576), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n572), .A2(new_n574), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n553), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n492), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  INV_X1    g405(.A(new_n292), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n551), .A2(new_n191), .ZN(new_n593));
  INV_X1    g407(.A(G472), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT89), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n593), .B(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n592), .A2(new_n596), .A3(new_n586), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n333), .A2(new_n336), .A3(new_n339), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n392), .B2(new_n393), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n391), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n360), .A2(new_n371), .B1(new_n380), .B2(new_n387), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT92), .A3(new_n390), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n604), .A3(KEYINPUT33), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT91), .B1(new_n603), .B2(new_n390), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n350), .A2(new_n359), .A3(new_n341), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT86), .B1(new_n366), .B2(new_n370), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n377), .A2(new_n379), .A3(new_n373), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT87), .B1(new_n384), .B2(new_n386), .ZN(new_n610));
  OAI22_X1  g424(.A1(new_n607), .A2(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT91), .ZN(new_n612));
  INV_X1    g426(.A(new_n390), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n600), .B1(new_n605), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G478), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n394), .A2(new_n396), .A3(new_n191), .ZN(new_n618));
  NAND2_X1  g432(.A1(G478), .A2(G902), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT93), .ZN(new_n621));
  OAI21_X1  g435(.A(G478), .B1(new_n616), .B2(G902), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n598), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(KEYINPUT94), .B(new_n598), .C1(new_n621), .C2(new_n624), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n467), .A2(KEYINPUT90), .A3(new_n485), .A4(new_n483), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT90), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n489), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n474), .A2(new_n477), .A3(new_n463), .A4(new_n479), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n191), .B1(new_n633), .B2(new_n481), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n448), .A2(new_n450), .B1(new_n464), .B2(new_n465), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n462), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n485), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n491), .B(new_n630), .C1(new_n632), .C2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n407), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n597), .A2(new_n629), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  NAND2_X1  g456(.A1(new_n598), .A2(new_n398), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n638), .A2(new_n407), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n597), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  INV_X1    g461(.A(new_n596), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n573), .A2(new_n568), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n584), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n582), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT95), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n492), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT37), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n566), .ZN(G12));
  NAND2_X1  g471(.A1(new_n630), .A2(new_n491), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n636), .A2(new_n485), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT90), .B1(new_n636), .B2(new_n485), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n292), .A2(new_n553), .A3(new_n661), .A4(new_n654), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n400), .B1(new_n402), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n598), .A2(new_n398), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n244), .ZN(G30));
  NAND2_X1  g482(.A1(new_n490), .A2(KEYINPUT96), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n488), .A2(new_n670), .A3(new_n489), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n669), .A2(KEYINPUT38), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT38), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n528), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n540), .A2(new_n541), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n675), .B1(new_n676), .B2(new_n499), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n677), .B2(G902), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n535), .A2(new_n552), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n491), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n340), .A2(new_n398), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n664), .B(KEYINPUT39), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n292), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n291), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n280), .A2(new_n287), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n188), .B(new_n685), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n686), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n653), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n674), .A2(new_n683), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT98), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n197), .ZN(G45));
  AND4_X1   g511(.A1(new_n623), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n623), .B1(new_n622), .B2(new_n618), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n340), .B(new_n665), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n662), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT99), .B(G146), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G48));
  OAI21_X1  g517(.A(new_n191), .B1(new_n285), .B2(new_n286), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n188), .A3(new_n287), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n553), .A2(new_n661), .A3(new_n587), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n629), .A2(new_n708), .A3(new_n639), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT41), .B(G113), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n709), .B(new_n711), .ZN(G15));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n644), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR2_X1   g528(.A1(new_n638), .A2(new_n706), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n553), .A3(new_n408), .A4(new_n654), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NOR3_X1   g531(.A1(new_n638), .A2(new_n682), .A3(new_n706), .ZN(new_n718));
  INV_X1    g532(.A(new_n542), .ZN(new_n719));
  INV_X1    g533(.A(new_n515), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n499), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n549), .B2(new_n550), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n593), .A2(G472), .B1(new_n533), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT101), .B1(new_n723), .B2(new_n587), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n533), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n528), .B(new_n529), .ZN(new_n726));
  AOI21_X1  g540(.A(G902), .B1(new_n726), .B2(new_n518), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n587), .B(new_n725), .C1(new_n727), .C2(new_n594), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n718), .B(new_n406), .C1(new_n724), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  OAI21_X1  g546(.A(new_n725), .B1(new_n727), .B2(new_n594), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n694), .ZN(new_n734));
  INV_X1    g548(.A(new_n700), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n715), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  NAND3_X1  g551(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n283), .A2(new_n284), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n283), .A2(KEYINPUT102), .A3(new_n284), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(G469), .A3(new_n270), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n193), .A3(new_n287), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n188), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n700), .A2(new_n738), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n535), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(KEYINPUT104), .B(new_n493), .C1(new_n532), .C2(new_n534), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n548), .A3(new_n552), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n587), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n744), .A2(new_n188), .ZN(new_n754));
  INV_X1    g568(.A(new_n738), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n625), .A3(new_n665), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n753), .B1(new_n756), .B2(new_n588), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n751), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  NOR4_X1   g573(.A1(new_n588), .A2(new_n666), .A3(new_n738), .A4(new_n745), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n252), .ZN(G36));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n340), .B1(new_n621), .B2(new_n624), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n763), .B2(KEYINPUT107), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n698), .A2(new_n699), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n765), .B(KEYINPUT43), .C1(new_n766), .C2(new_n340), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n767), .A3(new_n596), .A4(new_n653), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n738), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n741), .A2(KEYINPUT45), .A3(new_n270), .A4(new_n742), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT106), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n262), .A2(new_n266), .A3(new_n269), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n740), .B2(new_n739), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n774), .A2(new_n775), .A3(KEYINPUT45), .A4(new_n742), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  OAI22_X1  g592(.A1(new_n271), .A2(new_n279), .B1(new_n778), .B2(new_n190), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT105), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI221_X1 g595(.A(KEYINPUT105), .B1(new_n778), .B2(new_n190), .C1(new_n271), .C2(new_n279), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n193), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n772), .A2(new_n776), .B1(new_n781), .B2(new_n782), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n786), .B1(new_n787), .B2(new_n192), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n788), .A3(new_n287), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n188), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n684), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n768), .A2(new_n769), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n768), .A2(KEYINPUT108), .A3(new_n769), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n770), .B(new_n791), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT109), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n255), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n287), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n784), .A2(new_n193), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n804), .B2(new_n786), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n189), .B1(new_n805), .B2(new_n785), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n802), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n700), .A2(new_n738), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n553), .A2(new_n587), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n790), .A2(new_n801), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  NAND2_X1  g627(.A1(new_n399), .A2(new_n304), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n681), .B1(new_n488), .B2(new_n489), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n643), .B1(new_n766), .B2(new_n598), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n597), .A2(new_n406), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n655), .A3(new_n590), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n709), .A2(new_n713), .A3(new_n716), .A4(new_n731), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n723), .A2(KEYINPUT101), .A3(new_n587), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n728), .A2(new_n729), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n407), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n826), .A2(new_n718), .B1(new_n708), .B2(new_n644), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(KEYINPUT111), .A3(new_n709), .A4(new_n716), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n820), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n625), .A2(new_n723), .A3(new_n653), .A4(new_n665), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n661), .A2(new_n707), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n662), .A2(new_n666), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n701), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n582), .A2(new_n652), .A3(new_n665), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n582), .A2(KEYINPUT114), .A3(new_n652), .A4(new_n665), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n745), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n638), .A2(new_n682), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n679), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n833), .A2(KEYINPUT52), .A3(new_n834), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n842), .B(new_n736), .C1(new_n666), .C2(new_n662), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(new_n701), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n760), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n746), .A2(new_n734), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n340), .A2(new_n398), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n755), .A2(new_n850), .A3(new_n665), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n292), .A2(new_n553), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n755), .A2(KEYINPUT112), .A3(new_n850), .A4(new_n665), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n654), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n758), .A2(new_n848), .A3(new_n849), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n816), .A2(new_n829), .A3(new_n847), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n736), .B(new_n861), .C1(new_n666), .C2(new_n662), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(new_n834), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n820), .B1(new_n864), .B2(new_n846), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n857), .A2(new_n821), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n816), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n815), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n829), .A2(new_n847), .A3(new_n858), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT53), .B1(new_n864), .B2(new_n846), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n829), .A2(new_n871), .A3(new_n858), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(KEYINPUT54), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n750), .A2(new_n587), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n764), .A2(new_n767), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n738), .A2(new_n706), .A3(new_n401), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT48), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT117), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT116), .Z(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(new_n882), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n883), .B(new_n884), .C1(KEYINPUT117), .C2(new_n879), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n679), .A2(new_n586), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n877), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n629), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n885), .A2(G952), .A3(new_n304), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n764), .A2(new_n767), .A3(new_n400), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n724), .A2(new_n730), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n890), .A2(new_n891), .A3(new_n706), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n889), .B1(new_n661), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n868), .A2(new_n873), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n876), .A2(new_n734), .A3(new_n877), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n598), .A3(new_n766), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n674), .A2(new_n491), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n892), .A2(KEYINPUT50), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT50), .B1(new_n892), .B2(new_n897), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n895), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n890), .A2(new_n891), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n808), .A2(new_n811), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n705), .A2(new_n287), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n189), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n738), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n900), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT51), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n902), .A2(new_n904), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n910), .A2(new_n755), .A3(new_n901), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT115), .B(new_n909), .C1(new_n911), .C2(new_n900), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n814), .B1(new_n894), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n674), .A2(new_n766), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n340), .A2(new_n189), .A3(new_n681), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n903), .B(KEYINPUT49), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n915), .A2(new_n886), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n914), .A2(new_n918), .ZN(G75));
  NAND2_X1  g733(.A1(new_n864), .A2(new_n846), .ZN(new_n920));
  INV_X1    g734(.A(new_n820), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n866), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT53), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n829), .A2(new_n816), .A3(new_n847), .A4(new_n858), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n924), .A3(G902), .A4(new_n487), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n823), .A2(new_n828), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n847), .A2(new_n928), .A3(new_n921), .A4(new_n858), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n867), .B1(new_n929), .B2(new_n816), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(KEYINPUT118), .A3(G902), .A4(new_n487), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n635), .B(new_n462), .Z(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n927), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n304), .A2(G952), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n923), .A2(new_n924), .A3(G210), .A4(G902), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n939), .B2(new_n933), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n935), .A2(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n192), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n923), .A2(KEYINPUT54), .A3(new_n924), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT54), .B1(new_n923), .B2(new_n924), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n285), .A2(new_n286), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n787), .B(KEYINPUT120), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n930), .A2(G902), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n936), .B1(new_n948), .B2(new_n950), .ZN(G54));
  NAND4_X1  g765(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT58), .A4(G902), .ZN(new_n952));
  INV_X1    g766(.A(new_n335), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n952), .A2(new_n293), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n936), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n952), .B2(new_n293), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(G60));
  INV_X1    g771(.A(new_n616), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n619), .B(KEYINPUT59), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n958), .B(new_n960), .C1(new_n944), .C2(new_n945), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n868), .B2(new_n873), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n961), .B(new_n955), .C1(new_n962), .C2(new_n958), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(G63));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n577), .B(KEYINPUT60), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n923), .A2(new_n924), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n583), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n651), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n955), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n965), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n930), .A2(new_n651), .A3(new_n967), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n975), .A2(KEYINPUT61), .A3(new_n955), .A4(new_n970), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G66));
  INV_X1    g791(.A(new_n404), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n978), .B2(new_n460), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n829), .B2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT121), .ZN(new_n981));
  INV_X1    g795(.A(new_n635), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(G898), .B2(new_n304), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n981), .B(new_n983), .ZN(G69));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n985));
  OAI21_X1  g799(.A(G953), .B1(new_n264), .B2(new_n663), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT123), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n520), .A2(new_n522), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n326), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n860), .A2(new_n695), .A3(new_n834), .A4(new_n862), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT122), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(KEYINPUT122), .B2(new_n991), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT122), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n990), .A2(new_n995), .A3(KEYINPUT62), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n994), .A2(new_n796), .A3(new_n812), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n589), .A2(new_n818), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n998), .A2(new_n690), .A3(new_n738), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n304), .B(new_n989), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n789), .A2(new_n188), .A3(new_n685), .A4(new_n841), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n874), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n812), .A2(new_n796), .A3(new_n1003), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1002), .A2(new_n1001), .A3(new_n874), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n760), .B1(new_n757), .B2(new_n751), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n860), .A2(new_n834), .A3(new_n862), .ZN(new_n1008));
  OR3_X1    g822(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n304), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n663), .A2(G953), .ZN(new_n1011));
  INV_X1    g825(.A(new_n989), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n985), .B(new_n987), .C1(new_n1000), .C2(new_n1013), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n987), .A2(new_n985), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n987), .A2(new_n985), .ZN(new_n1016));
  AND4_X1   g830(.A1(new_n1015), .A2(new_n1000), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1014), .A2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(new_n928), .A2(new_n921), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1019), .A2(new_n857), .ZN(new_n1020));
  AOI22_X1  g834(.A1(new_n1020), .A2(new_n871), .B1(new_n869), .B2(KEYINPUT53), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT127), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n528), .A2(KEYINPUT126), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n546), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1026), .A2(new_n546), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1021), .A2(new_n1022), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n870), .A2(new_n872), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(KEYINPUT127), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n812), .A2(new_n796), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1033), .A2(new_n829), .A3(new_n1003), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n545), .B1(new_n1035), .B2(new_n1024), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n936), .B1(new_n1036), .B2(new_n498), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n997), .A2(new_n1019), .A3(new_n999), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n525), .B(new_n545), .C1(new_n1038), .C2(new_n1025), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1032), .A2(new_n1037), .A3(new_n1039), .ZN(G57));
endmodule


