//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT27), .B(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n206), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n212), .A3(new_n209), .ZN(new_n213));
  OR2_X1    g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(new_n213), .C1(KEYINPUT26), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT28), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n204), .A2(new_n216), .A3(new_n205), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n207), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  AND3_X1   g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(new_n209), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n227), .B2(KEYINPUT65), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n224), .A2(new_n229), .A3(new_n226), .A4(new_n209), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  NOR4_X1   g034(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n224), .A2(KEYINPUT25), .A3(new_n226), .A4(new_n209), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n218), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G120gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G113gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G127gat), .B(G134gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n249));
  INV_X1    g048(.A(G127gat), .ZN(new_n250));
  OR3_X1    g049(.A1(new_n250), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253));
  AND4_X1   g052(.A1(new_n253), .A2(new_n245), .A3(new_n248), .A4(new_n246), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT1), .B1(new_n242), .B2(new_n244), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n255), .B2(new_n248), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT70), .B(new_n252), .C1(new_n254), .C2(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n203), .B1(new_n240), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n207), .A2(new_n215), .A3(new_n217), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT25), .B1(new_n228), .B2(new_n230), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n238), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n265), .A2(KEYINPUT71), .A3(new_n259), .A4(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n240), .A2(new_n261), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT32), .ZN(new_n271));
  XNOR2_X1  g070(.A(G15gat), .B(G43gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT72), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n277), .B(KEYINPUT33), .C1(new_n268), .C2(new_n269), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n271), .B(new_n274), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n268), .A2(new_n269), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT34), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n274), .A2(KEYINPUT33), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n270), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT22), .ZN(new_n288));
  INV_X1    g087(.A(G211gat), .ZN(new_n289));
  INV_X1    g088(.A(G218gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n301));
  OAI21_X1  g100(.A(G141gat), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(G141gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT78), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n303), .B2(G141gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  INV_X1    g108(.A(G155gat), .ZN(new_n310));
  INV_X1    g109(.A(G162gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(new_n312), .B2(KEYINPUT2), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(G148gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n304), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n312), .A2(new_n309), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n299), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G228gat), .A2(G233gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n294), .B(KEYINPUT74), .Z(new_n325));
  AOI22_X1  g124(.A1(new_n308), .A2(new_n313), .B1(new_n319), .B2(new_n318), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n326), .B2(new_n298), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n322), .B(new_n324), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n323), .B(KEYINPUT84), .Z(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n297), .B2(new_n298), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n327), .A2(new_n295), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G22gat), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT85), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(KEYINPUT85), .A3(new_n336), .ZN(new_n340));
  XOR2_X1   g139(.A(G78gat), .B(G106gat), .Z(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT31), .B(G50gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n340), .A2(new_n344), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n282), .B1(new_n279), .B2(new_n284), .ZN(new_n348));
  NOR4_X1   g147(.A1(new_n286), .A2(new_n347), .A3(new_n348), .A4(KEYINPUT35), .ZN(new_n349));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT75), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n265), .B2(new_n296), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n354), .B(KEYINPUT76), .Z(new_n357));
  OAI22_X1  g156(.A1(new_n356), .A2(KEYINPUT77), .B1(new_n240), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n359));
  AOI211_X1 g158(.A(new_n359), .B(new_n355), .C1(new_n265), .C2(new_n296), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n358), .A2(new_n294), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n325), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n240), .A2(new_n354), .ZN(new_n363));
  INV_X1    g162(.A(new_n357), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n265), .B2(new_n296), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n352), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n240), .A2(new_n357), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n354), .B1(new_n240), .B2(KEYINPUT29), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(new_n359), .ZN(new_n371));
  INV_X1    g170(.A(new_n360), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n295), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n352), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n366), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(new_n375), .A3(KEYINPUT30), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n373), .A2(new_n366), .A3(new_n377), .A4(new_n374), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n376), .A2(KEYINPUT86), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT86), .B1(new_n376), .B2(new_n378), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  INV_X1    g182(.A(G85gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n245), .A2(new_n248), .A3(new_n246), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT69), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n255), .A2(new_n253), .A3(new_n248), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT70), .B1(new_n393), .B2(new_n252), .ZN(new_n394));
  INV_X1    g193(.A(new_n260), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n389), .B(new_n326), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n261), .A2(KEYINPUT80), .A3(new_n389), .A4(new_n326), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(KEYINPUT4), .C1(new_n257), .C2(new_n321), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(new_n326), .A3(new_n252), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n403), .B2(KEYINPUT4), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n398), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n326), .A2(new_n298), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n257), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT5), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n406), .A2(KEYINPUT82), .A3(new_n409), .A4(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n409), .A2(KEYINPUT4), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n411), .B1(new_n418), .B2(new_n403), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n326), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n257), .A2(new_n321), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n422), .A2(new_n403), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT5), .B1(new_n423), .B2(new_n410), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n388), .B1(new_n417), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n382), .B1(new_n427), .B2(KEYINPUT6), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n415), .B2(new_n416), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  NOR4_X1   g229(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n430), .A4(new_n388), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n388), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n381), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n349), .B1(new_n436), .B2(KEYINPUT90), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n430), .B1(new_n429), .B2(new_n388), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n387), .B(new_n425), .C1(new_n415), .C2(new_n416), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n440), .A2(new_n428), .A3(new_n431), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n441), .A2(new_n442), .A3(new_n381), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n202), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n441), .B2(new_n381), .ZN(new_n445));
  INV_X1    g244(.A(new_n428), .ZN(new_n446));
  INV_X1    g245(.A(new_n431), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n435), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n381), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT90), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT91), .A4(new_n349), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n279), .A2(new_n284), .ZN(new_n452));
  INV_X1    g251(.A(new_n282), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT73), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n285), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n348), .A2(KEYINPUT73), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n347), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n376), .A2(new_n378), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n448), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n451), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n410), .B1(new_n406), .B2(new_n409), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n387), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n423), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT39), .B1(new_n466), .B2(new_n411), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n469), .A2(KEYINPUT40), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(KEYINPUT40), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n381), .A2(new_n470), .A3(new_n433), .A4(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n373), .A2(new_n474), .A3(new_n366), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n352), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n373), .B2(new_n366), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n295), .B1(new_n371), .B2(new_n372), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n363), .A2(new_n362), .A3(new_n365), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT37), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n473), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(new_n352), .A3(new_n482), .A4(new_n475), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n478), .A2(new_n375), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n432), .A2(new_n435), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n347), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n472), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT36), .B1(new_n454), .B2(new_n285), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n456), .A2(new_n457), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(KEYINPUT36), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n448), .B2(new_n459), .ZN(new_n491));
  OR3_X1    g290(.A1(new_n487), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(G1gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G1gat), .B2(new_n494), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n497), .B(G8gat), .Z(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  INV_X1    g300(.A(G36gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT92), .B1(new_n506), .B2(new_n500), .ZN(new_n507));
  OAI22_X1  g306(.A1(new_n505), .A2(new_n507), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT93), .ZN(new_n513));
  INV_X1    g312(.A(new_n511), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n503), .A2(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n510), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n498), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(KEYINPUT17), .A3(new_n517), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n498), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT17), .B1(new_n513), .B2(new_n517), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n519), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT94), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT18), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n517), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n498), .A3(new_n521), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(new_n519), .A3(new_n520), .A4(new_n526), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n520), .B(KEYINPUT13), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n517), .A3(new_n498), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n537), .B2(new_n518), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT95), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(KEYINPUT95), .B(new_n535), .C1(new_n537), .C2(new_n518), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n528), .A2(new_n533), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  INV_X1    g343(.A(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT11), .B(G169gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n546), .B(new_n547), .Z(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT12), .Z(new_n549));
  AND3_X1   g348(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n543), .B1(new_n542), .B2(new_n549), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n550), .A2(new_n551), .B1(new_n542), .B2(new_n549), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(G71gat), .B(G78gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT97), .B(G57gat), .ZN(new_n556));
  INV_X1    g355(.A(G64gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n557), .A2(G57gat), .ZN(new_n559));
  AND2_X1   g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  OAI22_X1  g359(.A1(new_n558), .A2(new_n559), .B1(KEYINPUT9), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n555), .B1(new_n561), .B2(KEYINPUT98), .ZN(new_n562));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n555), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n384), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n384), .B2(new_n570), .ZN(new_n573));
  NAND3_X1  g372(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G99gat), .B(G106gat), .Z(new_n576));
  OAI21_X1  g375(.A(KEYINPUT102), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n568), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n575), .B(new_n576), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n568), .A2(new_n581), .A3(new_n577), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT10), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n568), .A2(KEYINPUT10), .A3(new_n579), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n554), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n582), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n554), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n553), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT99), .B(KEYINPUT21), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n562), .A2(new_n567), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(new_n250), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G155gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G183gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(new_n289), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n598), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n498), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n568), .B2(KEYINPUT21), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n602), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT41), .ZN(new_n608));
  INV_X1    g407(.A(G232gat), .ZN(new_n609));
  INV_X1    g408(.A(G233gat), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n529), .B2(new_n579), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n521), .A2(new_n581), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n613), .B2(new_n523), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  INV_X1    g417(.A(new_n615), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT100), .B(G134gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G162gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n616), .A2(new_n620), .A3(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n607), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n594), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n493), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n441), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n449), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  AOI21_X1  g435(.A(KEYINPUT42), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  OAI21_X1  g437(.A(G8gat), .B1(new_n631), .B2(new_n449), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n640), .B2(KEYINPUT42), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI211_X1 g442(.A(KEYINPUT103), .B(new_n637), .C1(new_n640), .C2(KEYINPUT42), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n490), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n631), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n286), .A2(new_n348), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n646), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n631), .A2(new_n486), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  NOR3_X1   g453(.A1(new_n487), .A2(new_n490), .A3(new_n491), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n445), .A2(new_n450), .A3(new_n349), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n656), .A2(new_n202), .B1(KEYINPUT35), .B2(new_n460), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n657), .B2(new_n451), .ZN(new_n658));
  INV_X1    g457(.A(new_n628), .ZN(new_n659));
  INV_X1    g458(.A(new_n607), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n661), .A2(new_n594), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n501), .A3(new_n441), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT45), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n658), .B2(new_n659), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n493), .A2(KEYINPUT44), .A3(new_n628), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n594), .A4(new_n607), .ZN(new_n668));
  OAI21_X1  g467(.A(G29gat), .B1(new_n668), .B2(new_n448), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(G1328gat));
  NAND4_X1  g469(.A1(new_n661), .A2(new_n502), .A3(new_n381), .A4(new_n594), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT46), .Z(new_n672));
  OAI21_X1  g471(.A(G36gat), .B1(new_n668), .B2(new_n449), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(G1329gat));
  OAI21_X1  g473(.A(G43gat), .B1(new_n668), .B2(new_n647), .ZN(new_n675));
  INV_X1    g474(.A(G43gat), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n661), .A2(new_n676), .A3(new_n649), .A4(new_n594), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT47), .B1(new_n678), .B2(KEYINPUT104), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n680), .B(new_n681), .C1(new_n675), .C2(new_n677), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n679), .A2(new_n682), .ZN(G1330gat));
  INV_X1    g482(.A(G50gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n662), .A2(new_n684), .A3(new_n347), .ZN(new_n685));
  OAI21_X1  g484(.A(G50gat), .B1(new_n668), .B2(new_n486), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT48), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1331gat));
  INV_X1    g488(.A(new_n593), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n552), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n629), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT105), .Z(new_n693));
  AND2_X1   g492(.A1(new_n493), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n441), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n556), .ZN(G1332gat));
  AOI21_X1  g495(.A(new_n449), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT106), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(G1333gat));
  NAND4_X1  g500(.A1(new_n493), .A2(G71gat), .A3(new_n490), .A4(new_n693), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT107), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n694), .A2(new_n649), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(G71gat), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g505(.A1(new_n694), .A2(new_n347), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT109), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(G78gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1335gat));
  NAND4_X1  g509(.A1(new_n666), .A2(new_n667), .A3(new_n607), .A4(new_n691), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(new_n384), .A3(new_n448), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n493), .A2(new_n553), .A3(new_n628), .A4(new_n607), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n690), .B1(new_n713), .B2(KEYINPUT51), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n659), .B1(new_n462), .B2(new_n492), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n715), .A2(new_n716), .A3(new_n553), .A4(new_n607), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n441), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n712), .B1(new_n384), .B2(new_n718), .ZN(G1336gat));
  NAND4_X1  g518(.A1(new_n714), .A2(new_n570), .A3(new_n381), .A4(new_n717), .ZN(new_n720));
  OAI21_X1  g519(.A(G92gat), .B1(new_n711), .B2(new_n449), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT52), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1337gat));
  INV_X1    g526(.A(G99gat), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n711), .A2(new_n728), .A3(new_n647), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n649), .A3(new_n717), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(G1338gat));
  NAND2_X1  g530(.A1(new_n713), .A2(KEYINPUT51), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n732), .A2(new_n347), .A3(new_n593), .A4(new_n717), .ZN(new_n733));
  INV_X1    g532(.A(G106gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n711), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(G106gat), .A3(new_n347), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n735), .A2(new_n737), .A3(KEYINPUT53), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1339gat));
  OR3_X1    g541(.A1(new_n583), .A2(new_n554), .A3(new_n584), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(KEYINPUT54), .A3(new_n585), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT54), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n745), .B(new_n554), .C1(new_n583), .C2(new_n584), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n746), .A2(KEYINPUT111), .A3(new_n590), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT111), .B1(new_n746), .B2(new_n590), .ZN(new_n748));
  OAI211_X1 g547(.A(KEYINPUT55), .B(new_n744), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n591), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT112), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n752), .A3(new_n591), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n751), .A2(new_n552), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n551), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n759));
  INV_X1    g558(.A(new_n548), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n519), .A2(new_n536), .A3(new_n534), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT113), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n532), .A2(new_n519), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n520), .B2(new_n763), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n593), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n628), .B1(new_n757), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n760), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n628), .B(new_n769), .C1(new_n551), .C2(new_n550), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n607), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n629), .A2(new_n553), .A3(new_n690), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n448), .A2(new_n381), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(new_n777), .A3(new_n773), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n458), .A2(new_n775), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n243), .A3(new_n552), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n286), .A2(new_n347), .A3(new_n348), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n775), .A2(new_n781), .A3(new_n776), .A4(new_n778), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n783), .A2(new_n552), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n785), .B2(new_n243), .ZN(G1340gat));
  NAND3_X1  g585(.A1(new_n779), .A2(new_n241), .A3(new_n593), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n783), .A2(new_n593), .A3(new_n784), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n241), .ZN(G1341gat));
  NAND4_X1  g588(.A1(new_n783), .A2(G127gat), .A3(new_n660), .A4(new_n784), .ZN(new_n790));
  INV_X1    g589(.A(new_n779), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n250), .B1(new_n791), .B2(new_n607), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n790), .A2(new_n792), .ZN(G1342gat));
  NAND3_X1  g592(.A1(new_n783), .A2(new_n628), .A3(new_n784), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(G134gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n659), .A2(G134gat), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT56), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n775), .A2(new_n458), .A3(new_n778), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n776), .A4(new_n796), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n779), .A2(KEYINPUT116), .A3(new_n800), .A4(new_n796), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n798), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT117), .B1(new_n795), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n798), .A2(new_n803), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n794), .A2(G134gat), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n804), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n810), .ZN(G1343gat));
  AND2_X1   g610(.A1(new_n775), .A2(new_n778), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n347), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n647), .A2(new_n776), .ZN(new_n815));
  INV_X1    g614(.A(new_n773), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n750), .B1(new_n755), .B2(new_n754), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n817), .A2(new_n552), .B1(new_n765), .B2(new_n593), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n818), .A2(new_n628), .B1(new_n768), .B2(new_n770), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n819), .B2(new_n607), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(new_n486), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n815), .B1(new_n821), .B2(KEYINPUT57), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n814), .A2(new_n822), .A3(new_n552), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G141gat), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n812), .A2(new_n347), .ZN(new_n827));
  INV_X1    g626(.A(new_n815), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n316), .A3(new_n552), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(new_n830), .A3(KEYINPUT58), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n824), .B(new_n829), .C1(new_n825), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1344gat));
  OR2_X1    g633(.A1(new_n300), .A2(new_n301), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n814), .A2(new_n822), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT59), .B(new_n835), .C1(new_n836), .C2(new_n593), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n775), .A2(KEYINPUT57), .A3(new_n347), .A4(new_n778), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n813), .B1(new_n820), .B2(new_n486), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n593), .A3(new_n828), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(G148gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n593), .A2(new_n835), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n837), .A2(new_n843), .B1(new_n844), .B2(new_n845), .ZN(G1345gat));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n660), .A3(new_n828), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n660), .A2(G155gat), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT119), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n310), .A2(new_n847), .B1(new_n836), .B2(new_n849), .ZN(G1346gat));
  NAND3_X1  g649(.A1(new_n836), .A2(G162gat), .A3(new_n628), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n311), .B1(new_n844), .B2(new_n659), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(G1347gat));
  NOR2_X1   g652(.A1(new_n441), .A2(new_n449), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT121), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n812), .A2(KEYINPUT122), .A3(new_n781), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n775), .A2(new_n781), .A3(new_n778), .A4(new_n855), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n552), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G169gat), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n775), .A2(new_n458), .A3(new_n778), .A4(new_n854), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n553), .A2(G169gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n861), .B1(new_n866), .B2(new_n867), .ZN(G1348gat));
  NAND3_X1  g667(.A1(new_n856), .A2(new_n593), .A3(new_n859), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G176gat), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n690), .A2(G176gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n864), .B2(new_n865), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT123), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1349gat));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n660), .A3(new_n859), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G183gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n799), .A2(new_n204), .A3(new_n660), .A4(new_n854), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n882));
  NAND2_X1  g681(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1350gat));
  NAND3_X1  g684(.A1(new_n856), .A2(new_n628), .A3(new_n859), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(G190gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n886), .B2(G190gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n628), .A2(new_n205), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n888), .A2(new_n889), .B1(new_n866), .B2(new_n890), .ZN(G1351gat));
  AND4_X1   g690(.A1(new_n647), .A2(new_n812), .A3(new_n347), .A4(new_n854), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n545), .A3(new_n552), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n855), .A2(new_n647), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n839), .B2(new_n840), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n552), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n545), .B2(new_n896), .ZN(G1352gat));
  INV_X1    g696(.A(G204gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n898), .A3(new_n593), .ZN(new_n899));
  XOR2_X1   g698(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n690), .B(new_n894), .C1(new_n839), .C2(new_n840), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n902), .B(new_n903), .C1(new_n898), .C2(new_n904), .ZN(G1353gat));
  NAND3_X1  g704(.A1(new_n892), .A2(new_n289), .A3(new_n660), .ZN(new_n906));
  INV_X1    g705(.A(new_n894), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n841), .A2(new_n660), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n289), .B1(new_n908), .B2(KEYINPUT126), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n910), .A3(new_n660), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n909), .A2(KEYINPUT63), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(G1354gat));
  AOI21_X1  g713(.A(G218gat), .B1(new_n892), .B2(new_n628), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n628), .A2(G218gat), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT127), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n895), .B2(new_n917), .ZN(G1355gat));
endmodule


