//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n865, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  NOR3_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n203), .A2(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT92), .B(G29gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT93), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n205), .A2(KEYINPUT91), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n207), .B1(new_n205), .B2(KEYINPUT91), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(KEYINPUT15), .A3(new_n209), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(G1gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n222), .B2(KEYINPUT95), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n226), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT97), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n214), .A2(new_n218), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT17), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n219), .A2(KEYINPUT97), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT96), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n229), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n202), .B(new_n230), .C1(new_n236), .C2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n232), .A2(new_n231), .A3(KEYINPUT17), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT97), .B1(new_n219), .B2(new_n234), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n240), .A3(new_n238), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n248), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n230), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n219), .A2(new_n229), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT98), .A3(new_n230), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n202), .B(KEYINPUT13), .Z(new_n252));
  INV_X1    g051(.A(KEYINPUT98), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n219), .A2(new_n253), .A3(new_n229), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n244), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT11), .B(G169gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT12), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n244), .A2(new_n263), .A3(new_n249), .A4(new_n255), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266));
  INV_X1    g065(.A(G169gat), .ZN(new_n267));
  INV_X1    g066(.A(G176gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT26), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT27), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT27), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT70), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n284), .A2(KEYINPUT28), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n290));
  AOI21_X1  g089(.A(G190gat), .B1(new_n280), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n280), .B2(new_n282), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n278), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n277), .ZN(new_n298));
  NAND3_X1  g097(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n274), .A2(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n267), .A2(new_n268), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT64), .B(G169gat), .ZN(new_n304));
  OR2_X1    g103(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT23), .A3(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n300), .B(new_n303), .C1(new_n304), .C2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n296), .B1(new_n301), .B2(new_n302), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n269), .A2(KEYINPUT23), .A3(new_n271), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n299), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n299), .A2(new_n312), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n298), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n296), .A2(new_n308), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT73), .B1(new_n295), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G127gat), .ZN(new_n319));
  INV_X1    g118(.A(G127gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G134gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n325));
  INV_X1    g124(.A(G113gat), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G120gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT72), .B1(new_n328), .B2(G113gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n326), .A3(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n323), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n328), .A2(G113gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n326), .A2(G120gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n322), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n300), .A2(new_n303), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n307), .A2(new_n304), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n296), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n315), .A2(new_n310), .A3(new_n309), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n272), .A2(new_n275), .B1(G183gat), .B2(G190gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n287), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n286), .B1(new_n280), .B2(new_n282), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n285), .A2(KEYINPUT28), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n289), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(new_n291), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n345), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n317), .A2(new_n339), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n344), .A2(new_n353), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT71), .B(G120gat), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n329), .B(new_n331), .C1(new_n358), .C2(new_n326), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n359), .A2(new_n323), .B1(new_n336), .B2(new_n337), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(KEYINPUT73), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n356), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT33), .ZN(new_n365));
  XNOR2_X1  g164(.A(G15gat), .B(G43gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n364), .B(KEYINPUT32), .C1(new_n365), .C2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n364), .B2(KEYINPUT32), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n365), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n370), .A2(KEYINPUT74), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT74), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n361), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT34), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n362), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n375), .A2(KEYINPUT76), .A3(new_n376), .A4(new_n362), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n363), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n356), .A2(KEYINPUT75), .A3(new_n361), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n376), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n374), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n381), .A2(new_n385), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n371), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n370), .A2(KEYINPUT74), .A3(new_n371), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n393), .B2(new_n369), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT36), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n396));
  INV_X1    g195(.A(G162gat), .ZN(new_n397));
  OR2_X1    g196(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT2), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n399), .ZN(new_n403));
  NOR2_X1   g202(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n404));
  OAI21_X1  g203(.A(G162gat), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n406));
  XOR2_X1   g205(.A(G155gat), .B(G162gat), .Z(new_n407));
  XNOR2_X1  g206(.A(G141gat), .B(G148gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n402), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(new_n408), .B2(KEYINPUT2), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n360), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n360), .A2(new_n410), .A3(new_n415), .A4(new_n411), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n410), .A2(new_n411), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n339), .A2(KEYINPUT80), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n333), .A2(new_n421), .A3(new_n338), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n410), .A2(new_n423), .A3(new_n411), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n419), .A2(new_n420), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n412), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n417), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT82), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n412), .ZN(new_n431));
  INV_X1    g230(.A(new_n426), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g232(.A(KEYINPUT82), .B(new_n426), .C1(new_n430), .C2(new_n412), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n428), .B(KEYINPUT5), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT0), .ZN(new_n438));
  XNOR2_X1  g237(.A(G57gat), .B(G85gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n413), .A2(new_n416), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT5), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n425), .A2(new_n442), .A3(new_n443), .A4(new_n426), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n435), .A2(new_n436), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n435), .A2(new_n444), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n440), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT77), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n295), .B2(new_n316), .ZN(new_n453));
  XNOR2_X1  g252(.A(G197gat), .B(G204gat), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT22), .ZN(new_n455));
  INV_X1    g254(.A(G211gat), .ZN(new_n456));
  INV_X1    g255(.A(G218gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G211gat), .B(G218gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT29), .B1(new_n344), .B2(new_n353), .ZN(new_n463));
  INV_X1    g262(.A(new_n451), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n453), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G64gat), .B(G92gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n466), .B(new_n467), .Z(new_n468));
  AOI21_X1  g267(.A(new_n451), .B1(new_n344), .B2(new_n353), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT29), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n295), .B2(new_n316), .ZN(new_n471));
  INV_X1    g270(.A(new_n452), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n465), .B(new_n468), .C1(new_n473), .C2(new_n462), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n465), .B1(new_n473), .B2(new_n462), .ZN(new_n477));
  INV_X1    g276(.A(new_n468), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n452), .B1(new_n357), .B2(new_n470), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n461), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n481), .A2(KEYINPUT30), .A3(new_n468), .A4(new_n465), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n476), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n441), .B1(new_n435), .B2(new_n444), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n435), .A2(new_n441), .A3(new_n444), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(KEYINPUT83), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n450), .B(new_n484), .C1(new_n487), .C2(KEYINPUT6), .ZN(new_n488));
  INV_X1    g287(.A(new_n418), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n462), .A2(new_n470), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(new_n423), .ZN(new_n491));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n462), .B1(new_n424), .B2(new_n470), .ZN(new_n493));
  OR3_X1    g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n460), .A2(new_n454), .A3(new_n458), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT29), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n462), .B2(new_n496), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n489), .B1(new_n498), .B2(new_n423), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n492), .B1(new_n499), .B2(new_n493), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G22gat), .ZN(new_n502));
  INV_X1    g301(.A(G22gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT31), .B(G50gat), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT84), .ZN(new_n506));
  XOR2_X1   g305(.A(G78gat), .B(G106gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n502), .A2(KEYINPUT86), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n512), .A2(new_n508), .B1(new_n502), .B2(new_n504), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n488), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n374), .A2(new_n386), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n393), .A2(new_n388), .A3(new_n369), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n395), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n512), .A2(new_n508), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n504), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n509), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n425), .A2(new_n442), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n432), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n430), .A2(new_n426), .A3(new_n412), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT87), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n430), .A2(new_n529), .A3(new_n426), .A4(new_n412), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n526), .A2(new_n531), .A3(KEYINPUT39), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n426), .B1(new_n425), .B2(new_n442), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n440), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT40), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n449), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(KEYINPUT40), .A3(new_n535), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n483), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n483), .A2(new_n541), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT40), .B1(new_n532), .B2(new_n535), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n485), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT88), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n524), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n445), .A2(new_n446), .B1(new_n448), .B2(new_n440), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n449), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n551), .B2(new_n446), .ZN(new_n552));
  INV_X1    g351(.A(new_n474), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n473), .A2(new_n461), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n453), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT38), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n468), .A2(new_n555), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(new_n477), .B2(new_n478), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n553), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT89), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n555), .B1(new_n481), .B2(new_n465), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n563), .B(KEYINPUT38), .C1(new_n560), .C2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n477), .A2(KEYINPUT37), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n468), .B1(new_n481), .B2(new_n465), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(new_n559), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n563), .B1(new_n569), .B2(KEYINPUT38), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n562), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n552), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT90), .B1(new_n548), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n540), .B1(new_n539), .B2(new_n542), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n544), .A2(new_n546), .A3(KEYINPUT88), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n514), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(KEYINPUT38), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT89), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n565), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT6), .B1(new_n550), .B2(new_n449), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n579), .B(new_n562), .C1(new_n580), .C2(new_n549), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n520), .B1(new_n573), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n516), .A2(new_n517), .A3(new_n524), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586));
  INV_X1    g385(.A(new_n488), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n516), .A2(new_n517), .A3(new_n524), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT35), .B1(new_n589), .B2(new_n488), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n265), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT99), .ZN(new_n593));
  AND2_X1   g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT103), .Z(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(KEYINPUT8), .A2(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G99gat), .B(G106gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT104), .Z(new_n608));
  NAND3_X1  g407(.A1(new_n247), .A2(new_n240), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n219), .A2(new_n607), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT105), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n613), .A2(new_n614), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n598), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n613), .A3(new_n597), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT100), .B1(G71gat), .B2(G78gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G57gat), .B(G64gat), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G71gat), .B(G78gat), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n627), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT101), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n627), .B(new_n628), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(KEYINPUT21), .ZN(new_n636));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n229), .B1(new_n635), .B2(KEYINPUT21), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT102), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n640), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n623), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT106), .B(KEYINPUT10), .Z(new_n649));
  INV_X1    g448(.A(new_n607), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n607), .A2(new_n630), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT107), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n653), .B2(new_n655), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n658), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n651), .A2(new_n652), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n666), .B(KEYINPUT108), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n656), .A2(new_n662), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(new_n663), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n648), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n593), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n552), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g476(.A1(new_n593), .A2(new_n483), .A3(new_n674), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(G8gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT42), .B2(new_n681), .ZN(G1325gat));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n518), .B1(new_n516), .B2(new_n517), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n395), .A2(KEYINPUT109), .A3(new_n519), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n675), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n387), .A2(new_n394), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n690), .B1(new_n675), .B2(new_n693), .ZN(G1326gat));
  NAND3_X1  g493(.A1(new_n593), .A2(new_n514), .A3(new_n674), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  XOR2_X1   g496(.A(new_n673), .B(KEYINPUT110), .Z(new_n698));
  INV_X1    g497(.A(new_n647), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n265), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n395), .A2(new_n515), .A3(new_n519), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n582), .B1(new_n576), .B2(new_n581), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n588), .A2(new_n590), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n623), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n701), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n622), .B1(new_n584), .B2(new_n591), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n515), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n573), .B2(new_n583), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n591), .B1(new_n714), .B2(new_n689), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n623), .A2(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n700), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n211), .B1(new_n720), .B2(new_n552), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n622), .A2(new_n699), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n673), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n593), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n552), .A2(new_n211), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n722), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n593), .A2(new_n724), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(KEYINPUT45), .A3(new_n726), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n721), .A2(new_n728), .A3(new_n730), .ZN(G1328gat));
  OAI21_X1  g530(.A(G36gat), .B1(new_n720), .B2(new_n484), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n484), .A2(G36gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT46), .B1(new_n725), .B2(new_n734), .ZN(new_n735));
  OR3_X1    g534(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n734), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n735), .A3(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n725), .B2(new_n692), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n709), .A2(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n689), .A2(new_n738), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n741), .A2(new_n700), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT47), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n739), .B(new_n746), .C1(new_n720), .C2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1330gat));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  INV_X1    g548(.A(G50gat), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n719), .B2(new_n514), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n725), .A2(G50gat), .A3(new_n524), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n729), .A2(new_n750), .A3(new_n514), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n741), .A2(new_n524), .A3(new_n700), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n754), .B(KEYINPUT48), .C1(new_n755), .C2(new_n750), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(G1331gat));
  NAND2_X1  g556(.A1(new_n573), .A2(new_n583), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n689), .A3(new_n515), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n265), .B1(new_n759), .B2(new_n706), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n648), .A2(new_n698), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n552), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g565(.A(new_n484), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n768), .A2(KEYINPUT112), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(KEYINPUT112), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1333gat));
  INV_X1    g573(.A(G71gat), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n689), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT113), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n691), .B(KEYINPUT114), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n762), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n763), .A2(new_n514), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  INV_X1    g584(.A(new_n723), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n760), .A2(new_n786), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n760), .A2(new_n792), .A3(KEYINPUT51), .A4(new_n786), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n794), .A2(new_n602), .A3(new_n764), .A4(new_n673), .ZN(new_n795));
  INV_X1    g594(.A(new_n265), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n699), .A3(new_n673), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n741), .A2(new_n552), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n795), .B1(new_n800), .B2(new_n801), .ZN(G1336gat));
  NOR3_X1   g601(.A1(new_n698), .A2(G92gat), .A3(new_n484), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n741), .A2(new_n484), .A3(new_n797), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n603), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n797), .B1(new_n712), .B2(new_n718), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n483), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n787), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n809), .A2(G92gat), .B1(new_n810), .B2(new_n803), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n805), .ZN(G1337gat));
  INV_X1    g611(.A(G99gat), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n794), .A2(new_n813), .A3(new_n691), .A4(new_n673), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n741), .A2(new_n689), .A3(new_n797), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n813), .ZN(G1338gat));
  NOR3_X1   g615(.A1(new_n698), .A2(G106gat), .A3(new_n524), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n760), .B2(new_n786), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n715), .A2(new_n790), .A3(new_n265), .A4(new_n723), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT117), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(G106gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n808), .B2(new_n514), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT53), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n794), .A2(new_n817), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n741), .A2(new_n524), .A3(new_n797), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n825), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(G1339gat));
  NOR4_X1   g631(.A1(new_n622), .A2(new_n265), .A3(new_n699), .A4(new_n673), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n202), .B1(new_n248), .B2(new_n230), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n252), .B1(new_n251), .B2(new_n254), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n260), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n264), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n658), .C1(new_n653), .C2(new_n655), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n667), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n656), .B2(new_n662), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n661), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n842), .A2(KEYINPUT55), .B1(new_n661), .B2(new_n668), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n622), .A2(new_n837), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n264), .A2(new_n673), .A3(new_n836), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n262), .B2(new_n264), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n843), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n849), .B2(new_n622), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n833), .B1(new_n850), .B2(new_n699), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n589), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n552), .A2(new_n483), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n265), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n326), .A2(KEYINPUT118), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n326), .A2(KEYINPUT118), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n854), .B2(new_n698), .ZN(new_n861));
  INV_X1    g660(.A(new_n358), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n673), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n854), .B2(new_n863), .ZN(G1341gat));
  NOR2_X1   g663(.A1(new_n854), .A2(new_n699), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(new_n320), .ZN(G1342gat));
  NOR2_X1   g665(.A1(new_n623), .A2(new_n483), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n318), .A3(new_n764), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT56), .Z(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n854), .B2(new_n623), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  INV_X1    g670(.A(new_n851), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n764), .A3(new_n514), .A4(new_n689), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n483), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n796), .A2(G141gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT57), .B1(new_n851), .B2(new_n524), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(new_n255), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n242), .B2(new_n243), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n263), .B1(new_n880), .B2(new_n249), .ZN(new_n881));
  INV_X1    g680(.A(new_n264), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n845), .B(new_n843), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n847), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n623), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n647), .B1(new_n886), .B2(new_n846), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n878), .B(new_n514), .C1(new_n887), .C2(new_n833), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n689), .A2(new_n853), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n877), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G141gat), .B1(new_n890), .B2(new_n796), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g692(.A(G148gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n874), .A2(new_n894), .A3(new_n673), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n888), .A3(new_n673), .A4(new_n889), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(G148gat), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n896), .B2(G148gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(G1345gat));
  NAND4_X1  g699(.A1(new_n874), .A2(new_n398), .A3(new_n399), .A4(new_n647), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n890), .A2(new_n699), .B1(new_n404), .B2(new_n403), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1346gat));
  OAI21_X1  g702(.A(G162gat), .B1(new_n890), .B2(new_n623), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n867), .A2(new_n397), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n873), .B2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n764), .A2(new_n484), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n780), .A2(new_n514), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n872), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n796), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n852), .A2(new_n907), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(KEYINPUT119), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n796), .A2(new_n304), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n673), .A3(new_n915), .ZN(new_n919));
  INV_X1    g718(.A(new_n910), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n698), .B1(new_n305), .B2(new_n306), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n919), .A2(new_n268), .B1(new_n920), .B2(new_n921), .ZN(G1349gat));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n923), .A3(new_n647), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT120), .B1(new_n910), .B2(new_n699), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(G183gat), .A3(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n699), .A2(new_n347), .A3(new_n346), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n913), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n926), .B2(new_n929), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(G1350gat));
  NAND2_X1  g732(.A1(new_n622), .A2(new_n285), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n920), .A2(new_n622), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(G190gat), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n935), .B2(G190gat), .ZN(new_n938));
  OAI22_X1  g737(.A1(new_n916), .A2(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  NAND2_X1  g738(.A1(new_n877), .A2(new_n888), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT124), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n877), .A2(new_n888), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n908), .B1(new_n688), .B2(new_n687), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n265), .A2(G197gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n908), .A2(new_n524), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n872), .A2(new_n689), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n265), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n947), .A2(new_n950), .ZN(G1352gat));
  INV_X1    g750(.A(G204gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n952), .A3(new_n673), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT62), .Z(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n945), .B2(new_n698), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n949), .A2(new_n456), .A3(new_n647), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n944), .A2(new_n647), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n877), .A2(new_n888), .A3(new_n958), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g763(.A(KEYINPUT125), .B(new_n957), .C1(new_n960), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1354gat));
  AOI21_X1  g765(.A(G218gat), .B1(new_n949), .B2(new_n622), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n945), .A2(new_n457), .A3(new_n623), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(G1355gat));
endmodule


