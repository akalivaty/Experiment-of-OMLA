//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1047, new_n1048;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n208));
  NOR2_X1   g007(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(KEYINPUT76), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n218), .A3(G148gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n219), .A2(new_n204), .ZN(new_n220));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n214), .B(new_n215), .C1(new_n220), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G197gat), .B(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G211gat), .A2(G218gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT22), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n229), .A3(new_n232), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(KEYINPUT71), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n228), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n214), .B1(new_n220), .B2(new_n225), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT29), .B1(new_n236), .B2(new_n237), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G228gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n243), .B(KEYINPUT81), .C1(new_n244), .C2(KEYINPUT3), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n242), .A2(new_n247), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G22gat), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n219), .A2(new_n204), .B1(new_n224), .B2(new_n223), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n212), .B1(new_n207), .B2(new_n210), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT29), .B1(new_n256), .B2(new_n215), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n245), .B1(new_n257), .B2(new_n239), .ZN(new_n258));
  NAND2_X1  g057(.A1(G228gat), .A2(G233gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n252), .A2(new_n253), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n253), .B1(new_n252), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g061(.A(G78gat), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n252), .A2(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G22gat), .ZN(new_n265));
  INV_X1    g064(.A(G78gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n252), .A2(new_n253), .A3(new_n260), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT31), .B(G50gat), .ZN(new_n269));
  INV_X1    g068(.A(G106gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n263), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n263), .B2(new_n268), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT82), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n271), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n261), .A2(new_n262), .A3(G78gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n268), .A3(new_n271), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT82), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT79), .ZN(new_n284));
  XOR2_X1   g083(.A(G1gat), .B(G29gat), .Z(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G225gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G113gat), .ZN(new_n293));
  INV_X1    g092(.A(G113gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G120gat), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT1), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G127gat), .A2(G134gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(G127gat), .A2(G134gat), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT68), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301));
  INV_X1    g100(.A(G127gat), .ZN(new_n302));
  INV_X1    g101(.A(G134gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n304), .B2(new_n297), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n296), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT69), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n297), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n296), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n310), .B(new_n296), .C1(new_n300), .C2(new_n305), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n307), .A2(new_n256), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n311), .A2(new_n309), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n315), .A2(KEYINPUT4), .A3(new_n307), .A4(new_n256), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(new_n254), .B2(new_n255), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n309), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT68), .B1(new_n298), .B2(new_n299), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n301), .A3(new_n297), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n310), .B1(new_n321), .B2(new_n296), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n226), .B(new_n317), .C1(new_n318), .C2(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n314), .A2(new_n316), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n243), .B1(new_n318), .B2(new_n322), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n312), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n291), .ZN(new_n328));
  OAI211_X1 g127(.A(KEYINPUT77), .B(new_n243), .C1(new_n318), .C2(new_n322), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n291), .A2(new_n324), .B1(new_n330), .B2(KEYINPUT5), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n291), .A4(new_n323), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n284), .B(new_n290), .C1(new_n331), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT6), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(KEYINPUT5), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n332), .ZN(new_n339));
  INV_X1    g138(.A(new_n334), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n284), .B1(new_n341), .B2(new_n290), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n283), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n290), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n334), .B1(new_n332), .B2(new_n338), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT79), .B1(new_n346), .B2(new_n289), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n347), .A2(KEYINPUT80), .A3(new_n336), .A4(new_n335), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n345), .A2(new_n336), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n241), .A2(new_n238), .ZN(new_n357));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT27), .B(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(KEYINPUT28), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G183gat), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT27), .B1(new_n363), .B2(KEYINPUT67), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n366), .A3(G183gat), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n364), .A2(new_n367), .A3(new_n361), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n368), .B2(KEYINPUT28), .ZN(new_n369));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n371), .A2(KEYINPUT26), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n371), .B1(KEYINPUT23), .B2(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(KEYINPUT23), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT66), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT66), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n371), .A2(new_n382), .A3(KEYINPUT23), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n379), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT65), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT65), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n387), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n370), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT25), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n385), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n375), .A2(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n394), .A2(KEYINPUT25), .A3(new_n396), .A4(new_n380), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n378), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n359), .B1(new_n399), .B2(new_n227), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401));
  INV_X1    g200(.A(G169gat), .ZN(new_n402));
  INV_X1    g201(.A(G176gat), .ZN(new_n403));
  AND4_X1   g202(.A1(new_n382), .A2(new_n402), .A3(new_n403), .A4(KEYINPUT23), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n382), .B1(new_n371), .B2(KEYINPUT23), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n396), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n386), .A2(new_n388), .B1(new_n370), .B2(new_n390), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n401), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n408), .A2(new_n397), .B1(new_n369), .B2(new_n377), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(new_n358), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT72), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n358), .B1(new_n409), .B2(KEYINPUT29), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n357), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n359), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n412), .A2(new_n239), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n356), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n357), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n413), .B1(new_n412), .B2(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n227), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT72), .B1(new_n421), .B2(new_n358), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n417), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n424), .A4(new_n355), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT73), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n418), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n414), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n417), .B1(new_n428), .B2(new_n419), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(KEYINPUT73), .A3(KEYINPUT30), .A4(new_n355), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n427), .A2(KEYINPUT74), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT74), .B1(new_n427), .B2(new_n430), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n355), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n431), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n282), .B1(new_n352), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n318), .A2(new_n322), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n409), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT70), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n399), .B1(new_n322), .B2(new_n318), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n446), .B(KEYINPUT64), .Z(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n409), .A2(new_n440), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n444), .A2(new_n445), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(new_n450), .A3(new_n443), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT34), .B1(new_n452), .B2(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT33), .B1(new_n452), .B2(new_n447), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n452), .A2(new_n447), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n451), .B(new_n453), .C1(new_n455), .C2(new_n458), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n460), .B2(new_n464), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n439), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT36), .A3(new_n465), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n202), .B1(new_n438), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n275), .A2(new_n281), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n347), .A2(new_n336), .A3(new_n335), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n344), .B1(new_n474), .B2(new_n283), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n350), .B1(new_n475), .B2(new_n348), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n427), .A2(new_n430), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n427), .A2(KEYINPUT74), .A3(new_n430), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n435), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n473), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n468), .A2(new_n470), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(KEYINPUT83), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n356), .B1(new_n429), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n356), .C1(new_n429), .C2(new_n485), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT86), .B(KEYINPUT37), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n429), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n474), .A2(new_n344), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n355), .B(new_n494), .C1(new_n429), .C2(new_n490), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n428), .A2(new_n419), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n239), .B1(new_n412), .B2(new_n416), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT37), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n497), .A2(new_n500), .B1(new_n429), .B2(new_n355), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n495), .A2(new_n351), .A3(new_n496), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n272), .A2(new_n273), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT84), .B1(new_n324), .B2(new_n291), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n314), .A2(new_n316), .A3(new_n323), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n328), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT39), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n327), .A2(new_n329), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(new_n291), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n505), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n514), .A3(new_n290), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT40), .A4(new_n290), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n517), .A2(new_n345), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n477), .A2(new_n435), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n504), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n472), .A2(new_n484), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n496), .A2(new_n351), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n466), .A2(new_n467), .ZN(new_n526));
  INV_X1    g325(.A(new_n520), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n469), .A2(new_n503), .A3(new_n465), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n476), .A2(new_n481), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G50gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G43gat), .ZN(new_n535));
  INV_X1    g334(.A(G43gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G50gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n537), .A3(KEYINPUT89), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT15), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(G29gat), .ZN(new_n545));
  INV_X1    g344(.A(G36gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT90), .ZN(new_n548));
  NOR3_X1   g347(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n543), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n552), .A2(new_n553), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n543), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n547), .A2(KEYINPUT90), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n549), .A2(new_n550), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT91), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n542), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n537), .A2(KEYINPUT92), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n535), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n537), .A2(KEYINPUT92), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n547), .A2(new_n543), .B1(G29gat), .B2(G36gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n542), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT17), .B1(new_n560), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n542), .ZN(new_n570));
  INV_X1    g369(.A(new_n559), .ZN(new_n571));
  NAND2_X1  g370(.A1(G29gat), .A2(G36gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n558), .B2(KEYINPUT91), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n567), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT16), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(G1gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(G1gat), .B2(new_n578), .ZN(new_n581));
  INV_X1    g380(.A(G8gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n567), .ZN(new_n585));
  INV_X1    g384(.A(new_n583), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n585), .A2(new_n586), .B1(G229gat), .B2(G233gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(KEYINPUT18), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n586), .B1(new_n569), .B2(new_n576), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n585), .A2(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n589), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n594), .B(KEYINPUT13), .Z(new_n597));
  INV_X1    g396(.A(new_n593), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n585), .A2(new_n586), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n591), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G197gat), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT11), .B(G169gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n591), .A2(new_n596), .A3(new_n607), .A4(new_n600), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT94), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n601), .A2(new_n612), .A3(new_n608), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n611), .A2(KEYINPUT95), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT95), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G85gat), .A2(G92gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT7), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G99gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n270), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n619), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n618), .A2(new_n627), .A3(new_n622), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n585), .A2(new_n629), .B1(KEYINPUT41), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n626), .A2(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n577), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n640), .B(new_n632), .C1(new_n635), .C2(new_n636), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(KEYINPUT103), .A3(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n637), .A2(KEYINPUT103), .A3(new_n638), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n631), .A2(KEYINPUT41), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT101), .Z(new_n645));
  XNOR2_X1  g444(.A(G134gat), .B(G162gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G57gat), .B(G64gat), .Z(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(KEYINPUT96), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT9), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n650), .B2(KEYINPUT96), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G71gat), .B(G78gat), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT97), .ZN(new_n658));
  INV_X1    g457(.A(new_n655), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n650), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n656), .A2(KEYINPUT100), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n651), .B2(new_n653), .ZN(new_n663));
  INV_X1    g462(.A(new_n660), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n665), .A3(KEYINPUT21), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n583), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n656), .A2(new_n660), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT98), .B(KEYINPUT21), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G231gat), .A2(G233gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G127gat), .B(G155gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(G183gat), .B(G211gat), .Z(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n677), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n679), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n670), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n679), .A2(new_n682), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n680), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n669), .A3(new_n683), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n632), .ZN(new_n691));
  INV_X1    g490(.A(new_n636), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT104), .B1(new_n694), .B2(new_n640), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n637), .A2(new_n696), .A3(new_n638), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n695), .A2(new_n697), .A3(new_n647), .A4(new_n641), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n649), .A2(new_n690), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT105), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n649), .A2(new_n698), .A3(new_n690), .A4(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(G230gat), .A2(G233gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n671), .A2(new_n633), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT10), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n629), .A2(new_n656), .A3(new_n660), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n633), .A2(new_n706), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n661), .A2(new_n709), .A3(new_n665), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n661), .A2(new_n709), .A3(new_n665), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n713), .A2(KEYINPUT106), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n704), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n705), .A2(new_n707), .ZN(new_n716));
  INV_X1    g515(.A(new_n704), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(G120gat), .B(G148gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT107), .ZN(new_n721));
  XNOR2_X1  g520(.A(G176gat), .B(G204gat), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n721), .B(new_n722), .Z(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n715), .A2(new_n718), .A3(new_n723), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n703), .A2(new_n727), .ZN(new_n728));
  AND4_X1   g527(.A1(KEYINPUT108), .A2(new_n533), .A3(new_n616), .A4(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n616), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n523), .B2(new_n532), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT108), .B1(new_n731), .B2(new_n728), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n352), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT109), .B(G1gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1324gat));
  XOR2_X1   g535(.A(KEYINPUT16), .B(G8gat), .Z(new_n737));
  OAI211_X1 g536(.A(new_n520), .B(new_n737), .C1(new_n729), .C2(new_n732), .ZN(new_n738));
  INV_X1    g537(.A(new_n732), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(KEYINPUT108), .A3(new_n728), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n527), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n738), .B1(new_n741), .B2(new_n582), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1325gat));
  XNOR2_X1  g545(.A(new_n483), .B(KEYINPUT110), .ZN(new_n747));
  OAI21_X1  g546(.A(G15gat), .B1(new_n733), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n526), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n749), .A2(G15gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n733), .B2(new_n750), .ZN(G1326gat));
  OAI21_X1  g550(.A(new_n473), .B1(new_n729), .B2(new_n732), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(KEYINPUT111), .B(new_n473), .C1(new_n729), .C2(new_n732), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT43), .B(G22gat), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n754), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1327gat));
  INV_X1    g558(.A(new_n727), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n690), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n611), .A2(new_n613), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n611), .A2(KEYINPUT112), .A3(new_n613), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT113), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n522), .A2(new_n482), .A3(new_n483), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n532), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n649), .A2(new_n698), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n771), .A2(KEYINPUT114), .A3(new_n772), .A4(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n533), .A2(new_n773), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n769), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n545), .B1(new_n781), .B2(new_n476), .ZN(new_n782));
  INV_X1    g581(.A(new_n773), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n762), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n731), .A2(new_n545), .A3(new_n476), .A4(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n785), .B(KEYINPUT45), .ZN(new_n790));
  AOI211_X1 g589(.A(new_n352), .B(new_n769), .C1(new_n778), .C2(new_n780), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n545), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(G1328gat));
  AOI21_X1  g592(.A(new_n546), .B1(new_n781), .B2(new_n520), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n731), .A2(new_n546), .A3(new_n520), .A4(new_n784), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT46), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT116), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n795), .B(new_n799), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n527), .B(new_n769), .C1(new_n778), .C2(new_n780), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n798), .B(new_n800), .C1(new_n801), .C2(new_n546), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n797), .A2(new_n802), .ZN(G1329gat));
  AND4_X1   g602(.A1(new_n536), .A2(new_n731), .A3(new_n526), .A4(new_n784), .ZN(new_n804));
  INV_X1    g603(.A(new_n747), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(G43gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n536), .B1(new_n781), .B2(new_n471), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n807), .A2(KEYINPUT47), .B1(new_n808), .B2(new_n810), .ZN(G1330gat));
  AND4_X1   g610(.A1(new_n534), .A2(new_n731), .A3(new_n473), .A4(new_n784), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n781), .A2(new_n473), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(G50gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n534), .B1(new_n781), .B2(new_n504), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT48), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n818), .ZN(G1331gat));
  AND3_X1   g618(.A1(new_n703), .A2(new_n760), .A3(new_n767), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n771), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n476), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g623(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n520), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT118), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n821), .A2(KEYINPUT119), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT119), .B1(new_n821), .B2(new_n827), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n830), .B(new_n831), .ZN(G1333gat));
  OAI21_X1  g631(.A(G71gat), .B1(new_n821), .B2(new_n747), .ZN(new_n833));
  INV_X1    g632(.A(G71gat), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n526), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT120), .B(KEYINPUT50), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n836), .B(new_n837), .Z(G1334gat));
  NOR2_X1   g637(.A1(new_n821), .A2(new_n282), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(new_n266), .ZN(G1335gat));
  INV_X1    g639(.A(new_n690), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n767), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n760), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n778), .B2(new_n780), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G85gat), .B1(new_n846), .B2(new_n352), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n783), .B1(new_n532), .B2(new_n770), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n848), .A2(KEYINPUT51), .A3(new_n843), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT51), .B1(new_n848), .B2(new_n843), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n760), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n476), .A2(new_n620), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(G1336gat));
  AOI21_X1  g652(.A(new_n621), .B1(new_n845), .B2(new_n520), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n527), .A2(G92gat), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT52), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n857), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n527), .B(new_n844), .C1(new_n778), .C2(new_n780), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n621), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(G1337gat));
  OAI21_X1  g662(.A(G99gat), .B1(new_n846), .B2(new_n747), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n526), .A2(new_n624), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n851), .B2(new_n865), .ZN(G1338gat));
  NOR2_X1   g665(.A1(new_n503), .A2(G106gat), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n473), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(G106gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n270), .B1(new_n845), .B2(new_n504), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n851), .B2(new_n868), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n871), .A2(new_n872), .B1(new_n873), .B2(new_n874), .ZN(G1339gat));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n713), .A2(KEYINPUT106), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n877), .A2(new_n717), .A3(new_n708), .A4(new_n711), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n715), .A2(KEYINPUT54), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n881), .B(new_n704), .C1(new_n712), .C2(new_n714), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n724), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n876), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n879), .A2(KEYINPUT55), .A3(new_n724), .A4(new_n882), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n884), .A2(new_n726), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n765), .A2(new_n766), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n594), .B1(new_n584), .B2(new_n593), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n598), .A2(new_n599), .A3(new_n597), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n605), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n610), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n727), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n773), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n884), .A2(new_n726), .A3(new_n885), .ZN(new_n895));
  AOI211_X1 g694(.A(new_n891), .B(new_n895), .C1(new_n649), .C2(new_n698), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n841), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n700), .A2(new_n702), .A3(new_n727), .A4(new_n767), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n473), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n900), .A2(new_n476), .A3(new_n526), .A4(new_n527), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n294), .A3(new_n730), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n899), .A2(new_n352), .A3(new_n529), .ZN(new_n903));
  INV_X1    g702(.A(new_n767), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n527), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n294), .B2(new_n905), .ZN(G1340gat));
  NOR3_X1   g705(.A1(new_n901), .A2(new_n292), .A3(new_n727), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n527), .A3(new_n760), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n292), .B2(new_n908), .ZN(G1341gat));
  OAI21_X1  g708(.A(G127gat), .B1(new_n901), .B2(new_n841), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n903), .A2(new_n302), .A3(new_n527), .A4(new_n690), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1342gat));
  NOR2_X1   g711(.A1(new_n783), .A2(new_n520), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n903), .A2(new_n303), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g714(.A(G134gat), .B1(new_n901), .B2(new_n783), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G1343gat));
  AND2_X1   g717(.A1(new_n216), .A2(new_n218), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n614), .A2(new_n615), .A3(new_n895), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n783), .B1(new_n921), .B2(new_n892), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n773), .A2(new_n610), .A3(new_n886), .A4(new_n890), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n690), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND4_X1   g723(.A1(new_n700), .A2(new_n702), .A3(new_n727), .A4(new_n767), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n473), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT57), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n897), .A2(new_n898), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n504), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n471), .A2(new_n352), .A3(new_n520), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n920), .B1(new_n932), .B2(new_n730), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT58), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n352), .B1(new_n897), .B2(new_n898), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n805), .A2(new_n503), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n616), .A2(new_n205), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT121), .ZN(new_n938));
  AND4_X1   g737(.A1(new_n527), .A2(new_n935), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n933), .A2(new_n934), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT95), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n763), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n611), .A2(KEYINPUT95), .A3(new_n613), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n945), .A3(new_n886), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n773), .B1(new_n946), .B2(new_n893), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n841), .B1(new_n947), .B2(new_n896), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n282), .B1(new_n948), .B2(new_n898), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n931), .B1(new_n949), .B2(new_n929), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT57), .B(new_n503), .C1(new_n897), .C2(new_n898), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n950), .A2(new_n767), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n940), .B1(new_n952), .B2(new_n919), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n942), .B1(new_n953), .B2(KEYINPUT58), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n927), .A2(new_n904), .A3(new_n930), .A4(new_n931), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n939), .B1(new_n955), .B2(new_n920), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(KEYINPUT122), .A3(new_n934), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n941), .B1(new_n954), .B2(new_n957), .ZN(G1344gat));
  INV_X1    g757(.A(KEYINPUT59), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n959), .B(G148gat), .C1(new_n932), .C2(new_n727), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n931), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n931), .A2(new_n962), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n963), .A2(new_n964), .A3(new_n727), .ZN(new_n965));
  AND4_X1   g764(.A1(new_n730), .A2(new_n700), .A3(new_n702), .A4(new_n727), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n929), .B(new_n473), .C1(new_n924), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n503), .B1(new_n897), .B2(new_n898), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n965), .B(new_n967), .C1(new_n929), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G148gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n961), .B1(new_n970), .B2(KEYINPUT59), .ZN(new_n971));
  AOI211_X1 g770(.A(KEYINPUT124), .B(new_n959), .C1(new_n969), .C2(G148gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n960), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n935), .A2(new_n936), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n974), .A2(new_n520), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(new_n203), .A3(new_n760), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(G1345gat));
  OAI21_X1  g776(.A(G155gat), .B1(new_n932), .B2(new_n841), .ZN(new_n978));
  INV_X1    g777(.A(G155gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n975), .A2(new_n979), .A3(new_n690), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1346gat));
  OAI21_X1  g780(.A(G162gat), .B1(new_n932), .B2(new_n783), .ZN(new_n982));
  INV_X1    g781(.A(G162gat), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n913), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n982), .B1(new_n974), .B2(new_n984), .ZN(G1347gat));
  NOR3_X1   g784(.A1(new_n476), .A2(new_n749), .A3(new_n527), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n900), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n987), .A2(new_n402), .A3(new_n730), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n476), .B1(new_n897), .B2(new_n898), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n520), .B1(new_n989), .B2(new_n990), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(new_n529), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n994), .A2(new_n995), .A3(new_n904), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n988), .B1(new_n996), .B2(new_n402), .ZN(G1348gat));
  OAI21_X1  g796(.A(G176gat), .B1(new_n987), .B2(new_n727), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n994), .A2(new_n995), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n760), .A2(new_n403), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(G1349gat));
  OAI21_X1  g800(.A(G183gat), .B1(new_n987), .B2(new_n841), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n690), .A2(new_n360), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1002), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(KEYINPUT60), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT60), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n1006), .B(new_n1002), .C1(new_n999), .C2(new_n1003), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1005), .A2(new_n1007), .ZN(G1350gat));
  NAND3_X1  g807(.A1(new_n900), .A2(new_n773), .A3(new_n986), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1009), .A2(new_n1010), .A3(G190gat), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1010), .B1(new_n1009), .B2(G190gat), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n773), .A2(new_n361), .ZN(new_n1013));
  OAI22_X1  g812(.A1(new_n1011), .A2(new_n1012), .B1(new_n999), .B2(new_n1013), .ZN(G1351gat));
  NAND3_X1  g813(.A1(new_n747), .A2(new_n352), .A3(new_n520), .ZN(new_n1015));
  INV_X1    g814(.A(new_n1015), .ZN(new_n1016));
  OAI211_X1 g815(.A(new_n967), .B(new_n1016), .C1(new_n929), .C2(new_n968), .ZN(new_n1017));
  INV_X1    g816(.A(G197gat), .ZN(new_n1018));
  NOR3_X1   g817(.A1(new_n1017), .A2(new_n1018), .A3(new_n730), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n994), .A2(new_n904), .A3(new_n936), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1019), .B1(new_n1020), .B2(new_n1018), .ZN(G1352gat));
  NOR2_X1   g820(.A1(new_n727), .A2(G204gat), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n994), .A2(new_n936), .A3(new_n1022), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n1017), .A2(new_n727), .ZN(new_n1024));
  AOI22_X1  g823(.A1(new_n1023), .A2(KEYINPUT62), .B1(new_n1024), .B2(G204gat), .ZN(new_n1025));
  NOR3_X1   g824(.A1(new_n1023), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1026));
  INV_X1    g825(.A(KEYINPUT126), .ZN(new_n1027));
  OAI21_X1  g826(.A(KEYINPUT125), .B1(new_n899), .B2(new_n476), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n1028), .A2(new_n520), .A3(new_n936), .A4(new_n991), .ZN(new_n1029));
  INV_X1    g828(.A(new_n1022), .ZN(new_n1030));
  NOR2_X1   g829(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT62), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1027), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g832(.A(new_n1025), .B1(new_n1026), .B2(new_n1033), .ZN(G1353gat));
  NOR3_X1   g833(.A1(new_n1029), .A2(G211gat), .A3(new_n841), .ZN(new_n1035));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1036));
  OAI21_X1  g835(.A(KEYINPUT57), .B1(new_n899), .B2(new_n503), .ZN(new_n1037));
  NAND4_X1  g836(.A1(new_n1037), .A2(new_n690), .A3(new_n967), .A4(new_n1016), .ZN(new_n1038));
  AOI21_X1  g837(.A(KEYINPUT63), .B1(new_n1038), .B2(G211gat), .ZN(new_n1039));
  AOI21_X1  g838(.A(new_n1035), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1038), .A2(G211gat), .ZN(new_n1041));
  INV_X1    g840(.A(KEYINPUT63), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1038), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n1043), .A2(KEYINPUT127), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1040), .A2(new_n1045), .ZN(G1354gat));
  OAI21_X1  g845(.A(G218gat), .B1(new_n1017), .B2(new_n783), .ZN(new_n1047));
  OR2_X1    g846(.A1(new_n783), .A2(G218gat), .ZN(new_n1048));
  OAI21_X1  g847(.A(new_n1047), .B1(new_n1029), .B2(new_n1048), .ZN(G1355gat));
endmodule


