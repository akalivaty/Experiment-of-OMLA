

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n638), .A2(n523), .ZN(n641) );
  XOR2_X1 U549 ( .A(n753), .B(KEYINPUT100), .Z(n515) );
  XOR2_X2 U550 ( .A(KEYINPUT92), .B(n686), .Z(n765) );
  NOR2_X1 U551 ( .A1(n728), .A2(n727), .ZN(n729) );
  INV_X1 U552 ( .A(n979), .ZN(n756) );
  XNOR2_X1 U553 ( .A(n522), .B(n521), .ZN(n525) );
  XNOR2_X1 U554 ( .A(KEYINPUT78), .B(KEYINPUT4), .ZN(n521) );
  INV_X1 U555 ( .A(KEYINPUT80), .ZN(n531) );
  OR2_X1 U556 ( .A1(n712), .A2(n999), .ZN(n516) );
  BUF_X1 U557 ( .A(n688), .Z(n722) );
  OR2_X1 U558 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U559 ( .A1(n757), .A2(n756), .ZN(n758) );
  INV_X1 U560 ( .A(KEYINPUT75), .ZN(n584) );
  XNOR2_X1 U561 ( .A(n584), .B(KEYINPUT13), .ZN(n585) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n684) );
  XNOR2_X1 U563 ( .A(n586), .B(n585), .ZN(n587) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  NOR2_X1 U565 ( .A1(G651), .A2(G543), .ZN(n643) );
  NOR2_X2 U566 ( .A1(G2105), .A2(n537), .ZN(n879) );
  NOR2_X1 U567 ( .A1(G651), .A2(n638), .ZN(n651) );
  NOR2_X1 U568 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U569 ( .A(n531), .B(KEYINPUT8), .ZN(n532) );
  OR2_X1 U570 ( .A1(n548), .A2(n547), .ZN(n683) );
  XNOR2_X1 U571 ( .A(G168), .B(n532), .ZN(G286) );
  INV_X1 U572 ( .A(G651), .ZN(n523) );
  NOR2_X1 U573 ( .A1(G543), .A2(n523), .ZN(n517) );
  XOR2_X2 U574 ( .A(KEYINPUT1), .B(n517), .Z(n645) );
  NAND2_X1 U575 ( .A1(G63), .A2(n645), .ZN(n519) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  NAND2_X1 U577 ( .A1(G51), .A2(n651), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U579 ( .A(KEYINPUT6), .B(n520), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G89), .A2(n643), .ZN(n522) );
  NAND2_X1 U581 ( .A1(G76), .A2(n641), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U583 ( .A(n526), .B(KEYINPUT5), .Z(n527) );
  XOR2_X1 U584 ( .A(KEYINPUT79), .B(n529), .Z(n530) );
  XOR2_X1 U585 ( .A(KEYINPUT7), .B(n530), .Z(G168) );
  XOR2_X1 U586 ( .A(KEYINPUT17), .B(n533), .Z(n534) );
  XNOR2_X2 U587 ( .A(n534), .B(KEYINPUT64), .ZN(n880) );
  NAND2_X1 U588 ( .A1(n880), .A2(G138), .ZN(n541) );
  INV_X1 U589 ( .A(G2104), .ZN(n537) );
  AND2_X1 U590 ( .A1(n537), .A2(G2105), .ZN(n875) );
  NAND2_X1 U591 ( .A1(G126), .A2(n875), .ZN(n536) );
  AND2_X1 U592 ( .A1(G2105), .A2(G2104), .ZN(n876) );
  NAND2_X1 U593 ( .A1(G114), .A2(n876), .ZN(n535) );
  AND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G102), .A2(n879), .ZN(n538) );
  AND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U598 ( .A1(n875), .A2(G125), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G101), .A2(n879), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT23), .B(n542), .Z(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U602 ( .A1(G137), .A2(n880), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n876), .A2(G113), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U605 ( .A(n683), .ZN(G160) );
  NAND2_X1 U606 ( .A1(G64), .A2(n645), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G52), .A2(n651), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U609 ( .A(KEYINPUT66), .B(n551), .ZN(n558) );
  NAND2_X1 U610 ( .A1(n643), .A2(G90), .ZN(n552) );
  XNOR2_X1 U611 ( .A(KEYINPUT67), .B(n552), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n641), .A2(G77), .ZN(n553) );
  XOR2_X1 U613 ( .A(KEYINPUT68), .B(n553), .Z(n554) );
  NOR2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n556), .B(KEYINPUT9), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(G171) );
  NAND2_X1 U617 ( .A1(n880), .A2(G135), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n559), .B(KEYINPUT82), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G99), .A2(n879), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G111), .A2(n876), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n875), .A2(G123), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT18), .B(n562), .Z(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n918) );
  XNOR2_X1 U626 ( .A(G2096), .B(n918), .ZN(n567) );
  OR2_X1 U627 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  NAND2_X1 U631 ( .A1(G75), .A2(n641), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G88), .A2(n643), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G50), .A2(n651), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT86), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n645), .A2(G62), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n574), .A2(n573), .ZN(G166) );
  NAND2_X1 U639 ( .A1(G94), .A2(G452), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U643 ( .A(G223), .B(KEYINPUT72), .Z(n819) );
  NAND2_X1 U644 ( .A1(n819), .A2(G567), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT73), .ZN(n578) );
  XNOR2_X1 U646 ( .A(KEYINPUT11), .B(n578), .ZN(G234) );
  NAND2_X1 U647 ( .A1(n645), .A2(G56), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT14), .B(n579), .Z(n588) );
  NAND2_X1 U649 ( .A1(n643), .A2(G81), .ZN(n580) );
  XOR2_X1 U650 ( .A(KEYINPUT12), .B(n580), .Z(n583) );
  NAND2_X1 U651 ( .A1(n641), .A2(G68), .ZN(n581) );
  XOR2_X1 U652 ( .A(n581), .B(KEYINPUT74), .Z(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n586) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n651), .A2(G43), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n974) );
  INV_X1 U657 ( .A(G860), .ZN(n612) );
  OR2_X1 U658 ( .A1(n974), .A2(n612), .ZN(n591) );
  XNOR2_X1 U659 ( .A(KEYINPUT76), .B(n591), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U662 ( .A1(G54), .A2(n651), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G79), .A2(n641), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G92), .A2(n643), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G66), .A2(n645), .ZN(n594) );
  XNOR2_X1 U667 ( .A(KEYINPUT77), .B(n594), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X2 U670 ( .A(n599), .B(KEYINPUT15), .ZN(n970) );
  INV_X1 U671 ( .A(n970), .ZN(n702) );
  INV_X1 U672 ( .A(G868), .ZN(n662) );
  NAND2_X1 U673 ( .A1(n702), .A2(n662), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G65), .A2(n645), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT70), .ZN(n609) );
  NAND2_X1 U677 ( .A1(G78), .A2(n641), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G91), .A2(n643), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G53), .A2(n651), .ZN(n605) );
  XNOR2_X1 U681 ( .A(KEYINPUT71), .B(n605), .ZN(n606) );
  NOR2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(G299) );
  NAND2_X1 U684 ( .A1(G868), .A2(G286), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G299), .A2(n662), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n612), .A2(G559), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n613), .A2(n970), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n974), .ZN(n615) );
  XOR2_X1 U691 ( .A(KEYINPUT81), .B(n615), .Z(n618) );
  NAND2_X1 U692 ( .A1(G868), .A2(n970), .ZN(n616) );
  NOR2_X1 U693 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U695 ( .A1(n970), .A2(G559), .ZN(n660) );
  XNOR2_X1 U696 ( .A(n974), .B(n660), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n619), .A2(G860), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G67), .A2(n645), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G55), .A2(n651), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G80), .A2(n641), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G93), .A2(n643), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U704 ( .A(KEYINPUT83), .B(n624), .Z(n625) );
  OR2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n663) );
  XOR2_X1 U706 ( .A(n627), .B(n663), .Z(G145) );
  NAND2_X1 U707 ( .A1(G72), .A2(n641), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G85), .A2(n643), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U710 ( .A(KEYINPUT65), .B(n630), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G60), .A2(n645), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G47), .A2(n651), .ZN(n631) );
  AND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U715 ( .A1(G49), .A2(n651), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n645), .A2(n637), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G73), .A2(n641), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n642), .Z(n650) );
  NAND2_X1 U723 ( .A1(n643), .A2(G86), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT84), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G61), .A2(n645), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U727 ( .A(KEYINPUT85), .B(n648), .Z(n649) );
  NOR2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n651), .A2(G48), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(G305) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(G290), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(G288), .ZN(n657) );
  XNOR2_X1 U733 ( .A(G166), .B(G299), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n655), .B(n974), .ZN(n656) );
  XNOR2_X1 U735 ( .A(n657), .B(n656), .ZN(n659) );
  XOR2_X1 U736 ( .A(G305), .B(n663), .Z(n658) );
  XNOR2_X1 U737 ( .A(n659), .B(n658), .ZN(n893) );
  XOR2_X1 U738 ( .A(n893), .B(n660), .Z(n661) );
  NAND2_X1 U739 ( .A1(G868), .A2(n661), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n667), .ZN(n669) );
  XOR2_X1 U745 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n668) );
  XNOR2_X1 U746 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U747 ( .A1(G2072), .A2(n670), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U751 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U752 ( .A1(G96), .A2(n673), .ZN(n824) );
  NAND2_X1 U753 ( .A1(n824), .A2(G2106), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U755 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G108), .A2(n675), .ZN(n825) );
  NAND2_X1 U757 ( .A1(n825), .A2(G567), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n826) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n678) );
  XNOR2_X1 U760 ( .A(KEYINPUT88), .B(n678), .ZN(n679) );
  NOR2_X1 U761 ( .A1(n826), .A2(n679), .ZN(n821) );
  NAND2_X1 U762 ( .A1(n821), .A2(G36), .ZN(n680) );
  XOR2_X1 U763 ( .A(KEYINPUT89), .B(n680), .Z(G176) );
  INV_X1 U764 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U765 ( .A(G1986), .B(G290), .ZN(n969) );
  INV_X1 U766 ( .A(G40), .ZN(n682) );
  OR2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n684), .A2(n681), .ZN(n814) );
  NAND2_X1 U769 ( .A1(n969), .A2(n814), .ZN(n800) );
  NOR2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n688), .A2(G8), .ZN(n686) );
  INV_X1 U773 ( .A(n765), .ZN(n751) );
  XOR2_X1 U774 ( .A(KEYINPUT94), .B(KEYINPUT28), .Z(n692) );
  INV_X1 U775 ( .A(n688), .ZN(n712) );
  NAND2_X1 U776 ( .A1(n712), .A2(G2072), .ZN(n687) );
  XOR2_X1 U777 ( .A(KEYINPUT27), .B(n687), .Z(n690) );
  NAND2_X1 U778 ( .A1(G1956), .A2(n722), .ZN(n689) );
  NAND2_X1 U779 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U780 ( .A1(n693), .A2(G299), .ZN(n691) );
  XNOR2_X1 U781 ( .A(n692), .B(n691), .ZN(n710) );
  NOR2_X1 U782 ( .A1(G299), .A2(n693), .ZN(n694) );
  XOR2_X1 U783 ( .A(n694), .B(KEYINPUT97), .Z(n708) );
  XOR2_X1 U784 ( .A(G1996), .B(KEYINPUT95), .Z(n947) );
  NAND2_X1 U785 ( .A1(n712), .A2(n947), .ZN(n695) );
  XNOR2_X1 U786 ( .A(n695), .B(KEYINPUT26), .ZN(n696) );
  INV_X1 U787 ( .A(G1341), .ZN(n999) );
  NAND2_X1 U788 ( .A1(n696), .A2(n516), .ZN(n697) );
  NOR2_X1 U789 ( .A1(n974), .A2(n697), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n712), .A2(G1348), .ZN(n699) );
  NOR2_X1 U791 ( .A1(G2067), .A2(n722), .ZN(n698) );
  NOR2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n702), .A2(n703), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n705) );
  OR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U797 ( .A(n706), .B(KEYINPUT96), .ZN(n707) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U800 ( .A(n711), .B(KEYINPUT29), .ZN(n716) );
  XNOR2_X1 U801 ( .A(G1961), .B(KEYINPUT93), .ZN(n1008) );
  NAND2_X1 U802 ( .A1(n722), .A2(n1008), .ZN(n714) );
  XNOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .ZN(n941) );
  NAND2_X1 U804 ( .A1(n712), .A2(n941), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n726) );
  NAND2_X1 U806 ( .A1(G171), .A2(n726), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n738) );
  INV_X1 U808 ( .A(G8), .ZN(n721) );
  NOR2_X1 U809 ( .A1(n751), .A2(G1971), .ZN(n718) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n722), .ZN(n717) );
  NOR2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n719), .A2(G303), .ZN(n720) );
  OR2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n731) );
  AND2_X1 U814 ( .A1(n738), .A2(n731), .ZN(n730) );
  NOR2_X1 U815 ( .A1(n751), .A2(G1966), .ZN(n741) );
  NOR2_X1 U816 ( .A1(G2084), .A2(n722), .ZN(n737) );
  NOR2_X1 U817 ( .A1(n741), .A2(n737), .ZN(n723) );
  NAND2_X1 U818 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U819 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n725), .A2(G168), .ZN(n728) );
  NOR2_X1 U821 ( .A1(G171), .A2(n726), .ZN(n727) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n729), .Z(n739) );
  NAND2_X1 U823 ( .A1(n730), .A2(n739), .ZN(n735) );
  INV_X1 U824 ( .A(n731), .ZN(n733) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n732) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U827 ( .A(n736), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U828 ( .A1(G8), .A2(n737), .ZN(n743) );
  AND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X2 U833 ( .A(n746), .B(KEYINPUT98), .ZN(n761) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n754), .A2(n747), .ZN(n967) );
  NAND2_X1 U837 ( .A1(n761), .A2(n967), .ZN(n749) );
  NAND2_X1 U838 ( .A1(G288), .A2(G1976), .ZN(n748) );
  XOR2_X1 U839 ( .A(KEYINPUT99), .B(n748), .Z(n963) );
  NAND2_X1 U840 ( .A1(n749), .A2(n963), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U842 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  AND2_X1 U843 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n755), .A2(n765), .ZN(n757) );
  XNOR2_X1 U845 ( .A(G1981), .B(G305), .ZN(n979) );
  NAND2_X1 U846 ( .A1(n515), .A2(n758), .ZN(n770) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n759), .B(KEYINPUT24), .ZN(n760) );
  AND2_X1 U849 ( .A1(n760), .A2(n765), .ZN(n768) );
  INV_X1 U850 ( .A(n761), .ZN(n764) );
  NAND2_X1 U851 ( .A1(G166), .A2(G8), .ZN(n762) );
  NOR2_X1 U852 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n798) );
  XNOR2_X1 U857 ( .A(KEYINPUT37), .B(G2067), .ZN(n812) );
  NAND2_X1 U858 ( .A1(G104), .A2(n879), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G140), .A2(n880), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n773), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G128), .A2(n875), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G116), .A2(n876), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n779), .ZN(n890) );
  NOR2_X1 U868 ( .A1(n812), .A2(n890), .ZN(n921) );
  NAND2_X1 U869 ( .A1(n814), .A2(n921), .ZN(n810) );
  XNOR2_X1 U870 ( .A(KEYINPUT90), .B(n814), .ZN(n795) );
  NAND2_X1 U871 ( .A1(G95), .A2(n879), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G119), .A2(n875), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n876), .A2(G107), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G131), .A2(n880), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n784) );
  OR2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n861) );
  NAND2_X1 U878 ( .A1(G1991), .A2(n861), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G129), .A2(n875), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G117), .A2(n876), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n879), .A2(G105), .ZN(n788) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U885 ( .A1(G141), .A2(n880), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n855) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n855), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n915) );
  NAND2_X1 U889 ( .A1(n795), .A2(n915), .ZN(n804) );
  XOR2_X1 U890 ( .A(KEYINPUT91), .B(n804), .Z(n796) );
  AND2_X1 U891 ( .A1(n810), .A2(n796), .ZN(n797) );
  AND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n817) );
  NOR2_X1 U894 ( .A1(G1991), .A2(n861), .ZN(n801) );
  XNOR2_X1 U895 ( .A(KEYINPUT103), .B(n801), .ZN(n922) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n802) );
  XOR2_X1 U897 ( .A(n802), .B(KEYINPUT102), .Z(n803) );
  NAND2_X1 U898 ( .A1(n922), .A2(n803), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n855), .A2(G1996), .ZN(n806) );
  XNOR2_X1 U901 ( .A(n806), .B(KEYINPUT101), .ZN(n912) );
  NAND2_X1 U902 ( .A1(n807), .A2(n912), .ZN(n809) );
  XOR2_X1 U903 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n808) );
  XNOR2_X1 U904 ( .A(n809), .B(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n812), .A2(n890), .ZN(n916) );
  NAND2_X1 U907 ( .A1(n813), .A2(n916), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n818), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U913 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U916 ( .A(KEYINPUT105), .B(n823), .Z(G188) );
  INV_X1 U918 ( .A(G120), .ZN(G236) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  INV_X1 U923 ( .A(n826), .ZN(G319) );
  XOR2_X1 U924 ( .A(KEYINPUT41), .B(G1961), .Z(n828) );
  XNOR2_X1 U925 ( .A(G1996), .B(G1991), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U927 ( .A(n829), .B(KEYINPUT109), .Z(n831) );
  XNOR2_X1 U928 ( .A(G1981), .B(G1966), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U930 ( .A(G1976), .B(G1971), .Z(n833) );
  XNOR2_X1 U931 ( .A(G1986), .B(G1956), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U933 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U934 ( .A(KEYINPUT108), .B(G2474), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(G229) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(G2678), .Z(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2072), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2090), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2096), .B(G2100), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U945 ( .A(G2078), .B(G2084), .Z(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(G227) );
  NAND2_X1 U947 ( .A1(G124), .A2(n875), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n879), .A2(G100), .ZN(n849) );
  NAND2_X1 U950 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U951 ( .A1(n876), .A2(G112), .ZN(n852) );
  NAND2_X1 U952 ( .A1(G136), .A2(n880), .ZN(n851) );
  NAND2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U954 ( .A1(n854), .A2(n853), .ZN(G162) );
  XNOR2_X1 U955 ( .A(n855), .B(G162), .ZN(n857) );
  XNOR2_X1 U956 ( .A(G164), .B(G160), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n865) );
  XNOR2_X1 U958 ( .A(KEYINPUT111), .B(KEYINPUT114), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n918), .B(KEYINPUT46), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT110), .B(n860), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n861), .B(KEYINPUT48), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U964 ( .A(n865), .B(n864), .Z(n888) );
  NAND2_X1 U965 ( .A1(G103), .A2(n879), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G139), .A2(n880), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U968 ( .A1(n876), .A2(G115), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n868), .B(KEYINPUT112), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G127), .A2(n875), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(n871), .ZN(n872) );
  XNOR2_X1 U973 ( .A(KEYINPUT113), .B(n872), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n929) );
  NAND2_X1 U975 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U978 ( .A1(G106), .A2(n879), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G142), .A2(n880), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n929), .B(n886), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n890), .B(n889), .Z(n891) );
  NOR2_X1 U986 ( .A1(G37), .A2(n891), .ZN(n892) );
  XOR2_X1 U987 ( .A(KEYINPUT115), .B(n892), .Z(G395) );
  XNOR2_X1 U988 ( .A(G286), .B(n893), .ZN(n895) );
  XNOR2_X1 U989 ( .A(G171), .B(n970), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U991 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U992 ( .A(G2451), .B(G2430), .Z(n898) );
  XNOR2_X1 U993 ( .A(G2438), .B(G2443), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n904) );
  XOR2_X1 U995 ( .A(G2435), .B(G2454), .Z(n900) );
  XNOR2_X1 U996 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U998 ( .A(G2446), .B(G2427), .Z(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1011 ( .A(G2090), .B(G162), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(KEYINPUT51), .ZN(n928) );
  INV_X1 U1014 ( .A(n915), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n926) );
  XNOR2_X1 U1016 ( .A(G160), .B(G2084), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n934) );
  XOR2_X1 U1023 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1026 ( .A(KEYINPUT50), .B(n932), .Z(n933) );
  NOR2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n935), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n957) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n957), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n937), .A2(G29), .ZN(n1019) );
  XOR2_X1 U1032 ( .A(G29), .B(KEYINPUT120), .Z(n960) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(G1991), .B(G25), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n946) );
  XOR2_X1 U1036 ( .A(G2072), .B(G33), .Z(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(G28), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G27), .B(n941), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G32), .B(n947), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1044 ( .A(KEYINPUT53), .B(n950), .Z(n953) );
  XOR2_X1 U1045 ( .A(KEYINPUT54), .B(G34), .Z(n951) );
  XNOR2_X1 U1046 ( .A(G2084), .B(n951), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(KEYINPUT118), .B(G2090), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G35), .B(n954), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n958) );
  XOR2_X1 U1051 ( .A(n958), .B(n957), .Z(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n961), .ZN(n1017) );
  XNOR2_X1 U1054 ( .A(G16), .B(KEYINPUT56), .ZN(n987) );
  NAND2_X1 U1055 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G1956), .B(G299), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n985) );
  XOR2_X1 U1061 ( .A(G1348), .B(n970), .Z(n972) );
  XOR2_X1 U1062 ( .A(G171), .B(G1961), .Z(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT122), .B(n973), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(G1341), .B(KEYINPUT123), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n983) );
  XOR2_X1 U1068 ( .A(G168), .B(G1966), .Z(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT57), .B(n980), .Z(n981) );
  XNOR2_X1 U1071 ( .A(n981), .B(KEYINPUT121), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n1015) );
  INV_X1 U1075 ( .A(G16), .ZN(n1013) );
  XOR2_X1 U1076 ( .A(G1986), .B(G24), .Z(n991) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n993), .B(n992), .ZN(n1007) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(G4), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G20), .B(G1956), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(KEYINPUT124), .B(n999), .Z(n1000) );
  XNOR2_X1 U1090 ( .A(G19), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1096 ( .A(G5), .B(n1008), .Z(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(n1020), .B(KEYINPUT126), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1021), .ZN(G150) );
  INV_X1 U1105 ( .A(G150), .ZN(G311) );
endmodule

