//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT88), .ZN(new_n211));
  NAND2_X1  g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT88), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n204), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n218), .A2(new_n203), .A3(new_n210), .A4(new_n212), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT89), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n215), .A2(new_n219), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT90), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n220), .B2(new_n221), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT96), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(G85gat), .A3(G92gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233));
  INV_X1    g032(.A(G85gat), .ZN(new_n234));
  INV_X1    g033(.A(G92gat), .ZN(new_n235));
  AOI22_X1  g034(.A1(KEYINPUT8), .A2(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n229), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G99gat), .B(G106gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n228), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n238), .B(new_n239), .ZN(new_n242));
  AND2_X1   g041(.A1(G232gat), .A2(G233gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n220), .A2(new_n242), .B1(KEYINPUT41), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(G190gat), .B(G218gat), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n243), .A2(KEYINPUT41), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(G162gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n245), .A2(new_n246), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT98), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n247), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(KEYINPUT97), .ZN(new_n255));
  INV_X1    g054(.A(new_n251), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n245), .B(new_n246), .C1(KEYINPUT98), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n255), .B1(new_n254), .B2(new_n257), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G22gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT16), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(G1gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(G1gat), .B2(new_n262), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(G8gat), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267));
  NOR2_X1   g066(.A1(G71gat), .A2(G78gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n268), .B(KEYINPUT93), .Z(new_n269));
  INV_X1    g068(.A(G57gat), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n270), .A2(G64gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(G64gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT9), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G71gat), .ZN(new_n274));
  INV_X1    g073(.A(G78gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n269), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n278));
  OR3_X1    g077(.A1(new_n270), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT94), .B1(new_n270), .B2(G64gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n281), .B2(new_n271), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G211gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G127gat), .B(G155gat), .Z(new_n287));
  OR2_X1    g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n287), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n267), .ZN(new_n290));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n288), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n288), .B2(new_n289), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT95), .B(G183gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OR3_X1    g098(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n294), .B2(new_n295), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n242), .A2(new_n282), .A3(new_n276), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT10), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n240), .A2(new_n283), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n304), .A3(new_n303), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n305), .A2(new_n307), .B1(G230gat), .B2(G233gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G230gat), .A2(G233gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n306), .B2(new_n303), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT99), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G120gat), .B(G148gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT100), .ZN(new_n313));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  OR2_X1    g114(.A1(new_n310), .A2(KEYINPUT99), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n311), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n315), .B1(new_n311), .B2(new_n316), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n261), .A2(new_n302), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT101), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT101), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n261), .A2(new_n302), .A3(new_n323), .A4(new_n320), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n265), .B(G8gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n225), .B2(new_n227), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n223), .A2(new_n327), .B1(new_n326), .B2(new_n220), .ZN(new_n328));
  NAND2_X1  g127(.A1(G229gat), .A2(G233gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n329), .B(KEYINPUT91), .Z(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(KEYINPUT18), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n266), .A2(new_n224), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n220), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n330), .B(KEYINPUT13), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT18), .B1(new_n328), .B2(new_n330), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G113gat), .B(G141gat), .ZN(new_n341));
  INV_X1    g140(.A(G197gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT11), .B(G169gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(KEYINPUT12), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n338), .B(new_n340), .C1(KEYINPUT92), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n331), .A2(KEYINPUT92), .A3(new_n336), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n349), .B(new_n346), .C1(new_n337), .C2(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n353), .B(KEYINPUT81), .Z(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356));
  INV_X1    g155(.A(G204gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G197gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(G211gat), .A2(G218gat), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n362), .A2(KEYINPUT22), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(G197gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(G204gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n368));
  NOR2_X1   g167(.A1(G211gat), .A2(G218gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G218gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n285), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G211gat), .A2(G218gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(KEYINPUT73), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT72), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n367), .B(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G141gat), .B(G148gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(G155gat), .B2(G162gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n380), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G141gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G148gat), .ZN(new_n386));
  INV_X1    g185(.A(G148gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G141gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G155gat), .B(G162gat), .ZN(new_n390));
  INV_X1    g189(.A(G155gat), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT2), .B1(new_n391), .B2(new_n250), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n356), .B1(new_n377), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n376), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n367), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n376), .A2(new_n363), .A3(new_n366), .A4(new_n361), .ZN(new_n401));
  AND4_X1   g200(.A1(new_n356), .A2(new_n397), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n370), .A2(new_n374), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n367), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n396), .B1(new_n367), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n394), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n384), .A2(new_n393), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n355), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(G228gat), .A3(G233gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n394), .B1(new_n377), .B2(KEYINPUT29), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n410), .A2(G22gat), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT31), .B(G50gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT83), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n377), .A2(new_n356), .A3(new_n397), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n409), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n413), .A2(new_n408), .ZN(new_n424));
  INV_X1    g223(.A(new_n412), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n423), .A2(new_n354), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G22gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(G22gat), .B(new_n419), .C1(new_n410), .C2(new_n414), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n415), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n427), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n420), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G127gat), .ZN(new_n434));
  INV_X1    g233(.A(G134gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G127gat), .A2(G134gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT1), .ZN(new_n439));
  INV_X1    g238(.A(G120gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G113gat), .ZN(new_n441));
  INV_X1    g240(.A(G113gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G120gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n438), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G113gat), .B(G120gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n438), .B1(new_n447), .B2(KEYINPUT68), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(new_n443), .A3(KEYINPUT68), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n439), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT69), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n444), .A2(new_n453), .B1(new_n436), .B2(new_n437), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT1), .B1(new_n447), .B2(KEYINPUT68), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT69), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n446), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n384), .A2(new_n393), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT75), .B1(new_n458), .B2(new_n394), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT75), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n408), .A2(new_n460), .A3(KEYINPUT3), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n457), .A2(new_n395), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n451), .B1(new_n448), .B2(new_n450), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n454), .A2(KEYINPUT69), .A3(new_n455), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND4_X1   g265(.A1(new_n463), .A2(new_n466), .A3(new_n446), .A4(new_n458), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n445), .B1(new_n464), .B2(new_n465), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n463), .B1(new_n468), .B2(new_n458), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n462), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n408), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n466), .A2(new_n446), .A3(new_n458), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(KEYINPUT76), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT76), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n477), .A3(new_n408), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n473), .B(KEYINPUT39), .C1(new_n479), .C2(new_n472), .ZN(new_n480));
  XNOR2_X1  g279(.A(G57gat), .B(G85gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT79), .ZN(new_n482));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT78), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n482), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n475), .A2(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n463), .A3(new_n458), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n471), .B1(new_n491), .B2(new_n462), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT39), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n480), .A2(new_n494), .A3(KEYINPUT40), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n462), .B(new_n471), .C1(new_n467), .C2(new_n469), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n491), .A2(KEYINPUT5), .A3(new_n471), .A4(new_n462), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n472), .A3(new_n478), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n488), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(KEYINPUT29), .ZN(new_n504));
  AND2_X1   g303(.A1(G169gat), .A2(G176gat), .ZN(new_n505));
  INV_X1    g304(.A(G169gat), .ZN(new_n506));
  INV_X1    g305(.A(G176gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT23), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G183gat), .A2(G190gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(G183gat), .A2(G190gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT23), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n510), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n510), .A2(new_n516), .A3(new_n519), .A4(new_n517), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G183gat), .ZN(new_n527));
  INV_X1    g326(.A(G190gat), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT28), .B(new_n528), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT66), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n505), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n541));
  NOR2_X1   g340(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n508), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n511), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n534), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n504), .B1(new_n526), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n524), .B1(new_n521), .B2(new_n522), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n534), .A2(new_n544), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n547), .A2(new_n548), .A3(new_n503), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n377), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n526), .A2(new_n545), .A3(new_n502), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n547), .A2(new_n548), .B1(KEYINPUT29), .B2(new_n503), .ZN(new_n552));
  INV_X1    g351(.A(new_n377), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G8gat), .B(G36gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT74), .ZN(new_n557));
  XNOR2_X1  g356(.A(G64gat), .B(G92gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OR3_X1    g359(.A1(new_n555), .A2(KEYINPUT30), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n560), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n550), .A2(new_n554), .A3(new_n559), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT30), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n495), .A2(new_n501), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n480), .A2(new_n494), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT40), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n433), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n559), .B1(new_n555), .B2(KEYINPUT37), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n571), .A3(new_n554), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT86), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT38), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT86), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n550), .A2(new_n554), .A3(new_n575), .A4(new_n571), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n570), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n570), .A2(new_n573), .A3(new_n576), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT87), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT38), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n578), .B2(KEYINPUT38), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n563), .B(new_n577), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n498), .A2(new_n500), .A3(new_n499), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n487), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n586), .A3(new_n501), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT85), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n501), .A2(new_n586), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT6), .B1(new_n584), .B2(new_n487), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(KEYINPUT85), .A3(new_n501), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n569), .B1(new_n583), .B2(new_n594), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n430), .A2(KEYINPUT84), .A3(new_n432), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n420), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n423), .A2(new_n354), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n424), .A2(new_n425), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n601), .B2(G22gat), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n426), .A2(new_n427), .A3(new_n418), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n431), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n432), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n597), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT80), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n501), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n501), .A2(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n611), .A3(new_n592), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n591), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n564), .A2(new_n561), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n526), .A2(new_n545), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n457), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G227gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT64), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n547), .A2(new_n548), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n618), .A3(new_n457), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n627), .A2(KEYINPUT32), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT34), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n621), .A2(new_n626), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(new_n622), .ZN(new_n631));
  AOI211_X1 g430(.A(KEYINPUT34), .B(new_n624), .C1(new_n621), .C2(new_n626), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G15gat), .B(G43gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G71gat), .B(G99gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  AND2_X1   g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n627), .A2(KEYINPUT32), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n630), .A2(new_n629), .A3(new_n623), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n621), .A2(new_n626), .B1(G227gat), .B2(G233gat), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n640), .B(new_n641), .C1(new_n629), .C2(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n633), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n639), .B1(new_n633), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT36), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n595), .A2(new_n616), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n594), .A2(new_n606), .A3(new_n646), .A4(new_n614), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT35), .ZN(new_n653));
  NOR4_X1   g452(.A1(new_n433), .A2(new_n644), .A3(new_n645), .A4(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n614), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n612), .B2(new_n591), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n652), .A2(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n352), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n325), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n613), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n655), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(G8gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n659), .A2(new_n671), .A3(new_n650), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n660), .A2(new_n646), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(G1326gat));
  INV_X1    g473(.A(KEYINPUT84), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n604), .B2(new_n605), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n596), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n659), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n592), .A2(KEYINPUT85), .A3(new_n501), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT85), .B1(new_n592), .B2(new_n501), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n682), .A2(new_n683), .A3(new_n590), .ZN(new_n684));
  INV_X1    g483(.A(new_n639), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT70), .B1(new_n466), .B2(new_n446), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n618), .B(new_n445), .C1(new_n464), .C2(new_n465), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n625), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NOR4_X1   g488(.A1(new_n468), .A2(new_n547), .A3(new_n548), .A4(KEYINPUT70), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n622), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT34), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n640), .B1(new_n692), .B2(new_n641), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n685), .B1(new_n686), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n633), .A2(new_n643), .A3(new_n639), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n606), .A2(new_n694), .A3(new_n614), .A4(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n653), .B1(new_n684), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n654), .A2(new_n656), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT36), .B1(new_n694), .B2(new_n695), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n677), .A2(new_n656), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n567), .A2(KEYINPUT40), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n606), .B1(new_n565), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n577), .A2(new_n563), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n578), .A2(KEYINPUT38), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT87), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(new_n580), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n684), .B2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n697), .B(new_n698), .C1(new_n701), .C2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n260), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n258), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n261), .B1(new_n651), .B2(new_n657), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n320), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n302), .A2(new_n718), .A3(new_n352), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n681), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AOI211_X1 g519(.A(KEYINPUT44), .B(new_n261), .C1(new_n651), .C2(new_n657), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n715), .B1(new_n709), .B2(new_n711), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n681), .B(new_n719), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n613), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n714), .A2(new_n719), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(G29gat), .A3(new_n613), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(G1328gat));
  OAI21_X1  g530(.A(G36gat), .B1(new_n725), .B2(new_n614), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n727), .A2(G36gat), .A3(new_n614), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1329gat));
  INV_X1    g534(.A(new_n650), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n720), .B2(new_n724), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(KEYINPUT104), .A3(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n650), .B1(new_n741), .B2(new_n723), .ZN(new_n742));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n646), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n727), .A2(G43gat), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT105), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n738), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G43gat), .B1(new_n740), .B2(new_n650), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(KEYINPUT47), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1330gat));
  OAI21_X1  g552(.A(G50gat), .B1(new_n740), .B2(new_n606), .ZN(new_n754));
  INV_X1    g553(.A(new_n727), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n677), .A2(new_n756), .A3(G50gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n677), .B2(G50gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n754), .A2(KEYINPUT48), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n759), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n608), .B1(new_n720), .B2(new_n724), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n760), .B1(new_n763), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n351), .A2(new_n320), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n709), .A2(new_n302), .A3(new_n261), .A4(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n613), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(new_n270), .ZN(G1332gat));
  INV_X1    g571(.A(new_n770), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT49), .B(G64gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(new_n655), .A3(new_n774), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n770), .A2(new_n614), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT108), .ZN(G1333gat));
  OAI21_X1  g577(.A(new_n274), .B1(new_n770), .B2(new_n745), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n736), .A2(G71gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g581(.A1(new_n770), .A2(new_n677), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(new_n275), .ZN(G1335gat));
  INV_X1    g583(.A(new_n302), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n717), .A2(new_n785), .A3(new_n765), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G85gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n712), .A2(new_n302), .A3(new_n351), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT51), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n661), .A3(new_n718), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n789), .A2(new_n661), .B1(new_n792), .B2(new_n234), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n718), .A2(new_n235), .A3(new_n655), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT109), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n235), .B1(new_n787), .B2(new_n655), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n787), .B2(new_n655), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n786), .A2(KEYINPUT110), .A3(new_n614), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n801), .A2(new_n235), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n799), .B2(new_n803), .ZN(G1337gat));
  NAND2_X1  g603(.A1(new_n787), .A2(G99gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n718), .A3(new_n646), .ZN(new_n807));
  INV_X1    g606(.A(G99gat), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n806), .A2(new_n736), .B1(new_n807), .B2(new_n808), .ZN(G1338gat));
  INV_X1    g608(.A(G106gat), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n810), .A3(new_n718), .A4(new_n433), .ZN(new_n811));
  OR2_X1    g610(.A1(KEYINPUT111), .A2(KEYINPUT53), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT53), .B(G106gat), .C1(new_n786), .C2(new_n677), .ZN(new_n814));
  OAI21_X1  g613(.A(G106gat), .B1(new_n786), .B2(new_n606), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n811), .B2(KEYINPUT111), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n813), .A2(new_n814), .B1(new_n816), .B2(new_n817), .ZN(G1339gat));
  NOR2_X1   g617(.A1(new_n321), .A2(new_n351), .ZN(new_n819));
  AND4_X1   g618(.A1(G230gat), .A2(new_n305), .A3(G233gat), .A4(new_n307), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n308), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  INV_X1    g621(.A(new_n315), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n308), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n823), .A4(new_n825), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n317), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n826), .A2(KEYINPUT113), .A3(new_n827), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n352), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n340), .A2(new_n336), .A3(new_n331), .A4(new_n347), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT114), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n328), .A2(new_n330), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n345), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n718), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT115), .B1(new_n841), .B2(new_n320), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n261), .B1(new_n835), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n834), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n711), .A3(new_n842), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n819), .B1(new_n850), .B2(new_n785), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(new_n608), .A3(new_n745), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n613), .A2(new_n655), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n352), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n851), .A2(new_n613), .A3(new_n696), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n351), .A2(new_n442), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT116), .Z(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n856), .A2(new_n440), .A3(new_n718), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  INV_X1    g663(.A(new_n854), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n718), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n866), .B2(G120gat), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT118), .B(new_n440), .C1(new_n865), .C2(new_n718), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n856), .B2(new_n302), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n785), .A2(new_n434), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n865), .B2(new_n871), .ZN(G1342gat));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n435), .A3(new_n711), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT56), .Z(new_n874));
  OAI21_X1  g673(.A(G134gat), .B1(new_n854), .B2(new_n261), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1343gat));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n851), .B2(new_n606), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n351), .A2(new_n832), .A3(new_n828), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n842), .A2(new_n718), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n261), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n849), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n785), .ZN(new_n884));
  INV_X1    g683(.A(new_n819), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT57), .A4(new_n608), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n302), .B1(new_n882), .B2(new_n849), .ZN(new_n889));
  OAI211_X1 g688(.A(KEYINPUT57), .B(new_n608), .C1(new_n889), .C2(new_n819), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT119), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n878), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n650), .A2(new_n853), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n351), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n851), .A2(new_n606), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n896), .A2(new_n893), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n385), .A3(new_n351), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  NAND3_X1  g702(.A1(new_n322), .A2(new_n324), .A3(new_n352), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT57), .B(new_n677), .C1(new_n884), .C2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n896), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n893), .B(KEYINPUT120), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n718), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n897), .A2(new_n387), .A3(new_n718), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n893), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n387), .B1(new_n913), .B2(new_n718), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n910), .B(new_n911), .C1(new_n914), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g714(.A(G155gat), .B1(new_n897), .B2(new_n302), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n912), .A2(new_n785), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G155gat), .ZN(G1346gat));
  NAND3_X1  g717(.A1(new_n897), .A2(new_n250), .A3(new_n711), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT121), .ZN(new_n920));
  OAI21_X1  g719(.A(G162gat), .B1(new_n912), .B2(new_n261), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n851), .A2(new_n661), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n745), .A2(new_n433), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n655), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n506), .A3(new_n351), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n661), .A2(new_n614), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n852), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n352), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n930), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n926), .B2(new_n718), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n929), .A2(new_n507), .A3(new_n320), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n926), .A2(new_n302), .A3(new_n527), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n929), .B2(new_n785), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n929), .B2(new_n261), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT123), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n942), .B(G190gat), .C1(new_n929), .C2(new_n261), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(KEYINPUT61), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n528), .A3(new_n711), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(KEYINPUT123), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(G1351gat));
  NAND3_X1  g747(.A1(new_n650), .A2(new_n433), .A3(new_n655), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT124), .Z(new_n950));
  NAND4_X1  g749(.A1(new_n923), .A2(new_n342), .A3(new_n351), .A4(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n896), .A2(new_n877), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n928), .A2(new_n650), .ZN(new_n953));
  NOR4_X1   g752(.A1(new_n952), .A2(new_n352), .A3(new_n905), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n954), .B2(new_n342), .ZN(G1352gat));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n923), .A2(new_n357), .A3(new_n950), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n957), .A2(new_n320), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n958), .B2(KEYINPUT62), .ZN(new_n959));
  OR4_X1    g758(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT62), .A4(new_n320), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(KEYINPUT62), .B1(new_n957), .B2(new_n320), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n953), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n907), .A2(new_n718), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n961), .A2(new_n964), .A3(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n907), .A2(new_n302), .A3(new_n965), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n923), .A2(new_n950), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n302), .A2(new_n285), .ZN(new_n973));
  OAI22_X1  g772(.A1(new_n970), .A2(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  NAND4_X1  g773(.A1(new_n923), .A2(new_n371), .A3(new_n711), .A4(new_n950), .ZN(new_n975));
  NOR4_X1   g774(.A1(new_n952), .A2(new_n261), .A3(new_n905), .A4(new_n953), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n371), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n979), .B(new_n975), .C1(new_n976), .C2(new_n371), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1355gat));
endmodule


