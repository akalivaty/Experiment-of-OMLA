//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  XNOR2_X1  g000(.A(KEYINPUT73), .B(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT69), .B(G953), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G210), .A3(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT2), .B(G113), .Z(new_n196));
  XNOR2_X1  g010(.A(G116), .B(G119), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G137), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n202), .A2(new_n204), .A3(new_n208), .A4(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n213), .A2(KEYINPUT0), .A3(G128), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n211), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(KEYINPUT0), .B2(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n211), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n210), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n220), .B2(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n220), .A2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n218), .A2(G143), .ZN(new_n228));
  OAI211_X1 g042(.A(G128), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n201), .A2(G137), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n203), .A2(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G128), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n219), .B(new_n221), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n209), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n199), .A2(new_n225), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT71), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(KEYINPUT71), .A3(new_n237), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n195), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n229), .A2(new_n234), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n209), .A2(new_n232), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT68), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n225), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n198), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n244), .A2(new_n199), .A3(new_n225), .A4(new_n246), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n247), .A2(KEYINPUT72), .A3(new_n198), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(KEYINPUT28), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n188), .B1(new_n241), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n240), .A2(new_n238), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT66), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n235), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT0), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n233), .A3(KEYINPUT64), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n222), .A2(new_n262), .B1(KEYINPUT0), .B2(G128), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n211), .A2(new_n216), .B1(new_n219), .B2(new_n221), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT65), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n215), .A2(new_n223), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n210), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n199), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n250), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n256), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n255), .A2(new_n271), .A3(new_n194), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n244), .A2(new_n225), .A3(new_n246), .A4(KEYINPUT30), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n198), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n260), .C2(new_n268), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT66), .B1(new_n242), .B2(new_n243), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n235), .A2(new_n258), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n268), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n277), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n194), .B1(new_n285), .B2(new_n250), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n254), .B1(new_n274), .B2(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n224), .A2(KEYINPUT65), .B1(new_n209), .B2(new_n207), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n267), .A2(new_n288), .B1(new_n257), .B2(new_n259), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT67), .B1(new_n289), .B2(KEYINPUT30), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n282), .A2(new_n279), .A3(new_n283), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n276), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n194), .A2(new_n250), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT31), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n255), .A2(new_n271), .ZN(new_n295));
  INV_X1    g109(.A(new_n194), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  INV_X1    g112(.A(new_n293), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n285), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n287), .A2(G472), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n302), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT81), .ZN(new_n311));
  INV_X1    g125(.A(G107), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G104), .ZN(new_n313));
  INV_X1    g127(.A(G104), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT81), .A3(G107), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n312), .A2(KEYINPUT3), .A3(G104), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT3), .B1(new_n312), .B2(G104), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n313), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G101), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n314), .B2(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n312), .A2(KEYINPUT3), .A3(G104), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT82), .B(G101), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n313), .A4(new_n315), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(KEYINPUT4), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT83), .ZN(new_n327));
  INV_X1    g141(.A(G101), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n313), .A2(new_n315), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(new_n323), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND4_X1   g146(.A1(new_n327), .A2(new_n318), .A3(new_n331), .A4(G101), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n198), .B(new_n326), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n314), .A2(G107), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n312), .A2(G104), .ZN(new_n336));
  OAI21_X1  g150(.A(G101), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n325), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n197), .A2(KEYINPUT5), .ZN(new_n339));
  INV_X1    g153(.A(G116), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n340), .A2(KEYINPUT5), .A3(G119), .ZN(new_n341));
  INV_X1    g155(.A(G113), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n339), .A2(new_n343), .B1(new_n196), .B2(new_n197), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n334), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n334), .A2(new_n345), .A3(new_n347), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n229), .A2(new_n234), .ZN(new_n353));
  INV_X1    g167(.A(G125), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n215), .A2(new_n223), .A3(G125), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n352), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT87), .B(G224), .ZN(new_n361));
  INV_X1    g175(.A(G953), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n360), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n346), .A2(new_n365), .A3(new_n348), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n351), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n355), .A2(new_n356), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT86), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(KEYINPUT7), .A3(new_n363), .A4(new_n358), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n347), .B(KEYINPUT8), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n338), .A2(new_n344), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n338), .A2(new_n344), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT88), .B(KEYINPUT7), .Z(new_n375));
  NAND2_X1  g189(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n357), .B2(new_n359), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n370), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n378), .B2(new_n350), .ZN(new_n379));
  OAI21_X1  g193(.A(G210), .B1(G237), .B2(G902), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n367), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n367), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n310), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n354), .A2(G140), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n354), .A2(KEYINPUT77), .A3(G140), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT16), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n391), .A2(new_n218), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n218), .B1(new_n391), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n384), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G146), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n218), .A3(new_n393), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(KEYINPUT89), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n362), .A2(KEYINPUT69), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT69), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n401), .A2(new_n403), .A3(G214), .A4(new_n190), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n220), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n189), .A2(G143), .A3(G214), .A4(new_n190), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G131), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n406), .A3(new_n208), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(KEYINPUT17), .A3(G131), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n396), .A2(new_n400), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(KEYINPUT18), .A2(G131), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n414), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n386), .A2(new_n387), .A3(new_n218), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n389), .A2(new_n390), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n218), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n314), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n413), .A2(new_n424), .A3(new_n421), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G902), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT90), .B(G475), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G122), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT14), .B1(new_n437), .B2(G116), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n340), .B2(G122), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT92), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n340), .A2(G122), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT92), .B1(new_n442), .B2(KEYINPUT14), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n441), .B(G107), .C1(new_n439), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(G116), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n445), .A2(new_n442), .A3(new_n312), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n220), .A2(G128), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n220), .A2(G128), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n448), .A2(new_n449), .A3(G134), .ZN(new_n450));
  OAI21_X1  g264(.A(G134), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n446), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n312), .B1(new_n445), .B2(new_n442), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n449), .B1(new_n457), .B2(new_n447), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n448), .A2(KEYINPUT13), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n201), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n454), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n446), .A2(new_n455), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(KEYINPUT91), .A3(new_n463), .A4(new_n450), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n453), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  INV_X1    g280(.A(G217), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n466), .A2(new_n467), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n453), .A2(new_n461), .A3(new_n464), .A4(new_n468), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n436), .B1(new_n472), .B2(new_n187), .ZN(new_n473));
  AOI211_X1 g287(.A(new_n188), .B(new_n435), .C1(new_n470), .C2(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n362), .A2(G952), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(G234), .B2(G237), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n189), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(G898), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n473), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(G475), .A2(G902), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n408), .A2(new_n410), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT19), .B1(new_n386), .B2(new_n387), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n419), .B2(KEYINPUT19), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n398), .B1(new_n485), .B2(G146), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n421), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n425), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n482), .B1(new_n488), .B2(new_n427), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT20), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI211_X1 g305(.A(KEYINPUT20), .B(new_n482), .C1(new_n488), .C2(new_n427), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n433), .B(new_n480), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n383), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT74), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n233), .B2(G119), .ZN(new_n497));
  INV_X1    g311(.A(G119), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT74), .A3(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n233), .A2(G119), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G110), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT24), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT24), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G110), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT75), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT75), .B1(new_n503), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n498), .B2(G128), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n233), .A2(KEYINPUT23), .A3(G119), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n498), .A2(G128), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n502), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n417), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n398), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n394), .A2(new_n395), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n506), .A2(new_n507), .ZN(new_n517));
  INV_X1    g331(.A(new_n501), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(new_n512), .A3(new_n511), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(G110), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n520), .B2(G110), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n515), .B1(new_n516), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT22), .B(G137), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n520), .A2(G110), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n522), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n534), .B(new_n519), .C1(new_n394), .C2(new_n395), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n515), .A3(new_n529), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n467), .B1(new_n187), .B2(G234), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G902), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT79), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n531), .A2(KEYINPUT79), .A3(new_n536), .A4(new_n538), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n537), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n531), .A2(new_n187), .A3(new_n536), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT78), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT25), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n495), .B(new_n543), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n535), .A2(new_n515), .A3(new_n529), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n529), .B1(new_n535), .B2(new_n515), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(new_n188), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n548), .B1(new_n554), .B2(KEYINPUT78), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n550), .A3(new_n537), .ZN(new_n556));
  INV_X1    g370(.A(new_n543), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT80), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G221), .B1(new_n466), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n224), .B(new_n326), .C1(new_n332), .C2(new_n333), .ZN(new_n562));
  INV_X1    g376(.A(new_n210), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n242), .A2(new_n325), .A3(new_n337), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT10), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n325), .A2(new_n337), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n353), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT10), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n562), .A2(new_n563), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n325), .A2(new_n337), .B1(new_n234), .B2(new_n229), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT84), .B(new_n210), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT85), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT12), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n567), .A2(new_n353), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n563), .B1(new_n564), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT85), .B1(new_n576), .B2(KEYINPUT84), .ZN(new_n577));
  OAI211_X1 g391(.A(KEYINPUT85), .B(new_n210), .C1(new_n568), .C2(new_n571), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n570), .B(new_n574), .C1(new_n577), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n189), .A2(G227), .ZN(new_n582));
  XOR2_X1   g396(.A(G110), .B(G140), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n564), .B(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n562), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n210), .ZN(new_n588));
  INV_X1    g402(.A(new_n584), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n570), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n590), .A3(G469), .ZN(new_n591));
  NAND2_X1  g405(.A1(G469), .A2(G902), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n563), .B1(new_n586), .B2(new_n562), .ZN(new_n594));
  INV_X1    g408(.A(new_n570), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n584), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n572), .A2(new_n573), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n579), .A3(new_n578), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n598), .A2(new_n570), .A3(new_n589), .A4(new_n574), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n188), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G469), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n561), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n309), .A2(new_n494), .A3(new_n559), .A4(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(new_n324), .Z(G3));
  NAND2_X1  g419(.A1(new_n301), .A2(new_n187), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n606), .A2(G472), .B1(new_n302), .B2(new_n301), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n559), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n472), .A2(KEYINPUT33), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n472), .A2(KEYINPUT33), .ZN(new_n611));
  OAI211_X1 g425(.A(G478), .B(new_n187), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n470), .A2(new_n471), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n434), .B1(new_n613), .B2(new_n188), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n426), .B2(new_n427), .ZN(new_n616));
  OAI22_X1  g430(.A1(new_n491), .A2(new_n492), .B1(new_n616), .B2(new_n431), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n383), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(KEYINPUT93), .B(new_n310), .C1(new_n381), .C2(new_n382), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n479), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n609), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  OAI21_X1  g440(.A(KEYINPUT95), .B1(new_n491), .B2(KEYINPUT94), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n628), .B(new_n629), .C1(new_n489), .C2(new_n490), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n627), .A2(new_n492), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n492), .B1(new_n627), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n473), .A2(new_n474), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n433), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n609), .A2(new_n623), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(new_n310), .ZN(new_n640));
  INV_X1    g454(.A(new_n382), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n367), .A2(new_n379), .A3(new_n380), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n493), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n603), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(G472), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n301), .B2(new_n187), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n526), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n538), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n556), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n648), .A2(new_n652), .A3(new_n307), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  AND2_X1   g470(.A1(new_n556), .A2(new_n651), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n306), .B2(new_n308), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n603), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n621), .A2(new_n622), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n477), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n476), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR4_X1   g480(.A1(new_n631), .A2(new_n632), .A3(new_n635), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n660), .A2(new_n661), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  XNOR2_X1  g483(.A(new_n665), .B(KEYINPUT39), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n603), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  INV_X1    g486(.A(KEYINPUT97), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n301), .A2(new_n305), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n285), .A2(new_n250), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n194), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n251), .A2(new_n252), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n429), .B1(new_n680), .B2(new_n194), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n308), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT96), .Z(new_n684));
  NOR2_X1   g498(.A1(new_n381), .A2(new_n382), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT38), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n617), .A2(new_n634), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n686), .A2(new_n640), .A3(new_n652), .A4(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n674), .A2(new_n675), .A3(new_n684), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NOR2_X1   g504(.A1(new_n618), .A2(new_n666), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n660), .A2(new_n661), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NAND2_X1  g507(.A1(new_n556), .A2(new_n557), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n495), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT80), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n308), .B2(new_n306), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n600), .A2(new_n601), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n602), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n561), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n698), .A2(new_n619), .A3(new_n623), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND4_X1  g518(.A1(new_n698), .A2(new_n636), .A3(new_n623), .A4(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NAND4_X1  g520(.A1(new_n661), .A2(new_n658), .A3(new_n644), .A4(new_n701), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT98), .B(G119), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G21));
  INV_X1    g523(.A(new_n479), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n699), .A2(new_n560), .A3(new_n602), .A4(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n294), .A2(new_n300), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n253), .A2(new_n255), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n296), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n303), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n711), .A2(new_n715), .A3(new_n694), .A4(new_n647), .ZN(new_n716));
  INV_X1    g530(.A(new_n687), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT99), .B1(new_n661), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT99), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n719), .B(new_n687), .C1(new_n621), .C2(new_n622), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n723), .B(new_n716), .C1(new_n718), .C2(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND2_X1  g540(.A1(new_n661), .A2(new_n701), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n715), .A2(new_n647), .A3(new_n657), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n691), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n590), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n585), .A2(new_n590), .ZN(new_n735));
  OAI211_X1 g549(.A(G469), .B(new_n734), .C1(new_n735), .C2(new_n733), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n592), .B(KEYINPUT101), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n600), .B2(new_n601), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n561), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n381), .A2(new_n382), .A3(new_n640), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n309), .A2(new_n740), .A3(new_n559), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n691), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n732), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT103), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n746), .B(new_n732), .C1(new_n742), .C2(new_n743), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n308), .A2(KEYINPUT104), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n306), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n308), .A2(KEYINPUT104), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n694), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n740), .A2(new_n741), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(KEYINPUT42), .A3(new_n691), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  INV_X1    g570(.A(new_n667), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n742), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n201), .ZN(G36));
  OAI21_X1  g573(.A(new_n734), .B1(new_n735), .B2(new_n733), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(G469), .B1(new_n735), .B2(KEYINPUT45), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n738), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n602), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(KEYINPUT105), .A3(new_n602), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n765), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT106), .B1(new_n765), .B2(KEYINPUT46), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n560), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n670), .ZN(new_n775));
  INV_X1    g589(.A(new_n617), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n615), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT43), .Z(new_n778));
  INV_X1    g592(.A(new_n607), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n652), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  INV_X1    g597(.A(new_n741), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n775), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  NAND2_X1  g601(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n773), .A2(new_n560), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n743), .A2(new_n309), .A3(new_n559), .A4(new_n784), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(KEYINPUT107), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(new_n684), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n700), .A2(KEYINPUT49), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n700), .A2(KEYINPUT49), .ZN(new_n802));
  INV_X1    g616(.A(new_n694), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n560), .A3(new_n310), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n801), .A2(new_n802), .A3(new_n777), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n686), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n702), .A2(new_n705), .A3(new_n707), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n722), .B2(new_n724), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n310), .B(new_n710), .C1(new_n381), .C2(new_n382), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n618), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n559), .A3(new_n603), .A4(new_n607), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n604), .A3(KEYINPUT108), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT108), .B1(new_n811), .B2(new_n604), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n617), .A2(new_n633), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n643), .A2(new_n815), .A3(new_n710), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n608), .A2(new_n816), .B1(new_n645), .B2(new_n653), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT109), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT109), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n811), .A2(new_n604), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n819), .B1(new_n822), .B2(new_n812), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n808), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n753), .A2(new_n691), .A3(new_n728), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n433), .A2(new_n633), .A3(new_n665), .ZN(new_n826));
  OR4_X1    g640(.A1(new_n631), .A2(new_n784), .A3(new_n632), .A4(new_n826), .ZN(new_n827));
  OAI221_X1 g641(.A(new_n825), .B1(new_n757), .B2(new_n742), .C1(new_n827), .C2(new_n659), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n755), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT110), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n822), .A2(new_n812), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT109), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n822), .A2(new_n819), .A3(new_n812), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n828), .B1(new_n748), .B2(new_n754), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT110), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n808), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n668), .A2(new_n692), .A3(new_n730), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n718), .A2(new_n720), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n657), .A2(new_n683), .A3(new_n665), .A4(new_n740), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(KEYINPUT111), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT111), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT52), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n845), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n840), .A4(new_n843), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n668), .A2(new_n730), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n853), .B2(KEYINPUT52), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT53), .B1(new_n839), .B2(new_n851), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT54), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(KEYINPUT112), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n850), .B1(new_n831), .B2(new_n838), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n861), .B2(KEYINPUT53), .ZN(new_n862));
  INV_X1    g676(.A(new_n824), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n858), .B1(new_n853), .B2(KEYINPUT52), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n851), .A2(new_n863), .A3(new_n836), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n857), .B1(new_n866), .B2(KEYINPUT54), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n701), .A2(new_n741), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT115), .Z(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n476), .A3(new_n778), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n728), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n715), .A2(new_n647), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n803), .A2(new_n778), .A3(new_n476), .A4(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n686), .A2(new_n640), .A3(new_n701), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT50), .Z(new_n881));
  AND4_X1   g695(.A1(new_n559), .A2(new_n869), .A3(new_n476), .A4(new_n800), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n776), .A3(new_n614), .A4(new_n612), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n873), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n788), .B(new_n791), .C1(new_n560), .C2(new_n700), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n875), .A2(new_n741), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT113), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT51), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n872), .A2(new_n752), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT48), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n882), .A2(new_n619), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n475), .B(KEYINPUT117), .Z(new_n894));
  INV_X1    g708(.A(new_n727), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n875), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT51), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n867), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n900), .A2(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n806), .B1(new_n902), .B2(new_n903), .ZN(G75));
  NAND2_X1  g718(.A1(new_n866), .A2(new_n188), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(new_n380), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n351), .A2(new_n366), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n364), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(G952), .B2(new_n189), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT56), .B1(new_n906), .B2(KEYINPUT119), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(KEYINPUT119), .B2(new_n906), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n914), .B2(new_n909), .ZN(G51));
  NOR2_X1   g729(.A1(new_n189), .A2(G952), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n596), .A2(new_n599), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT120), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n866), .B(KEYINPUT54), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n737), .B(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n905), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n764), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n916), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n488), .A2(new_n427), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n926), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n916), .ZN(G60));
  OR2_X1    g745(.A1(new_n610), .A2(new_n611), .ZN(new_n932));
  XOR2_X1   g746(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n933));
  NOR2_X1   g747(.A1(new_n434), .A2(new_n429), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n916), .B1(new_n919), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n867), .A2(new_n935), .ZN(new_n938));
  INV_X1    g752(.A(new_n932), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n937), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT60), .Z(new_n947));
  AND3_X1   g761(.A1(new_n866), .A2(KEYINPUT123), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT123), .B1(new_n866), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n650), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n865), .B1(new_n856), .B2(KEYINPUT112), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n861), .A2(new_n860), .A3(KEYINPUT53), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n531), .A2(new_n536), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n866), .A2(KEYINPUT123), .A3(new_n947), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n916), .B1(KEYINPUT124), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n950), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n950), .A2(new_n958), .A3(new_n964), .A4(new_n960), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(G66));
  INV_X1    g780(.A(new_n361), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n967), .B2(new_n478), .ZN(new_n968));
  INV_X1    g782(.A(new_n189), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n968), .B1(new_n863), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(G898), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n907), .B1(new_n971), .B2(new_n969), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n970), .B(new_n972), .Z(G69));
  AOI21_X1  g787(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n796), .A2(new_n797), .B1(new_n775), .B2(new_n785), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n689), .A2(new_n840), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT125), .Z(new_n980));
  INV_X1    g794(.A(new_n815), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n784), .B1(new_n981), .B2(new_n618), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n698), .A2(new_n982), .A3(new_n603), .A4(new_n670), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n977), .A2(new_n980), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n275), .B1(new_n278), .B2(new_n284), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(new_n485), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n969), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n976), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n189), .A2(G900), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n774), .A2(new_n670), .A3(new_n841), .A4(new_n752), .ZN(new_n991));
  INV_X1    g805(.A(new_n758), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n755), .A2(new_n991), .A3(new_n992), .A4(new_n840), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n798), .A2(new_n786), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n994), .B2(new_n189), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n987), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n969), .B1(new_n977), .B2(new_n993), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n998), .A2(KEYINPUT126), .A3(new_n990), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n975), .B(new_n989), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n995), .A2(new_n996), .ZN(new_n1002));
  OAI21_X1  g816(.A(KEYINPUT126), .B1(new_n998), .B2(new_n990), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1002), .A2(new_n1003), .A3(new_n987), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n975), .B1(new_n1004), .B2(new_n989), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1001), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n985), .B2(new_n824), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n679), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n994), .B2(new_n824), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n677), .A2(new_n194), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n916), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1008), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n679), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n855), .B2(new_n856), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1010), .A2(new_n1013), .A3(new_n1016), .ZN(G57));
endmodule


