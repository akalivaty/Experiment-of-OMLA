//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G155gat), .B(G162gat), .Z(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT2), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT73), .B(KEYINPUT2), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n207), .B1(new_n208), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G120gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(G120gat), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(G113gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT1), .B1(new_n229), .B2(new_n222), .ZN(new_n230));
  OAI22_X1  g029(.A1(new_n225), .A2(new_n228), .B1(new_n230), .B2(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n215), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n218), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n236));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n231), .B(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(new_n232), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n232), .A2(new_n231), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT4), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n239), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n239), .A3(new_n246), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n238), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n243), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n251), .A2(new_n235), .A3(new_n237), .A4(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n232), .B(new_n231), .ZN(new_n254));
  INV_X1    g053(.A(new_n237), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n236), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n206), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n260));
  INV_X1    g059(.A(new_n249), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(new_n247), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n257), .B(new_n205), .C1(new_n262), .C2(new_n238), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(KEYINPUT6), .B(new_n206), .C1(new_n250), .C2(new_n258), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n267), .A3(new_n271), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT71), .Z(new_n278));
  INV_X1    g077(.A(G169gat), .ZN(new_n279));
  INV_X1    g078(.A(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT23), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n288));
  MUX2_X1   g087(.A(G183gat), .B(new_n288), .S(G190gat), .Z(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  INV_X1    g089(.A(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n287), .A2(KEYINPUT64), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT64), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n283), .A2(new_n284), .A3(new_n286), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT26), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n299), .A3(new_n284), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n285), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT27), .B(G183gat), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n302), .A2(new_n303), .A3(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n305));
  AOI21_X1  g104(.A(G190gat), .B1(new_n305), .B2(KEYINPUT27), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT28), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n300), .B(new_n301), .C1(new_n304), .C2(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n290), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(KEYINPUT65), .B2(new_n290), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n287), .B1(new_n289), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n298), .B(new_n310), .C1(new_n295), .C2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(G226gat), .A3(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n314), .A2(new_n317), .B1(G226gat), .B2(G233gat), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT72), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n278), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n277), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n316), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G64gat), .B(G92gat), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n326), .B(new_n327), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n322), .B2(new_n324), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(KEYINPUT30), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n325), .A2(new_n333), .A3(new_n328), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n266), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT29), .B1(new_n216), .B2(new_n217), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(new_n277), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n276), .A2(KEYINPUT75), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n339), .B(new_n317), .C1(new_n277), .C2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n216), .B1(new_n341), .B2(new_n217), .ZN(new_n342));
  INV_X1    g141(.A(G228gat), .ZN(new_n343));
  INV_X1    g142(.A(G233gat), .ZN(new_n344));
  OAI22_X1  g143(.A1(new_n338), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT3), .B1(new_n277), .B2(new_n317), .ZN(new_n347));
  OAI221_X1 g146(.A(new_n346), .B1(new_n347), .B2(new_n216), .C1(new_n278), .C2(new_n337), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G22gat), .ZN(new_n350));
  INV_X1    g149(.A(G22gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G78gat), .B(G106gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT31), .B(G50gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(new_n345), .B2(new_n348), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(KEYINPUT76), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n358), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G227gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(new_n344), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n314), .A2(new_n241), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n314), .A2(new_n241), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT32), .ZN(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT69), .ZN(new_n373));
  INV_X1    g172(.A(G15gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G43gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n371), .B(new_n377), .C1(KEYINPUT33), .C2(new_n369), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n370), .A2(KEYINPUT32), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n369), .B2(KEYINPUT33), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n367), .A2(new_n366), .A3(new_n368), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT34), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n378), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n378), .B2(new_n381), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT70), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(new_n385), .B2(new_n383), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT36), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT36), .B1(new_n386), .B2(new_n387), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n363), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n264), .A2(new_n265), .A3(new_n329), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT37), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n328), .B1(new_n325), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n319), .A2(new_n278), .A3(new_n321), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n323), .B1(new_n316), .B2(new_n318), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT38), .B1(new_n401), .B2(KEYINPUT37), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  OR3_X1    g202(.A1(new_n396), .A2(new_n403), .A3(KEYINPUT79), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT79), .B1(new_n396), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(new_n397), .B2(new_n325), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT38), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(KEYINPUT80), .A3(KEYINPUT38), .ZN(new_n410));
  AND4_X1   g209(.A1(new_n404), .A2(new_n405), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n254), .A2(new_n255), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n234), .B1(new_n248), .B2(new_n249), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT39), .B(new_n412), .C1(new_n413), .C2(new_n237), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n235), .B1(new_n261), .B2(new_n247), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT39), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n255), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n205), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT40), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT78), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n205), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT40), .A4(new_n414), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n412), .A2(KEYINPUT39), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n415), .B2(new_n255), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n419), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n259), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n335), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n332), .A2(KEYINPUT77), .A3(new_n334), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n361), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n395), .B1(new_n411), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n433), .A2(new_n434), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT35), .B1(new_n359), .B2(new_n360), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n388), .A2(new_n390), .A3(new_n266), .A4(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n438), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n388), .A2(new_n390), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n266), .A2(new_n440), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n435), .A4(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n386), .A2(new_n387), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n361), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT35), .B1(new_n448), .B2(new_n336), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n437), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n351), .A2(G15gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n374), .A2(G22gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n454), .A3(new_n452), .ZN(new_n457));
  INV_X1    g256(.A(G1gat), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n456), .A2(new_n457), .B1(KEYINPUT16), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n457), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n460), .A2(new_n455), .A3(G1gat), .ZN(new_n461));
  OAI21_X1  g260(.A(G8gat), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(KEYINPUT16), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n460), .B2(new_n455), .ZN(new_n465));
  INV_X1    g264(.A(G8gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT21), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471));
  INV_X1    g270(.A(G57gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(G64gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(G64gat), .ZN(new_n474));
  INV_X1    g273(.A(G64gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(G71gat), .A2(G78gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G71gat), .A2(G78gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT92), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n482));
  INV_X1    g281(.A(new_n480), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(new_n478), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT9), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n481), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n480), .B(new_n479), .C1(new_n488), .C2(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n469), .B1(new_n470), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n470), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  XNOR2_X1  g293(.A(new_n491), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G127gat), .B(G155gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT94), .ZN(new_n497));
  NAND2_X1  g296(.A1(G231gat), .A2(G233gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(KEYINPUT93), .Z(new_n499));
  XNOR2_X1  g298(.A(new_n497), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G183gat), .B(G211gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n495), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G232gat), .A2(G233gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT95), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT41), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n507), .B(KEYINPUT96), .Z(new_n508));
  XOR2_X1   g307(.A(G134gat), .B(G162gat), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n512));
  INV_X1    g311(.A(G92gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT99), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT99), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G92gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n512), .A2(new_n514), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519));
  OAI211_X1 g318(.A(G85gat), .B(G92gat), .C1(new_n519), .C2(KEYINPUT97), .ZN(new_n520));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT97), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G99gat), .ZN(new_n525));
  INV_X1    g324(.A(G106gat), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT8), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G99gat), .B(G106gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n518), .A2(new_n524), .A3(new_n529), .A4(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT100), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(KEYINPUT100), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT14), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n543));
  NAND2_X1  g342(.A1(G29gat), .A2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT85), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(KEYINPUT83), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT83), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n376), .A2(G50gat), .ZN(new_n552));
  INV_X1    g351(.A(G50gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(G43gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT84), .B1(new_n553), .B2(G43gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT84), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n376), .A3(G50gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(G43gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n550), .A2(new_n555), .B1(new_n548), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n376), .A2(G50gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n562), .A3(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(KEYINPUT15), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n539), .A2(new_n541), .A3(new_n544), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n547), .A2(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n536), .B1(new_n567), .B2(KEYINPUT86), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n542), .A2(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n560), .A2(new_n548), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(new_n569), .A3(new_n546), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n566), .A3(new_n555), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT17), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n535), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n505), .A2(new_n506), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(new_n535), .B2(new_n573), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580));
  NOR3_X1   g379(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT17), .B1(new_n573), .B2(new_n574), .ZN(new_n583));
  AOI211_X1 g382(.A(KEYINPUT86), .B(new_n536), .C1(new_n571), .C2(new_n572), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n534), .B(new_n533), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n585), .B2(new_n578), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n511), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n580), .B1(new_n576), .B2(new_n579), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n582), .A3(new_n578), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n510), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n503), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n490), .B1(new_n532), .B2(new_n531), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n535), .B2(new_n490), .ZN(new_n594));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT101), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n490), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(new_n533), .B2(new_n534), .ZN(new_n601));
  INV_X1    g400(.A(new_n596), .ZN(new_n602));
  NOR4_X1   g401(.A1(new_n601), .A2(new_n593), .A3(new_n598), .A4(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n604), .A3(KEYINPUT103), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n601), .B2(new_n593), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n535), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n596), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT102), .B1(new_n594), .B2(new_n596), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(new_n603), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n605), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n604), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n613), .B1(new_n619), .B2(new_n609), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n592), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n469), .B1(new_n583), .B2(new_n584), .ZN(new_n624));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT88), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n468), .A2(new_n573), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n624), .A2(KEYINPUT18), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G113gat), .B(G141gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G169gat), .B(G197gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT89), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n567), .A2(new_n462), .A3(new_n467), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n627), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n626), .B(KEYINPUT13), .Z(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  AOI211_X1 g440(.A(KEYINPUT89), .B(new_n641), .C1(new_n627), .C2(new_n637), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n628), .B(new_n635), .C1(new_n640), .C2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT18), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT90), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(KEYINPUT90), .A3(new_n645), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n468), .A2(new_n573), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n462), .A2(new_n467), .B1(new_n572), .B2(new_n571), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n639), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT89), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n638), .A2(new_n636), .A3(new_n639), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n644), .A2(new_n645), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n628), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n647), .A2(new_n648), .B1(new_n634), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n623), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n451), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n266), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  INV_X1    g461(.A(new_n659), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G8gat), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n663), .A2(new_n435), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n466), .B1(new_n659), .B2(new_n439), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT42), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(KEYINPUT42), .B2(new_n666), .ZN(G1325gat));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n392), .A2(new_n670), .A3(new_n393), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n392), .B2(new_n393), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(G15gat), .B1(new_n663), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n374), .A3(new_n444), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n362), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT106), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(new_n591), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n437), .B2(new_n450), .ZN(new_n683));
  INV_X1    g482(.A(new_n503), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n657), .A2(new_n684), .A3(new_n621), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(G29gat), .A3(new_n266), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT45), .Z(new_n688));
  AND3_X1   g487(.A1(new_n442), .A2(new_n446), .A3(new_n449), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n429), .B1(new_n420), .B2(new_n424), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n362), .B1(new_n690), .B2(new_n439), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n404), .A2(new_n405), .A3(new_n409), .A4(new_n410), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n394), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n591), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n451), .A2(KEYINPUT44), .A3(new_n591), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n685), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n266), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n688), .A2(new_n700), .ZN(G1328gat));
  NOR3_X1   g500(.A1(new_n686), .A2(G36gat), .A3(new_n435), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT46), .ZN(new_n703));
  OAI21_X1  g502(.A(G36gat), .B1(new_n699), .B2(new_n435), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1329gat));
  AOI21_X1  g504(.A(new_n699), .B1(new_n393), .B2(new_n392), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n376), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n686), .A2(G43gat), .A3(new_n443), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n698), .A2(new_n673), .A3(new_n685), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n711), .B2(G43gat), .ZN(new_n712));
  OAI22_X1  g511(.A1(new_n707), .A2(new_n710), .B1(KEYINPUT47), .B2(new_n712), .ZN(G1330gat));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n696), .A2(new_n697), .A3(new_n362), .A4(new_n685), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n361), .A2(G50gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT107), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n686), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n714), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT48), .B1(new_n686), .B2(new_n719), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n698), .A2(KEYINPUT108), .A3(new_n362), .A4(new_n685), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n553), .B1(new_n715), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n722), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT109), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n728), .B(new_n722), .C1(new_n723), .C2(new_n725), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n721), .B1(new_n727), .B2(new_n729), .ZN(G1331gat));
  INV_X1    g529(.A(KEYINPUT90), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n655), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n634), .B1(new_n652), .B2(new_n653), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n628), .A3(new_n733), .A4(new_n648), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n656), .A2(new_n634), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR4_X1   g535(.A1(new_n736), .A2(new_n622), .A3(new_n503), .A4(new_n591), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n451), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n266), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n472), .ZN(G1332gat));
  INV_X1    g539(.A(new_n738), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n435), .B(KEYINPUT110), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT111), .Z(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  OR3_X1    g547(.A1(new_n738), .A2(G71gat), .A3(new_n443), .ZN(new_n749));
  OAI21_X1  g548(.A(G71gat), .B1(new_n738), .B2(new_n674), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g551(.A1(new_n741), .A2(new_n362), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g553(.A1(new_n512), .A2(new_n517), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n684), .A2(new_n736), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n622), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n696), .A2(new_n697), .A3(new_n660), .A4(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n694), .B2(new_n757), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n266), .A2(new_n755), .A3(new_n622), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n755), .A2(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT112), .Z(G1336gat));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n762), .A3(KEYINPUT113), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n768), .B(new_n760), .C1(new_n694), .C2(new_n757), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n743), .A2(G92gat), .A3(new_n622), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n767), .A2(KEYINPUT114), .A3(new_n769), .A4(new_n770), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n698), .A2(new_n439), .A3(new_n758), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n514), .A2(new_n516), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n773), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT52), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n698), .A2(new_n742), .A3(new_n758), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n776), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(new_n763), .B2(new_n770), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n783), .ZN(G1337gat));
  NAND4_X1  g583(.A1(new_n763), .A2(new_n525), .A3(new_n444), .A4(new_n621), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n698), .A2(new_n673), .A3(new_n758), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n525), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n698), .A2(new_n362), .A3(new_n758), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G106gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n361), .A2(G106gat), .A3(new_n622), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n767), .A2(new_n769), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT53), .B1(new_n763), .B2(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1339gat));
  NAND2_X1  g595(.A1(new_n607), .A2(new_n608), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n602), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n607), .A2(new_n596), .A3(new_n608), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n612), .B1(new_n609), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n605), .A2(new_n614), .A3(new_n617), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n736), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n626), .B1(new_n624), .B2(new_n627), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n638), .A2(new_n639), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n633), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n734), .A2(new_n621), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n591), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n734), .A2(new_n813), .A3(new_n810), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n734), .B2(new_n810), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n607), .A2(new_n596), .A3(new_n608), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n609), .A3(new_n801), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n801), .A3(new_n602), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n613), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n816), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n821), .A2(new_n591), .A3(new_n618), .A4(new_n806), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n814), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n503), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n623), .A2(new_n736), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n266), .A3(new_n362), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n444), .A3(new_n743), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n220), .A3(new_n657), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n447), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n742), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n736), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n831), .B1(new_n834), .B2(new_n220), .ZN(G1340gat));
  NOR3_X1   g634(.A1(new_n830), .A2(new_n223), .A3(new_n622), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n621), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n223), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n839), .A3(new_n684), .ZN(new_n840));
  OAI21_X1  g639(.A(G127gat), .B1(new_n830), .B2(new_n503), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1342gat));
  OR4_X1    g641(.A1(G134gat), .A2(new_n832), .A3(new_n439), .A4(new_n682), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n830), .B2(new_n682), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n828), .B2(new_n361), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n821), .A2(new_n618), .A3(new_n806), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n811), .B1(new_n657), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n682), .ZN(new_n852));
  INV_X1    g651(.A(new_n815), .ZN(new_n853));
  INV_X1    g652(.A(new_n822), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n734), .A2(new_n813), .A3(new_n810), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n684), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g656(.A(KEYINPUT57), .B(new_n362), .C1(new_n857), .C2(new_n825), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n743), .A2(new_n660), .A3(new_n393), .A4(new_n392), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n657), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n674), .A2(new_n362), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT116), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n828), .A2(new_n266), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n743), .A3(new_n866), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n657), .A2(G141gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n622), .B1(new_n860), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n827), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n824), .A2(KEYINPUT119), .A3(new_n826), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n362), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n848), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n858), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n827), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n362), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n873), .B(new_n883), .C1(new_n872), .C2(new_n860), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n871), .B1(new_n884), .B2(G148gat), .ZN(new_n885));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT59), .B(new_n886), .C1(new_n861), .C2(new_n621), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n621), .A2(new_n886), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n885), .A2(new_n887), .B1(new_n867), .B2(new_n888), .ZN(G1345gat));
  OAI21_X1  g688(.A(G155gat), .B1(new_n862), .B2(new_n503), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n684), .A2(new_n210), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n867), .B2(new_n891), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n862), .B2(new_n682), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n865), .A2(new_n866), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n435), .A2(new_n211), .A3(new_n591), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1347gat));
  OR3_X1    g695(.A1(new_n435), .A2(KEYINPUT120), .A3(new_n660), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT120), .B1(new_n435), .B2(new_n660), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n900), .A2(new_n361), .A3(new_n444), .A4(new_n827), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n279), .A3(new_n657), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n743), .A2(new_n448), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n828), .A2(new_n660), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n736), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n905), .A2(new_n910), .ZN(G1348gat));
  OAI21_X1  g710(.A(G176gat), .B1(new_n904), .B2(new_n622), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n280), .A3(new_n621), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n904), .B2(new_n503), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n503), .A2(new_n302), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n909), .A2(new_n292), .A3(new_n591), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n591), .A3(new_n903), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(G190gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n920), .B2(G190gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n926), .B(new_n919), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1351gat));
  NOR2_X1   g727(.A1(new_n864), .A2(new_n743), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n907), .ZN(new_n930));
  AOI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n736), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n899), .A2(new_n673), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n883), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n736), .A2(G197gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1352gat));
  INV_X1    g734(.A(G204gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n933), .B2(new_n621), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n929), .A2(new_n936), .A3(new_n621), .A4(new_n907), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT123), .ZN(G1353gat));
  NAND3_X1  g741(.A1(new_n930), .A2(new_n269), .A3(new_n684), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n880), .A2(new_n881), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n361), .B1(new_n827), .B2(new_n874), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n947), .B2(new_n876), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n684), .B(new_n932), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n883), .A2(new_n951), .A3(new_n684), .A4(new_n932), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n269), .B1(KEYINPUT125), .B2(new_n944), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n945), .ZN(new_n956));
  INV_X1    g755(.A(new_n954), .ZN(new_n957));
  AOI211_X1 g756(.A(new_n956), .B(new_n957), .C1(new_n950), .C2(new_n952), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n943), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n961), .B(new_n943), .C1(new_n955), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1354gat));
  AOI21_X1  g762(.A(G218gat), .B1(new_n930), .B2(new_n591), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT127), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n682), .A2(new_n270), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n933), .B2(new_n966), .ZN(G1355gat));
endmodule


