//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1312, new_n1313, new_n1314, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n207), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n210), .B(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G68), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(G50), .B(G58), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  NAND3_X1  g0039(.A1(new_n204), .A2(G13), .A3(G20), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT12), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(G20), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n246), .A2(G77), .B1(G20), .B2(new_n242), .ZN(new_n247));
  INV_X1    g0047(.A(G50), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n213), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n253), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G1), .B2(new_n205), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n244), .B(new_n254), .C1(new_n242), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT11), .B1(new_n251), .B2(new_n253), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT14), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G226), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G97), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G232), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n213), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n268), .A2(KEYINPUT66), .A3(new_n213), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  AND2_X1   g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(G274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n280), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n277), .A2(G238), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n271), .A2(new_n284), .A3(KEYINPUT13), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT13), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n281), .A2(new_n283), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n270), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n260), .B(G169), .C1(new_n285), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT13), .B1(new_n271), .B2(new_n284), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n286), .A3(new_n270), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G179), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n291), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n260), .B1(new_n294), .B2(G169), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n259), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n285), .A2(new_n288), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n259), .B1(new_n297), .B2(G190), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n261), .A2(G223), .A3(G1698), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n261), .A2(new_n262), .ZN(new_n304));
  INV_X1    g0104(.A(G222), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n302), .B1(new_n303), .B2(new_n261), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n269), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT67), .B(G226), .Z(new_n308));
  NAND3_X1  g0108(.A1(new_n277), .A2(new_n282), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n281), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G200), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT8), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n312), .A2(KEYINPUT68), .A3(G58), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(KEYINPUT68), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n246), .ZN(new_n316));
  INV_X1    g0116(.A(G58), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n248), .A2(new_n317), .A3(new_n242), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(G20), .B1(G150), .B2(new_n249), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n255), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n241), .A2(new_n248), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n256), .B2(new_n248), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT9), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n307), .A2(G190), .A3(new_n281), .A4(new_n309), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n320), .B2(new_n322), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n311), .A2(new_n324), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT71), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT72), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT10), .B1(new_n328), .B2(KEYINPUT72), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(KEYINPUT72), .B(KEYINPUT10), .C1(new_n328), .C2(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G244), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n277), .A2(new_n282), .ZN(new_n336));
  INV_X1    g0136(.A(G238), .ZN(new_n337));
  AND2_X1   g0137(.A1(KEYINPUT70), .A2(G107), .ZN(new_n338));
  NOR2_X1   g0138(.A1(KEYINPUT70), .A2(G107), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n265), .A2(new_n337), .B1(new_n261), .B2(new_n340), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n304), .A2(KEYINPUT69), .A3(new_n266), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT69), .B1(new_n304), .B2(new_n266), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n269), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n281), .B1(new_n335), .B2(new_n336), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(G179), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n246), .B1(G20), .B2(G77), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n314), .A2(new_n250), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n255), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n241), .A2(new_n303), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n256), .B2(new_n303), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(new_n346), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n344), .A2(new_n345), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n281), .B1(new_n336), .B2(new_n335), .ZN(new_n360));
  OAI21_X1  g0160(.A(G200), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n355), .C1(new_n362), .C2(new_n346), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n310), .A2(G179), .ZN(new_n364));
  INV_X1    g0164(.A(new_n323), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n310), .A2(new_n356), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n358), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n301), .A2(new_n334), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n249), .A2(G159), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT74), .ZN(new_n371));
  XNOR2_X1  g0171(.A(G58), .B(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n245), .ZN(new_n378));
  NAND2_X1  g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n205), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n378), .A2(KEYINPUT7), .A3(new_n205), .A4(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n376), .B1(new_n384), .B2(G68), .ZN(new_n385));
  AOI211_X1 g0185(.A(KEYINPUT73), .B(new_n242), .C1(new_n382), .C2(new_n383), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT16), .B(new_n375), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n242), .B1(new_n382), .B2(new_n383), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n374), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n390), .A3(new_n253), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n315), .A2(new_n241), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n315), .B2(new_n256), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT75), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(KEYINPUT75), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n277), .A2(G232), .A3(new_n282), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n281), .A2(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(G223), .A2(G1698), .ZN(new_n401));
  AND2_X1   g0201(.A1(KEYINPUT3), .A2(G33), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT3), .A2(G33), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n401), .B1(G226), .B2(new_n262), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n345), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n406), .B(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n400), .A2(G179), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n407), .A2(new_n356), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n397), .A2(new_n398), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n397), .A2(new_n414), .A3(new_n398), .A4(new_n411), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n299), .B1(new_n400), .B2(new_n406), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n406), .B(KEYINPUT76), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n281), .A2(new_n399), .A3(new_n362), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(new_n391), .A3(new_n394), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n419), .A2(new_n391), .A3(KEYINPUT17), .A4(new_n394), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n413), .A2(new_n415), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n369), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(G264), .B(G1698), .C1(new_n402), .C2(new_n403), .ZN(new_n427));
  OAI211_X1 g0227(.A(G257), .B(new_n262), .C1(new_n402), .C2(new_n403), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n378), .A2(G303), .A3(new_n379), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n269), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n204), .A2(G45), .ZN(new_n432));
  OR2_X1    g0232(.A1(KEYINPUT5), .A2(G41), .ZN(new_n433));
  NAND2_X1  g0233(.A1(KEYINPUT5), .A2(G41), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT66), .B1(new_n268), .B2(new_n213), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n274), .A2(new_n273), .A3(new_n275), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n435), .A2(G274), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n279), .A2(G1), .ZN(new_n439));
  INV_X1    g0239(.A(new_n434), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(new_n436), .A3(G270), .A4(new_n437), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n431), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G116), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n204), .A2(new_n445), .A3(G13), .A4(G20), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT80), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n204), .A2(G33), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n240), .A2(new_n449), .A3(new_n213), .A4(new_n252), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n252), .A2(new_n213), .B1(G20), .B2(new_n445), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n205), .C1(G33), .C2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(KEYINPUT20), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT20), .B1(new_n451), .B2(new_n454), .ZN(new_n457));
  OAI221_X1 g0257(.A(new_n448), .B1(new_n445), .B2(new_n450), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n444), .A2(new_n458), .A3(KEYINPUT81), .A4(G179), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n438), .A2(new_n443), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n431), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(new_n458), .A3(KEYINPUT21), .A4(G169), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n446), .A2(new_n447), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n446), .A2(new_n447), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n464), .A2(new_n465), .B1(new_n450), .B2(new_n445), .ZN(new_n466));
  INV_X1    g0266(.A(new_n457), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(new_n455), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n431), .A2(G179), .A3(new_n438), .A4(new_n443), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(new_n462), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT82), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n459), .A2(new_n462), .A3(new_n470), .A4(KEYINPUT82), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n461), .A2(new_n458), .A3(G169), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n458), .B1(new_n461), .B2(G200), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n362), .B2(new_n461), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n473), .A2(new_n474), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n205), .B(G87), .C1(new_n402), .C2(new_n403), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(KEYINPUT22), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n261), .A2(new_n205), .A3(G87), .A4(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(KEYINPUT22), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT23), .ZN(new_n491));
  INV_X1    g0291(.A(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(G20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n205), .A2(G33), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n445), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n340), .A2(G20), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(KEYINPUT23), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n489), .A2(new_n490), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n490), .B1(new_n489), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n253), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n450), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n241), .A2(KEYINPUT25), .A3(new_n492), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT25), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n240), .B2(G107), .ZN(new_n504));
  AOI22_X1  g0304(.A1(G107), .A2(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT84), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n277), .A2(new_n506), .A3(G264), .A4(new_n442), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n442), .A2(new_n436), .A3(G264), .A4(new_n437), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n261), .A2(G257), .A3(G1698), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n261), .A2(G250), .A3(new_n262), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G294), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n507), .A2(new_n509), .B1(new_n269), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n514), .A2(new_n362), .A3(new_n438), .ZN(new_n515));
  AOI21_X1  g0315(.A(G200), .B1(new_n514), .B2(new_n438), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n500), .B(new_n505), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(KEYINPUT4), .A2(G244), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n262), .B(new_n518), .C1(new_n402), .C2(new_n403), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n335), .B1(new_n378), .B2(new_n379), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n452), .C1(new_n520), .C2(KEYINPUT4), .ZN(new_n521));
  OAI21_X1  g0321(.A(G250), .B1(new_n402), .B2(new_n403), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n262), .B1(new_n522), .B2(KEYINPUT4), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n269), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n442), .A2(new_n436), .A3(G257), .A4(new_n437), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n525), .A2(KEYINPUT78), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(KEYINPUT78), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n524), .B(new_n438), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n530), .A2(new_n453), .A3(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(G97), .B(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n533), .A2(new_n205), .B1(new_n303), .B2(new_n250), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n340), .B1(new_n382), .B2(new_n383), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n253), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n450), .A2(G97), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n240), .A2(new_n453), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT77), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(KEYINPUT77), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n529), .B(new_n544), .C1(new_n362), .C2(new_n528), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n528), .A2(new_n356), .B1(new_n536), .B2(new_n543), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT78), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n525), .B(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G179), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n438), .A4(new_n524), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n517), .A2(new_n545), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n507), .A2(new_n509), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n513), .A2(new_n269), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n438), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n550), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n356), .B1(new_n514), .B2(new_n438), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n489), .A2(new_n497), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT24), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n489), .A2(new_n490), .A3(new_n497), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n255), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n505), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n557), .A2(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT70), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n492), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G87), .A2(G97), .ZN(new_n567));
  NAND2_X1  g0367(.A1(KEYINPUT70), .A2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n205), .B1(new_n264), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n205), .B(G68), .C1(new_n402), .C2(new_n403), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n570), .B1(new_n494), .B2(new_n453), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT79), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n571), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT79), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n574), .A4(new_n573), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n253), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n349), .A2(new_n240), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n501), .A2(G87), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G238), .B(new_n262), .C1(new_n402), .C2(new_n403), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(G1698), .C1(new_n402), .C2(new_n403), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G116), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n269), .ZN(new_n589));
  AOI21_X1  g0389(.A(G250), .B1(new_n204), .B2(G45), .ZN(new_n590));
  INV_X1    g0390(.A(G274), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n439), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n277), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(G190), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n588), .A2(new_n269), .B1(new_n277), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n299), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n589), .A2(new_n550), .A3(new_n593), .ZN(new_n598));
  AOI21_X1  g0398(.A(G169), .B1(new_n589), .B2(new_n593), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n450), .A2(new_n348), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n580), .A2(new_n602), .A3(new_n582), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n584), .A2(new_n597), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n564), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n553), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n426), .A2(new_n481), .A3(new_n606), .ZN(G372));
  INV_X1    g0407(.A(new_n367), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n395), .A2(new_n411), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(new_n414), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n300), .A2(new_n347), .A3(new_n357), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n611), .A2(new_n296), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n422), .A2(new_n423), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT88), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n334), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n332), .A2(KEYINPUT88), .A3(new_n333), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n608), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n426), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n600), .A2(new_n603), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT87), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n577), .A2(new_n574), .A3(new_n573), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n255), .B1(new_n624), .B2(KEYINPUT79), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n601), .B(new_n581), .C1(new_n625), .C2(new_n579), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n595), .A2(new_n550), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G169), .B2(new_n595), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n626), .A2(new_n628), .B1(new_n629), .B2(new_n596), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT26), .B1(new_n552), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n581), .B1(new_n625), .B2(new_n579), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n589), .A2(new_n593), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(KEYINPUT85), .A3(G200), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n595), .B2(new_n299), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n634), .A2(new_n636), .A3(new_n638), .A4(new_n583), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n594), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n636), .A2(new_n638), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT86), .B1(new_n642), .B2(new_n584), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n633), .B(new_n621), .C1(new_n641), .C2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n477), .A2(new_n459), .A3(new_n462), .A4(new_n470), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n556), .A2(G169), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n514), .A2(G179), .A3(new_n438), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(new_n500), .B2(new_n505), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n545), .B(new_n517), .C1(new_n646), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n552), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n632), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n619), .B1(new_n620), .B2(new_n652), .ZN(G369));
  NAND3_X1  g0453(.A1(new_n204), .A2(new_n205), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n468), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n646), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n480), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT89), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n564), .A2(new_n660), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT90), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n659), .B1(new_n562), .B2(new_n563), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n517), .A2(new_n564), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n471), .A2(new_n472), .B1(new_n476), .B2(new_n475), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n659), .B1(new_n673), .B2(new_n474), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n649), .A2(new_n660), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n208), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n569), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n211), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n621), .B1(new_n641), .B2(new_n643), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n553), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n473), .A2(new_n474), .A3(new_n564), .A4(new_n477), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT93), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT93), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n673), .A2(new_n692), .A3(new_n474), .A4(new_n564), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n552), .A2(new_n633), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n695), .B(new_n621), .C1(new_n641), .C2(new_n643), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n633), .B1(new_n552), .B2(new_n630), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n622), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n687), .B1(new_n699), .B2(new_n660), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n553), .A2(new_n605), .A3(new_n659), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT92), .A3(new_n481), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT92), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n649), .A2(new_n630), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n536), .A2(new_n543), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n524), .A2(new_n438), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n548), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n706), .B1(new_n708), .B2(G190), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(new_n529), .B1(new_n546), .B2(new_n551), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n705), .A2(new_n710), .A3(new_n517), .A4(new_n660), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n704), .B1(new_n711), .B2(new_n480), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n703), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n659), .A2(KEYINPUT31), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n469), .A2(new_n635), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n708), .A2(new_n715), .A3(KEYINPUT30), .A4(new_n514), .ZN(new_n716));
  AOI21_X1  g0516(.A(G179), .B1(new_n460), .B2(new_n431), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n556), .A2(new_n528), .A3(new_n635), .A4(new_n717), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n514), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n528), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n714), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT91), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n595), .A2(new_n460), .A3(G179), .A4(new_n431), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n554), .A2(new_n555), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n528), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n724), .B1(new_n727), .B2(KEYINPUT30), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT91), .B(new_n720), .C1(new_n721), .C2(new_n528), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n719), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n659), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n723), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n701), .B1(new_n713), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n652), .A2(KEYINPUT29), .A3(new_n659), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n700), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n686), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n204), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n681), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n666), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n664), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n213), .B1(G20), .B2(new_n356), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT95), .B1(new_n550), .B2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n205), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n550), .A2(KEYINPUT95), .A3(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n362), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G87), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n205), .A2(G190), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(G179), .A3(new_n299), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n205), .A2(new_n550), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(G190), .A3(new_n299), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n261), .B1(new_n759), .B2(new_n303), .C1(new_n317), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n758), .A2(new_n550), .A3(new_n299), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n763), .A2(KEYINPUT32), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT32), .ZN(new_n766));
  INV_X1    g0566(.A(new_n763), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(new_n767), .B2(G159), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n762), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n362), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n205), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n453), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n760), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(G68), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(new_n362), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n248), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n750), .A2(G190), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G107), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n757), .A2(new_n769), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n774), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  INV_X1    g0583(.A(G326), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n782), .A2(new_n783), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n761), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n261), .B1(new_n786), .B2(G322), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n771), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n759), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n767), .A2(G329), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n785), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  INV_X1    g0594(.A(new_n779), .ZN(new_n795));
  INV_X1    g0595(.A(G303), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n793), .B1(new_n794), .B2(new_n795), .C1(new_n796), .C2(new_n755), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n746), .B1(new_n781), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n742), .ZN(new_n799));
  OR3_X1    g0599(.A1(KEYINPUT94), .A2(G13), .A3(G33), .ZN(new_n800));
  OAI21_X1  g0600(.A(KEYINPUT94), .B1(G13), .B2(G33), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n745), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n402), .A2(new_n403), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n208), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n279), .B2(new_n212), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n235), .B2(new_n279), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n680), .A2(new_n807), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n811), .A2(G355), .B1(new_n445), .B2(new_n680), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n798), .A2(new_n799), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n804), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n664), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n744), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n777), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G150), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n782), .A2(new_n821), .B1(new_n764), .B2(new_n759), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G143), .C2(new_n786), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n779), .A2(G68), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n261), .B1(new_n771), .B2(new_n317), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G132), .B2(new_n767), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n755), .A2(new_n248), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n755), .A2(new_n492), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n261), .B(new_n772), .C1(G294), .C2(new_n786), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n779), .A2(G87), .ZN(new_n833));
  INV_X1    g0633(.A(new_n759), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n776), .A2(G303), .B1(new_n834), .B2(G116), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n774), .A2(G283), .B1(new_n767), .B2(G311), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n745), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n802), .A2(new_n745), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n839), .B(new_n742), .C1(G77), .C2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n659), .B1(new_n352), .B2(new_n354), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n363), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n358), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n347), .A2(new_n357), .A3(new_n660), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n842), .B1(new_n802), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n847), .B(KEYINPUT97), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n652), .A2(new_n659), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n363), .A2(new_n843), .B1(new_n347), .B2(new_n357), .ZN(new_n852));
  INV_X1    g0652(.A(new_n846), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n851), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n742), .B1(new_n855), .B2(new_n734), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(KEYINPUT98), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n734), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n856), .B2(KEYINPUT98), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n848), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n739), .A2(new_n204), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT31), .B1(new_n730), .B2(new_n659), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT104), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n713), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n259), .A2(new_n659), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n296), .A2(new_n300), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n296), .B2(new_n300), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n854), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n610), .A2(new_n424), .ZN(new_n879));
  INV_X1    g0679(.A(new_n657), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n397), .A2(new_n398), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n609), .A2(new_n420), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n397), .A2(new_n398), .A3(new_n880), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n412), .A2(new_n885), .A3(new_n886), .A4(new_n420), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT7), .B1(new_n807), .B2(new_n205), .ZN(new_n892));
  INV_X1    g0692(.A(new_n383), .ZN(new_n893));
  OAI21_X1  g0693(.A(G68), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT73), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n389), .A2(new_n376), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n374), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n897), .A2(KEYINPUT16), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n255), .B1(new_n897), .B2(KEYINPUT16), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n393), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n657), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n425), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n420), .B1(new_n900), .B2(new_n657), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n407), .A2(new_n356), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n409), .A2(new_n410), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n890), .B1(new_n887), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT103), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n902), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n902), .B2(new_n909), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n891), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n703), .A2(new_n712), .B1(new_n868), .B2(KEYINPUT104), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n874), .B1(new_n914), .B2(new_n867), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT105), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n878), .A2(new_n913), .A3(new_n916), .A4(KEYINPUT40), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n902), .A2(new_n909), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n425), .A2(new_n901), .B1(new_n887), .B2(new_n908), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(KEYINPUT38), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n915), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n870), .A2(new_n426), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n701), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n610), .A2(new_n880), .ZN(new_n928));
  INV_X1    g0728(.A(new_n872), .ZN(new_n929));
  INV_X1    g0729(.A(new_n873), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n644), .B1(new_n552), .B2(new_n650), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n660), .B(new_n854), .C1(new_n932), .C2(new_n632), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n846), .B(KEYINPUT101), .Z(new_n934));
  AND3_X1   g0734(.A1(new_n933), .A2(KEYINPUT102), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT102), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n920), .B(new_n931), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n901), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n613), .B1(KEYINPUT18), .B2(new_n412), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n939), .B2(new_n415), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n887), .A2(new_n908), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n890), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT38), .B1(new_n882), .B2(new_n888), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n887), .A2(new_n908), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT38), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT103), .B1(new_n946), .B2(new_n940), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n902), .A2(new_n909), .A3(new_n910), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n943), .B1(new_n949), .B2(KEYINPUT39), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n296), .A2(new_n659), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n928), .B(new_n937), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n426), .B1(new_n700), .B2(new_n735), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n619), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n863), .B1(new_n927), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n927), .ZN(new_n957));
  INV_X1    g0757(.A(new_n533), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(G116), .A3(new_n214), .A4(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n248), .A2(G68), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT100), .Z(new_n965));
  AOI211_X1 g0765(.A(new_n303), .B(new_n211), .C1(G58), .C2(G68), .ZN(new_n966));
  OAI211_X1 g0766(.A(G1), .B(new_n738), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n957), .A2(new_n963), .A3(new_n967), .ZN(G367));
  OAI21_X1  g0768(.A(new_n805), .B1(new_n208), .B2(new_n348), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n231), .A2(new_n808), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n742), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n756), .A2(G58), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n779), .A2(G77), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n261), .B1(new_n761), .B2(new_n821), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G159), .B2(new_n774), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n771), .A2(new_n242), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n763), .A2(new_n819), .B1(new_n759), .B2(new_n248), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(G143), .C2(new_n776), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n972), .A2(new_n973), .A3(new_n975), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n756), .A2(G116), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT46), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n980), .A2(new_n981), .B1(G294), .B2(new_n774), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n981), .B2(new_n980), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT113), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n261), .B1(new_n767), .B2(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n794), .B2(new_n759), .C1(new_n340), .C2(new_n771), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n779), .A2(G97), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n777), .A2(new_n790), .B1(new_n796), .B2(new_n761), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(KEYINPUT112), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(KEYINPUT112), .C2(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n983), .B2(new_n984), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n979), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n971), .B1(new_n994), .B2(new_n745), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n629), .A2(new_n659), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT106), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n622), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT107), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT107), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n688), .C2(new_n997), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n995), .B1(new_n815), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n710), .B1(new_n544), .B2(new_n660), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT108), .Z(new_n1004));
  NAND3_X1  g0804(.A1(new_n546), .A2(new_n551), .A3(new_n659), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n677), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT45), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1007), .B2(new_n677), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1010), .A2(new_n1014), .A3(new_n672), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n672), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n675), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n666), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1022), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n665), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n671), .A2(new_n674), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1023), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1017), .A2(KEYINPUT110), .A3(new_n1018), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1020), .A2(new_n736), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n736), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n681), .B(KEYINPUT41), .Z(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n741), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1006), .A2(new_n671), .A3(new_n674), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT42), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n552), .B1(new_n1004), .B2(new_n564), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n660), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1038), .A2(KEYINPUT42), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT109), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1001), .B(KEYINPUT43), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(KEYINPUT109), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n672), .A2(new_n1007), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1002), .B1(new_n1037), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT114), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(G387));
  AOI21_X1  g0857(.A(new_n682), .B1(new_n1031), .B2(new_n736), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n736), .B2(new_n1031), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n668), .A2(new_n670), .A3(new_n804), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n228), .A2(new_n279), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n811), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1061), .A2(new_n808), .B1(new_n683), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n314), .A2(G50), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  AOI21_X1  g0865(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n683), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1063), .A2(new_n1067), .B1(new_n492), .B2(new_n680), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n742), .B1(new_n1068), .B2(new_n806), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n261), .B1(new_n248), .B2(new_n761), .C1(new_n777), .C2(new_n764), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n771), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n349), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n242), .B2(new_n759), .C1(new_n821), .C2(new_n763), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1070), .B(new_n1073), .C1(new_n315), .C2(new_n774), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1074), .B(new_n988), .C1(new_n303), .C2(new_n755), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT115), .Z(new_n1076));
  AOI22_X1  g0876(.A1(new_n774), .A2(G311), .B1(new_n776), .B2(G322), .ZN(new_n1077));
  INV_X1    g0877(.A(G317), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1077), .B1(new_n796), .B2(new_n759), .C1(new_n1078), .C2(new_n761), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT48), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n794), .B2(new_n771), .C1(new_n788), .C2(new_n755), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT49), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n807), .B1(new_n784), .B2(new_n763), .C1(new_n795), .C2(new_n445), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1076), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT116), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n746), .B1(new_n1087), .B2(KEYINPUT116), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1069), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1031), .A2(new_n741), .B1(new_n1060), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1059), .A2(new_n1091), .ZN(G393));
  NAND2_X1  g0892(.A1(new_n1007), .A2(new_n804), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n805), .B1(new_n453), .B2(new_n208), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n238), .A2(new_n808), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n742), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n771), .A2(new_n303), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G50), .B2(new_n774), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n314), .B2(new_n759), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n807), .B(new_n1099), .C1(G143), .C2(new_n767), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n777), .A2(new_n821), .B1(new_n764), .B2(new_n761), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT51), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1103), .A2(new_n833), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1100), .B(new_n1105), .C1(new_n242), .C2(new_n755), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G116), .A2(new_n1071), .B1(new_n774), .B2(G303), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n788), .B2(new_n759), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n261), .B(new_n1108), .C1(G322), .C2(new_n767), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n777), .A2(new_n1078), .B1(new_n790), .B2(new_n761), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT52), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1110), .A2(new_n1111), .B1(G107), .B2(new_n779), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1109), .B(new_n1112), .C1(new_n1111), .C2(new_n1110), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n755), .A2(new_n794), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1106), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1096), .B1(new_n1115), .B2(new_n745), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1093), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1019), .A2(new_n1015), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n740), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT117), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n1117), .C1(new_n1118), .C2(new_n740), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1031), .A2(new_n736), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1033), .A2(new_n681), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1126), .ZN(G390));
  AOI21_X1  g0927(.A(new_n701), .B1(new_n914), .B2(new_n867), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT92), .B1(new_n702), .B2(new_n481), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n711), .A2(new_n704), .A3(new_n480), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n733), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(G330), .A3(new_n854), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n931), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n875), .A2(new_n1128), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n935), .A2(new_n936), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n931), .B1(new_n1128), .B2(new_n849), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1131), .A2(new_n931), .A3(G330), .A4(new_n854), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n659), .B1(new_n694), .B2(new_n698), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n853), .B1(new_n1138), .B2(new_n845), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT118), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n870), .A2(new_n426), .A3(G330), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n953), .A2(new_n619), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1128), .A2(new_n875), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n933), .A2(new_n934), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT102), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n933), .A2(KEYINPUT102), .A3(new_n934), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n870), .A2(new_n849), .A3(G330), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1133), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1149), .A2(new_n1154), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT118), .B1(new_n1158), .B2(new_n1144), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT39), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n913), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1161), .A2(new_n943), .B1(new_n951), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1137), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1138), .A2(new_n845), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n846), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n931), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1167), .A2(new_n951), .A3(new_n913), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1163), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1162), .A2(new_n951), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n950), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n951), .A3(new_n913), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1147), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1146), .B(new_n1159), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n942), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1160), .B2(new_n913), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n951), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1154), .B2(new_n931), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1137), .B(new_n1172), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n870), .A2(new_n875), .A3(G330), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n931), .B1(new_n734), .B2(new_n854), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1154), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(KEYINPUT118), .B(new_n1144), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1142), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1179), .B(new_n1181), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1174), .A2(new_n1187), .A3(new_n681), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n949), .A2(new_n1177), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n950), .A2(new_n1170), .B1(new_n1189), .B2(new_n1167), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1179), .B(new_n741), .C1(new_n1147), .C2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n742), .B1(new_n315), .B2(new_n841), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n261), .B(new_n1097), .C1(G116), .C2(new_n786), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n777), .A2(new_n794), .B1(new_n763), .B2(new_n788), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n782), .A2(new_n340), .B1(new_n759), .B2(new_n453), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n757), .A2(new_n826), .A3(new_n1193), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n756), .A2(G150), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT53), .ZN(new_n1199));
  INV_X1    g0999(.A(G132), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n261), .B1(new_n761), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n774), .A2(G137), .B1(new_n776), .B2(G128), .ZN(new_n1202));
  INV_X1    g1002(.A(G125), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT54), .B(G143), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n763), .C1(new_n759), .C2(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1201), .B(new_n1205), .C1(G159), .C2(new_n1071), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n248), .B2(new_n795), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1197), .B1(new_n1199), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1192), .B1(new_n1208), .B2(new_n745), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1176), .B2(new_n803), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1191), .A2(KEYINPUT119), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT119), .B1(new_n1191), .B2(new_n1210), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1188), .B1(new_n1211), .B2(new_n1212), .ZN(G378));
  XNOR2_X1  g1013(.A(new_n1144), .B(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1159), .A2(new_n1146), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n701), .B1(new_n921), .B2(new_n922), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n323), .A2(new_n657), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT55), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n618), .B2(new_n367), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n608), .B(new_n1221), .C1(new_n616), .C2(new_n617), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n917), .A2(new_n1219), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n917), .B2(new_n1219), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n952), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n917), .A2(new_n1219), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1231), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n937), .A2(new_n928), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n917), .A2(new_n1219), .A3(new_n1231), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1234), .A2(new_n1241), .A3(KEYINPUT57), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n681), .B1(new_n1218), .B2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1179), .B1(new_n1190), .B2(new_n1147), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1214), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1234), .A2(new_n1241), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1243), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1234), .A2(new_n1241), .A3(new_n741), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n779), .A2(G58), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n278), .B(new_n807), .C1(new_n761), .C2(new_n492), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(new_n976), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n776), .A2(G116), .B1(new_n834), .B2(new_n349), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n774), .A2(G97), .B1(new_n767), .B2(G283), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n756), .B2(G77), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT58), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G33), .A2(G41), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT120), .ZN(new_n1260));
  AOI211_X1 g1060(.A(G50), .B(new_n1260), .C1(new_n278), .C2(new_n807), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT121), .Z(new_n1263));
  AOI22_X1  g1063(.A1(G150), .A2(new_n1071), .B1(new_n786), .B2(G128), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1203), .A2(new_n777), .B1(new_n782), .B2(new_n1200), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G137), .B2(new_n834), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(new_n755), .C2(new_n1204), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1267), .A2(KEYINPUT59), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n767), .A2(G124), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1260), .B(new_n1269), .C1(new_n795), .C2(new_n764), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT122), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1267), .B2(KEYINPUT59), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1268), .A2(new_n1272), .B1(KEYINPUT58), .B2(new_n1257), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n746), .B1(new_n1263), .B2(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n799), .B(new_n1274), .C1(new_n248), .C2(new_n840), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1236), .B2(new_n803), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1250), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1249), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(G375));
  NAND2_X1  g1080(.A1(new_n1133), .A2(new_n802), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n776), .A2(G132), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1282), .B1(new_n819), .B2(new_n761), .C1(new_n782), .C2(new_n1204), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n771), .A2(new_n248), .B1(new_n759), .B2(new_n821), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n807), .B(new_n1284), .C1(G128), .C2(new_n767), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1251), .B(new_n1285), .C1(new_n755), .C2(new_n764), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1283), .B1(new_n1286), .B2(KEYINPUT126), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(KEYINPUT126), .B2(new_n1286), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n782), .A2(new_n445), .B1(new_n759), .B2(new_n340), .ZN(new_n1289));
  XOR2_X1   g1089(.A(new_n1289), .B(KEYINPUT125), .Z(new_n1290));
  AOI22_X1  g1090(.A1(new_n776), .A2(G294), .B1(new_n767), .B2(G303), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n261), .B1(new_n786), .B2(G283), .ZN(new_n1292));
  AND4_X1   g1092(.A1(new_n973), .A2(new_n1291), .A3(new_n1072), .A4(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1290), .B(new_n1293), .C1(new_n453), .C2(new_n755), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n746), .B1(new_n1288), .B2(new_n1294), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n799), .B(new_n1295), .C1(new_n242), .C2(new_n840), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1141), .A2(new_n741), .B1(new_n1281), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1158), .A2(new_n1144), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(new_n1035), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1301), .B2(new_n1244), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(G381));
  NAND3_X1  g1103(.A1(new_n1059), .A2(new_n817), .A3(new_n1091), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1123), .A2(new_n1126), .A3(new_n1305), .A4(new_n861), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1191), .A2(new_n1210), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1188), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1306), .A2(G381), .A3(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1056), .A2(new_n1279), .A3(new_n1310), .ZN(G407));
  NAND2_X1  g1111(.A1(new_n658), .A2(G213), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1279), .A2(new_n1308), .A3(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(G407), .A2(G213), .A3(new_n1314), .ZN(G409));
  OR2_X1    g1115(.A1(new_n1037), .A2(new_n1053), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G393), .A2(G396), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1055), .B1(new_n1317), .B2(new_n1304), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(G390), .A2(new_n1318), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1123), .A2(new_n1126), .B1(new_n1317), .B2(new_n1304), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1316), .B(new_n1002), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1320), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1054), .B(new_n1322), .C1(G390), .C2(new_n1318), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G378), .B(new_n1277), .C1(new_n1243), .C2(new_n1248), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1246), .A2(new_n1036), .A3(new_n1247), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1277), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1308), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1313), .B1(new_n1325), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1300), .A2(KEYINPUT60), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n681), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1244), .A2(KEYINPUT60), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1331), .B1(new_n1332), .B2(new_n1299), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n861), .B1(new_n1333), .B2(new_n1298), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1333), .A2(new_n861), .A3(new_n1298), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT62), .B1(new_n1329), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT127), .B1(new_n1339), .B2(new_n1312), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  AOI211_X1 g1141(.A(new_n1341), .B(new_n1313), .C1(new_n1325), .C2(new_n1328), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1337), .A2(KEYINPUT62), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1338), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1336), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1346), .A2(G2897), .A3(new_n1313), .A4(new_n1334), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1313), .A2(G2897), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1348), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1350), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT61), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1324), .B1(new_n1345), .B2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1343), .A2(KEYINPUT63), .A3(new_n1337), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1324), .A2(KEYINPUT61), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT63), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1329), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1337), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1357), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1350), .A2(new_n1358), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1355), .A2(new_n1356), .A3(new_n1360), .A4(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1354), .A2(new_n1362), .ZN(G405));
  OAI21_X1  g1163(.A(new_n1325), .B1(new_n1279), .B2(new_n1309), .ZN(new_n1364));
  XNOR2_X1  g1164(.A(new_n1364), .B(new_n1337), .ZN(new_n1365));
  XNOR2_X1  g1165(.A(new_n1365), .B(new_n1324), .ZN(G402));
endmodule


