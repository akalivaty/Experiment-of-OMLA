//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT26), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT27), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT27), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(G183gat), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n214), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT27), .B(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n221), .A2(G183gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT68), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n228), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n227), .B1(KEYINPUT28), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n209), .A2(new_n210), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G169gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n215), .A2(new_n228), .A3(KEYINPUT64), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n239), .B(new_n244), .C1(new_n248), .C2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT23), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT25), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n245), .A2(new_n247), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n216), .A2(new_n218), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(G190gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n253), .A2(new_n254), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n203), .B1(new_n236), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G113gat), .ZN(new_n263));
  INV_X1    g062(.A(G120gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G113gat), .A2(G120gat), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268));
  XOR2_X1   g067(.A(G127gat), .B(G134gat), .Z(new_n269));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n268), .A3(new_n266), .ZN(new_n272));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n265), .A2(new_n266), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n273), .C1(new_n274), .C2(KEYINPUT69), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n254), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n260), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n229), .A2(new_n230), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT68), .B1(new_n232), .B2(new_n233), .ZN(new_n281));
  AOI21_X1  g080(.A(G190gat), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n226), .B(new_n214), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(KEYINPUT70), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n276), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G227gat), .ZN(new_n287));
  INV_X1    g086(.A(G233gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n276), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n279), .A2(KEYINPUT70), .A3(new_n284), .A4(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G15gat), .B(G43gat), .Z(new_n296));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n292), .B(KEYINPUT32), .C1(new_n294), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n291), .ZN(new_n304));
  INV_X1    g103(.A(new_n289), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT34), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT71), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n289), .B(new_n308), .C1(new_n286), .C2(new_n291), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n299), .A3(new_n301), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT72), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n310), .A2(new_n299), .A3(new_n316), .A4(new_n301), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n315), .B1(new_n314), .B2(new_n317), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n202), .B(new_n312), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321));
  INV_X1    g120(.A(G228gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(new_n288), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n324));
  NAND2_X1  g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328));
  AND2_X1   g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G211gat), .B(G218gat), .Z(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n324), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n330), .A2(new_n331), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n334), .A3(new_n327), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT74), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G155gat), .B(G162gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G141gat), .ZN(new_n344));
  INV_X1    g143(.A(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(KEYINPUT78), .A2(KEYINPUT79), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n346), .A2(new_n349), .A3(new_n350), .A4(new_n347), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n341), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n343), .A2(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G155gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT80), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G155gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n350), .B1(new_n359), .B2(G162gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n341), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT3), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n340), .B1(new_n363), .B2(KEYINPUT29), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT80), .B(G155gat), .ZN(new_n365));
  INV_X1    g164(.A(G162gat), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT2), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n353), .B1(new_n367), .B2(KEYINPUT79), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n341), .A2(new_n342), .ZN(new_n369));
  INV_X1    g168(.A(new_n348), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n369), .A2(new_n370), .B1(new_n351), .B2(new_n341), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT29), .B1(new_n337), .B2(new_n338), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g175(.A(KEYINPUT84), .B(KEYINPUT29), .C1(new_n337), .C2(new_n338), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n323), .B1(new_n364), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n354), .A2(new_n362), .A3(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n354), .A2(new_n362), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n332), .B2(new_n335), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n380), .B(new_n323), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n336), .A2(new_n339), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n373), .B1(new_n368), .B2(new_n371), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(G22gat), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT3), .B1(new_n383), .B2(KEYINPUT84), .ZN(new_n390));
  INV_X1    g189(.A(new_n377), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n381), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n392), .A2(new_n387), .B1(new_n322), .B2(new_n288), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n374), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n364), .A2(new_n380), .A3(new_n323), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G22gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n389), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n389), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n321), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT85), .B(G50gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n398), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n379), .A2(new_n388), .A3(G22gat), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n396), .B1(new_n393), .B2(new_n395), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n321), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n397), .A3(new_n398), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n401), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n402), .B1(new_n401), .B2(new_n409), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G8gat), .B(G36gat), .Z(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT77), .ZN(new_n414));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n280), .A2(new_n281), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n283), .B1(new_n418), .B2(new_n228), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT65), .B(G169gat), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n420), .A2(new_n240), .B1(new_n237), .B2(new_n238), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n258), .A2(new_n251), .A3(new_n249), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT25), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT66), .B(G183gat), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n424), .A2(new_n228), .B1(new_n245), .B2(new_n247), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n256), .ZN(new_n426));
  OAI22_X1  g225(.A1(new_n419), .A2(new_n227), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n382), .ZN(new_n428));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT75), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n429), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n279), .B2(new_n284), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n432), .B1(new_n433), .B2(new_n431), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n434), .B2(KEYINPUT75), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n417), .B1(new_n435), .B2(new_n385), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n427), .B2(new_n382), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n429), .B1(new_n279), .B2(new_n284), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT75), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n433), .B2(new_n431), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n439), .A2(new_n417), .A3(new_n385), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n434), .A2(new_n340), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n416), .B1(new_n436), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n439), .A2(new_n385), .A3(new_n441), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT76), .ZN(new_n447));
  INV_X1    g246(.A(new_n416), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n443), .A4(new_n442), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n444), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n448), .A4(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT0), .ZN(new_n456));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n380), .A2(new_n386), .A3(new_n290), .ZN(new_n460));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n276), .B1(new_n368), .B2(new_n371), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n276), .B(KEYINPUT4), .C1(new_n368), .C2(new_n371), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n460), .A2(new_n461), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n354), .A2(new_n362), .A3(new_n271), .A4(new_n275), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n462), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n461), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n372), .A2(new_n290), .A3(KEYINPUT81), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n466), .A2(new_n472), .A3(KEYINPUT5), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n460), .A2(new_n474), .A3(new_n461), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n464), .A2(new_n465), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n464), .A2(KEYINPUT82), .A3(new_n465), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n459), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n473), .A2(new_n480), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT6), .B1(new_n484), .B2(new_n458), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n454), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n412), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n314), .A2(new_n317), .B1(new_n311), .B2(new_n302), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n320), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n464), .A2(KEYINPUT82), .A3(new_n465), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT82), .B1(new_n464), .B2(new_n465), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n460), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n470), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n498), .A2(KEYINPUT86), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT86), .B1(new_n498), .B2(new_n499), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n499), .A3(new_n470), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(KEYINPUT40), .A3(new_n458), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n481), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT88), .B(new_n459), .C1(new_n473), .C2(new_n480), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n458), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT87), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n508), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n454), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n401), .A2(new_n409), .A3(new_n402), .ZN(new_n518));
  INV_X1    g317(.A(new_n402), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n399), .A2(new_n400), .A3(new_n321), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n447), .A2(new_n524), .A3(new_n443), .A4(new_n442), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n416), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n451), .B2(new_n447), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT38), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT90), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n435), .A2(new_n340), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n524), .B1(new_n434), .B2(new_n385), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT38), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(new_n525), .A3(new_n416), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n532), .A2(new_n525), .A3(KEYINPUT89), .A4(new_n416), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n485), .A2(new_n506), .A3(new_n507), .ZN(new_n538));
  INV_X1    g337(.A(new_n483), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n538), .A2(new_n539), .A3(new_n449), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n541), .B(KEYINPUT38), .C1(new_n526), .C2(new_n527), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n529), .A2(new_n537), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n518), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n490), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT35), .B1(new_n546), .B2(new_n488), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n314), .A2(new_n317), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT35), .B1(new_n538), .B2(new_n539), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n552), .A2(new_n454), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n551), .A2(new_n553), .A3(new_n545), .A4(new_n312), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n493), .A2(new_n544), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G8gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT16), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(G1gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n556), .B1(new_n559), .B2(KEYINPUT95), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(G1gat), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI221_X1 g361(.A(new_n559), .B1(KEYINPUT95), .B2(new_n556), .C1(G1gat), .C2(new_n557), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT92), .B(G29gat), .ZN(new_n565));
  INV_X1    g364(.A(G36gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(G29gat), .A2(G36gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT14), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G43gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G50gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT94), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT93), .B1(new_n571), .B2(G50gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n571), .A3(G50gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  INV_X1    g376(.A(G50gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(G43gat), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n573), .A2(new_n574), .A3(new_n576), .A4(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n572), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n571), .A2(G50gat), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n583), .A2(new_n584), .A3(new_n581), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n567), .B2(new_n569), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n564), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(KEYINPUT17), .A3(new_n588), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n591), .A2(new_n592), .B1(new_n589), .B2(new_n564), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT96), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n593), .A2(KEYINPUT98), .A3(KEYINPUT18), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(new_n590), .ZN(new_n597));
  INV_X1    g396(.A(new_n564), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n592), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n589), .A2(new_n564), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(KEYINPUT18), .A3(new_n595), .A4(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n595), .A3(new_n600), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n589), .B(new_n564), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n595), .B(KEYINPUT13), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n604), .A2(new_n608), .A3(new_n610), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT91), .B(G197gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT11), .B(G169gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n611), .B2(new_n613), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n622), .A2(new_n609), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n615), .A2(new_n621), .B1(new_n604), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n555), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G183gat), .B(G211gat), .Z(new_n626));
  INV_X1    g425(.A(G64gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  INV_X1    g427(.A(G57gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(KEYINPUT100), .A2(G57gat), .A3(G64gat), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT9), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n632), .A2(G71gat), .A3(G78gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(G71gat), .A2(G78gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n630), .B(new_n631), .C1(new_n633), .C2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n629), .A2(new_n627), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(G57gat), .A2(G64gat), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(KEYINPUT99), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(G71gat), .A3(G78gat), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n641), .B(new_n643), .C1(G71gat), .C2(G78gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n636), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT101), .ZN(new_n646));
  OAI211_X1 g445(.A(G231gat), .B(G233gat), .C1(new_n646), .C2(KEYINPUT21), .ZN(new_n647));
  XNOR2_X1  g446(.A(G127gat), .B(G155gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT20), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n645), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT21), .ZN(new_n653));
  NAND2_X1  g452(.A1(G231gat), .A2(G233gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n647), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n650), .B1(new_n647), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n626), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  INV_X1    g459(.A(new_n626), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n656), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n564), .B1(new_n646), .B2(KEYINPUT21), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n659), .A2(new_n662), .A3(new_n666), .ZN(new_n669));
  NAND2_X1  g468(.A1(G85gat), .A2(G92gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT7), .ZN(new_n671));
  NAND2_X1  g470(.A1(G99gat), .A2(G106gat), .ZN(new_n672));
  INV_X1    g471(.A(G85gat), .ZN(new_n673));
  INV_X1    g472(.A(G92gat), .ZN(new_n674));
  AOI22_X1  g473(.A1(KEYINPUT8), .A2(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(G99gat), .B(G106gat), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n671), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n597), .A2(new_n592), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  AND2_X1   g482(.A1(G232gat), .A2(G233gat), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n589), .A2(new_n683), .B1(KEYINPUT41), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(G190gat), .B(G218gat), .Z(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n684), .A2(KEYINPUT41), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT103), .ZN(new_n691));
  XNOR2_X1  g490(.A(G134gat), .B(G162gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n688), .B2(new_n689), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n668), .A2(new_n669), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n678), .A2(KEYINPUT10), .A3(new_n680), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n652), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n645), .A2(KEYINPUT101), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n645), .A2(KEYINPUT101), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n681), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n683), .A2(new_n645), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT10), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(G230gat), .A2(G233gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT104), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n698), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n709), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT10), .B1(new_n703), .B2(new_n704), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT105), .B(new_n711), .C1(new_n712), .C2(new_n700), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n705), .A2(new_n711), .ZN(new_n714));
  XNOR2_X1  g513(.A(G120gat), .B(G148gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(G176gat), .B(G204gat), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n715), .B(new_n716), .Z(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n710), .A2(new_n713), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n707), .A2(new_n709), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n721), .B2(new_n714), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n697), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n625), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n487), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n454), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT16), .B(G8gat), .Z(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n556), .B2(new_n729), .ZN(new_n732));
  MUX2_X1   g531(.A(new_n731), .B(new_n732), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g532(.A1(new_n320), .A2(new_n492), .ZN(new_n734));
  OAI21_X1  g533(.A(G15gat), .B1(new_n726), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n551), .A2(new_n312), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(G15gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n726), .B2(new_n737), .ZN(G1326gat));
  NOR2_X1   g537(.A1(new_n726), .A2(new_n545), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT43), .B(G22gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  NAND2_X1  g540(.A1(new_n668), .A2(new_n669), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n695), .A2(new_n696), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n742), .A2(new_n743), .A3(new_n723), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n625), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n486), .A3(new_n565), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT45), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n555), .B2(new_n743), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n554), .A2(new_n547), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n523), .A2(new_n543), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n320), .A2(new_n489), .A3(new_n492), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n743), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n723), .B(KEYINPUT106), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(new_n624), .A3(new_n742), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n749), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n749), .A2(new_n755), .A3(KEYINPUT107), .A4(new_n757), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n760), .A2(new_n486), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n747), .B1(new_n565), .B2(new_n762), .ZN(G1328gat));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n517), .A3(new_n761), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G36gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n625), .A2(new_n566), .A3(new_n517), .A4(new_n744), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT46), .Z(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n765), .A2(new_n767), .A3(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1329gat));
  OAI211_X1 g571(.A(KEYINPUT47), .B(G43gat), .C1(new_n758), .C2(new_n734), .ZN(new_n773));
  INV_X1    g572(.A(new_n736), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n745), .A2(new_n571), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n773), .B(new_n775), .C1(new_n776), .C2(KEYINPUT47), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  INV_X1    g577(.A(new_n734), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n779), .A3(new_n761), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(G43gat), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n777), .B1(new_n781), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g581(.A(KEYINPUT48), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n545), .A2(G50gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n625), .A2(new_n744), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n785), .B2(KEYINPUT111), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT112), .B1(new_n758), .B2(new_n545), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G50gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n758), .A2(KEYINPUT112), .A3(new_n545), .ZN(new_n789));
  OAI221_X1 g588(.A(new_n786), .B1(KEYINPUT111), .B2(new_n785), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n760), .A2(new_n412), .A3(new_n761), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n791), .A2(G50gat), .B1(new_n745), .B2(new_n784), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(G1331gat));
  NAND3_X1  g593(.A1(new_n756), .A2(new_n624), .A3(new_n697), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT113), .Z(new_n796));
  NAND2_X1  g595(.A1(new_n753), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n486), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G57gat), .ZN(G1332gat));
  INV_X1    g599(.A(new_n798), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n454), .ZN(new_n802));
  NOR2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  AND2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n802), .B2(new_n803), .ZN(G1333gat));
  OAI21_X1  g605(.A(G71gat), .B1(new_n801), .B2(new_n734), .ZN(new_n807));
  INV_X1    g606(.A(G71gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n798), .A2(new_n808), .A3(new_n774), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(KEYINPUT50), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1334gat));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n412), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g615(.A1(new_n749), .A2(new_n755), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n615), .A2(new_n621), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n623), .A2(new_n604), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n742), .A3(new_n724), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G85gat), .B1(new_n822), .B2(new_n487), .ZN(new_n823));
  INV_X1    g622(.A(new_n742), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n753), .A2(new_n624), .A3(new_n824), .A4(new_n754), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n486), .A2(new_n673), .A3(new_n723), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(G1336gat));
  OAI21_X1  g630(.A(G92gat), .B1(new_n822), .B2(new_n454), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n517), .A2(new_n674), .A3(new_n756), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT115), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n832), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n832), .B(new_n837), .C1(new_n829), .C2(new_n835), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1337gat));
  OAI21_X1  g640(.A(G99gat), .B1(new_n822), .B2(new_n734), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n736), .A2(G99gat), .A3(new_n724), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n829), .B2(new_n843), .ZN(G1338gat));
  NAND3_X1  g643(.A1(new_n817), .A2(new_n412), .A3(new_n821), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G106gat), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  INV_X1    g646(.A(new_n756), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n545), .A2(new_n848), .A3(G106gat), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n846), .B(new_n847), .C1(new_n829), .C2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n829), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n849), .B(KEYINPUT117), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n852), .A2(new_n853), .B1(new_n845), .B2(G106gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n854), .B2(new_n847), .ZN(G1339gat));
  NAND3_X1  g654(.A1(new_n697), .A2(new_n624), .A3(new_n724), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT118), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n707), .B2(new_n709), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n710), .A2(new_n859), .A3(new_n713), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n717), .B1(new_n721), .B2(new_n858), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n720), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n593), .A2(new_n595), .B1(new_n611), .B2(new_n613), .ZN(new_n864));
  INV_X1    g663(.A(new_n620), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n819), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT55), .B1(new_n860), .B2(new_n861), .ZN(new_n868));
  NOR4_X1   g667(.A1(new_n863), .A2(new_n867), .A3(new_n743), .A4(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n867), .A2(new_n724), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n624), .A2(new_n863), .ZN(new_n872));
  INV_X1    g671(.A(new_n868), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n870), .B1(new_n874), .B2(new_n754), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n857), .B1(new_n875), .B2(new_n824), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n412), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n517), .A2(new_n487), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n774), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G113gat), .B1(new_n879), .B2(new_n624), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n876), .A2(new_n487), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n546), .A2(new_n517), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n624), .A2(G113gat), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT119), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n883), .B2(new_n885), .ZN(G1340gat));
  NOR3_X1   g685(.A1(new_n879), .A2(new_n264), .A3(new_n848), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(new_n723), .A3(new_n882), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n264), .B2(new_n888), .ZN(G1341gat));
  OAI21_X1  g688(.A(G127gat), .B1(new_n879), .B2(new_n824), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n824), .A2(G127gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n883), .B2(new_n891), .ZN(G1342gat));
  NOR3_X1   g691(.A1(new_n883), .A2(G134gat), .A3(new_n743), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n879), .B2(new_n743), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  NOR2_X1   g697(.A1(new_n779), .A2(new_n545), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n881), .A2(new_n454), .A3(new_n899), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n900), .A2(new_n344), .A3(new_n820), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n734), .A2(new_n878), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT120), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n545), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n860), .A2(new_n861), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT55), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT121), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n863), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n820), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n871), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n754), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n907), .B(new_n824), .C1(new_n917), .C2(new_n869), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n856), .B(KEYINPUT118), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n871), .B1(new_n872), .B2(new_n913), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n870), .B1(new_n921), .B2(new_n754), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n907), .B1(new_n922), .B2(new_n824), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT123), .B(new_n906), .C1(new_n920), .C2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n905), .B1(new_n876), .B2(new_n545), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n915), .A2(new_n916), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n869), .B1(new_n927), .B2(new_n743), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT122), .B1(new_n928), .B2(new_n742), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n919), .A3(new_n918), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT123), .B1(new_n930), .B2(new_n906), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n904), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G141gat), .B1(new_n932), .B2(new_n624), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n902), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n936), .B(new_n904), .C1(new_n926), .C2(new_n931), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n820), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n901), .B1(new_n938), .B2(G141gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(G1344gat));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n723), .A3(new_n937), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n345), .A2(KEYINPUT59), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n876), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(KEYINPUT57), .A3(new_n412), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n856), .B1(new_n928), .B2(new_n742), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n412), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n946), .B1(KEYINPUT57), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(new_n723), .A3(new_n904), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT59), .B1(new_n950), .B2(new_n345), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n900), .A2(new_n345), .A3(new_n723), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1345gat));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n937), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n359), .B1(new_n955), .B2(new_n824), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n900), .A2(new_n365), .A3(new_n742), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1346gat));
  OAI21_X1  g757(.A(G162gat), .B1(new_n955), .B2(new_n743), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n900), .A2(new_n366), .A3(new_n754), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT125), .Z(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n454), .A2(new_n486), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n877), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n774), .ZN(new_n966));
  OAI21_X1  g765(.A(G169gat), .B1(new_n966), .B2(new_n624), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n964), .A2(new_n491), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n420), .A3(new_n820), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1348gat));
  OAI21_X1  g769(.A(G176gat), .B1(new_n966), .B2(new_n848), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n210), .A3(new_n723), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  OAI21_X1  g772(.A(new_n259), .B1(new_n966), .B2(new_n824), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n968), .A2(new_n418), .A3(new_n742), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n968), .A2(new_n228), .A3(new_n754), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n965), .A2(new_n774), .A3(new_n754), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n979), .A2(new_n980), .A3(G190gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n979), .B2(G190gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1351gat));
  AND2_X1   g782(.A1(new_n734), .A2(new_n963), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n949), .A2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(G197gat), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n985), .A2(new_n986), .A3(new_n624), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n945), .A2(new_n899), .A3(new_n963), .ZN(new_n988));
  AOI21_X1  g787(.A(G197gat), .B1(new_n988), .B2(new_n820), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(new_n989), .ZN(G1352gat));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n991));
  AOI21_X1  g790(.A(G204gat), .B1(new_n991), .B2(KEYINPUT62), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n988), .A2(new_n723), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n949), .A2(new_n756), .A3(new_n984), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(G204gat), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n996), .A2(KEYINPUT127), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(G1353gat));
  INV_X1    g799(.A(G211gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n988), .A2(new_n1001), .A3(new_n742), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n949), .A2(new_n742), .A3(new_n984), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(G1354gat));
  OAI21_X1  g805(.A(G218gat), .B1(new_n985), .B2(new_n743), .ZN(new_n1007));
  INV_X1    g806(.A(G218gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n988), .A2(new_n1008), .A3(new_n754), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1007), .A2(new_n1009), .ZN(G1355gat));
endmodule


