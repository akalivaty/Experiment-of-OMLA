//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT69), .B(G902), .Z(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT77), .ZN(new_n193));
  XNOR2_X1  g007(.A(G110), .B(G140), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT3), .B1(new_n197), .B2(G107), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n198), .A2(new_n201), .A3(KEYINPUT78), .A4(new_n202), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G101), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT79), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n197), .A2(KEYINPUT3), .A3(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n200), .A2(G104), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n211), .A2(KEYINPUT80), .A3(new_n212), .A4(new_n198), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n198), .A2(new_n201), .A3(new_n212), .A4(new_n202), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n205), .A2(new_n218), .A3(G101), .A4(new_n206), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n208), .A2(KEYINPUT4), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n205), .A2(new_n221), .A3(G101), .A4(new_n206), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT0), .A4(G128), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G128), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n200), .A2(G104), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n212), .B1(new_n234), .B2(new_n202), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n214), .A2(new_n215), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n214), .A2(new_n215), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n235), .B1(new_n213), .B2(new_n216), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT82), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT10), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n224), .A2(new_n226), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n225), .B2(G146), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(G128), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n224), .B(new_n226), .C1(KEYINPUT1), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(KEYINPUT66), .A3(new_n249), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n244), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n241), .A2(new_n243), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n247), .A2(new_n249), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n256), .B(KEYINPUT10), .C1(new_n242), .C2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n257), .B(new_n236), .C1(new_n237), .C2(new_n238), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT81), .B1(new_n259), .B2(new_n244), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n233), .B(new_n255), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G131), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n264), .A2(new_n267), .A3(new_n270), .A4(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n272), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT82), .B1(new_n217), .B2(new_n236), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n240), .B(new_n235), .C1(new_n213), .C2(new_n216), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n277), .A2(new_n254), .B1(new_n220), .B2(new_n232), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n259), .A2(new_n244), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n256), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n259), .A2(KEYINPUT81), .A3(new_n244), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n274), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n196), .B1(new_n273), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n239), .A2(new_n250), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n259), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT12), .B1(new_n286), .B2(new_n272), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT12), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n288), .B(new_n274), .C1(new_n285), .C2(new_n259), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT83), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n278), .A2(new_n282), .A3(new_n274), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n217), .A2(new_n257), .A3(new_n236), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n257), .B1(new_n217), .B2(new_n236), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n272), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n288), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT83), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n290), .A2(new_n291), .A3(new_n298), .A4(new_n195), .ZN(new_n299));
  AOI211_X1 g113(.A(G469), .B(new_n190), .C1(new_n284), .C2(new_n299), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n261), .A2(new_n272), .B1(new_n289), .B2(new_n287), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n196), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n261), .A2(new_n272), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n291), .A3(new_n195), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(G469), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(G469), .A2(G902), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n188), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT16), .ZN(new_n314));
  OR3_X1    g128(.A1(new_n312), .A2(KEYINPUT16), .A3(G140), .ZN(new_n315));
  AOI21_X1  g129(.A(G146), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(G237), .A2(G953), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(G143), .A3(G214), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(G143), .B1(new_n318), .B2(G214), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT17), .B(G131), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n314), .A2(new_n315), .A3(G146), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n317), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G131), .B1(new_n320), .B2(new_n321), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n327));
  INV_X1    g141(.A(G237), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n191), .A3(G214), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n225), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n270), .A3(new_n319), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n317), .A2(new_n322), .A3(new_n324), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT90), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT18), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n270), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n320), .B2(new_n321), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n311), .A2(new_n313), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G146), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n223), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n330), .B(new_n319), .C1(new_n337), .C2(new_n270), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT88), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n339), .A2(new_n344), .A3(new_n345), .A4(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n334), .A2(new_n336), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n197), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n347), .A2(new_n349), .ZN(new_n354));
  INV_X1    g168(.A(new_n336), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n354), .B(new_n352), .C1(new_n355), .C2(new_n333), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n309), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G475), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n342), .B(KEYINPUT19), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n360), .A2(new_n223), .B1(new_n326), .B2(new_n331), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n324), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT73), .A4(G146), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n352), .B1(new_n354), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT89), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n347), .A2(new_n349), .B1(new_n361), .B2(new_n365), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(new_n352), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n371), .A3(new_n356), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n372), .B2(new_n374), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n359), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G478), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n379), .A2(KEYINPUT15), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n248), .A2(G143), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT13), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n225), .A2(G128), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT92), .A3(new_n382), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT92), .B1(new_n383), .B2(new_n382), .ZN(new_n386));
  OAI221_X1 g200(.A(new_n381), .B1(new_n382), .B2(new_n383), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  INV_X1    g202(.A(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G116), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G122), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n200), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n390), .A2(new_n391), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT91), .B1(new_n389), .B2(G116), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G107), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n383), .A2(new_n381), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT93), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT93), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n383), .A2(new_n381), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n263), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n388), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n394), .A2(KEYINPUT14), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT94), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n394), .A2(KEYINPUT14), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n392), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G107), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n402), .A2(G134), .A3(new_n404), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n414), .A3(new_n395), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n187), .A2(new_n416), .A3(G953), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n407), .B2(new_n415), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n189), .B(new_n380), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n407), .A2(new_n415), .ZN(new_n423));
  INV_X1    g237(.A(new_n417), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n418), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n380), .B1(new_n426), .B2(new_n189), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n308), .A2(new_n378), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT65), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n230), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n227), .B(KEYINPUT65), .C1(new_n228), .C2(new_n229), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n272), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n265), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n263), .A2(G137), .ZN(new_n436));
  OAI21_X1  g250(.A(G131), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n271), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n257), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G116), .B(G119), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT2), .B(G113), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n446), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n444), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n247), .A2(KEYINPUT66), .A3(new_n249), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT66), .B1(new_n247), .B2(new_n249), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n439), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n231), .A2(new_n272), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(KEYINPUT30), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n443), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n457));
  NAND2_X1  g271(.A1(new_n318), .A2(G210), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT26), .B(G101), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n450), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n453), .A2(new_n462), .A3(new_n454), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n456), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT31), .ZN(new_n465));
  INV_X1    g279(.A(new_n461), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n441), .A2(new_n450), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n453), .A2(KEYINPUT28), .A3(new_n462), .A4(new_n454), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n466), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT31), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n456), .A2(new_n473), .A3(new_n461), .A4(new_n463), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(G472), .A2(G902), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT32), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n438), .B1(new_n252), .B2(new_n253), .ZN(new_n481));
  INV_X1    g295(.A(new_n454), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n450), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n463), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT68), .B(new_n450), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(KEYINPUT28), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n468), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n461), .A2(KEYINPUT29), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n461), .B1(new_n468), .B2(new_n471), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n456), .A2(new_n466), .A3(new_n463), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n490), .B(new_n189), .C1(new_n493), .C2(KEYINPUT29), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n478), .A2(new_n480), .B1(G472), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(KEYINPUT72), .A2(G110), .ZN(new_n496));
  NOR2_X1   g310(.A1(KEYINPUT72), .A2(G110), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n248), .B(G119), .C1(KEYINPUT71), .C2(KEYINPUT23), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n500));
  INV_X1    g314(.A(G119), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(G128), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n501), .B2(G128), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n498), .B(new_n499), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n501), .B2(G128), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(G128), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n248), .A2(KEYINPUT70), .A3(G119), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT24), .B(G110), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(new_n363), .A3(new_n364), .A4(new_n343), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n510), .A2(new_n511), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G110), .ZN(new_n517));
  INV_X1    g331(.A(new_n324), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n515), .B(new_n517), .C1(new_n518), .C2(new_n316), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT75), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT22), .B(G137), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT74), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n514), .A2(new_n519), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT76), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n514), .A3(new_n519), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n521), .A2(new_n532), .A3(new_n526), .A4(new_n528), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n530), .A2(new_n189), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT25), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n533), .A2(new_n531), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n537), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n530), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n416), .B1(new_n189), .B2(G234), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n530), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n542), .A2(G902), .A3(new_n540), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n495), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n191), .A2(G952), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(G234), .B2(G237), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n191), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT21), .B(G898), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G214), .B1(G237), .B2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G210), .B1(G237), .B2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n247), .A2(new_n312), .A3(new_n249), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n227), .B(G125), .C1(new_n228), .C2(new_n229), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n191), .A2(G224), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT85), .A3(KEYINPUT7), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT85), .B1(new_n560), .B2(KEYINPUT7), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n557), .B2(new_n558), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n565), .B2(new_n562), .ZN(new_n566));
  INV_X1    g380(.A(G113), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n393), .A2(G119), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT5), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n445), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n449), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n242), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G122), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT8), .Z(new_n576));
  OR2_X1    g390(.A1(new_n445), .A2(new_n568), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n577), .A2(new_n570), .B1(new_n444), .B2(new_n448), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n576), .B1(new_n578), .B2(new_n239), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n566), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n241), .A2(new_n243), .A3(new_n578), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n222), .A2(new_n450), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT4), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n212), .B1(new_n203), .B2(new_n204), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n218), .B1(new_n584), .B2(new_n206), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n581), .A2(new_n586), .A3(new_n575), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n556), .B1(new_n588), .B2(new_n309), .ZN(new_n589));
  AOI211_X1 g403(.A(KEYINPUT86), .B(G902), .C1(new_n580), .C2(new_n587), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n586), .ZN(new_n592));
  INV_X1    g406(.A(new_n575), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT6), .A3(new_n587), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n592), .A2(new_n596), .A3(new_n593), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n559), .B(new_n560), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n555), .B1(new_n591), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n601), .B(new_n554), .C1(new_n589), .C2(new_n590), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n551), .B(new_n553), .C1(new_n600), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n430), .A2(new_n546), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n475), .A2(new_n189), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n477), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n308), .A2(new_n545), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n609), .A2(new_n603), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n418), .B2(KEYINPUT95), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n426), .B(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n190), .A2(new_n379), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n426), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n379), .B1(new_n616), .B2(new_n190), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n378), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT96), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n377), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n372), .A2(new_n376), .A3(new_n374), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n429), .A3(new_n359), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n610), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n540), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n521), .A2(new_n528), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n634), .B(new_n635), .Z(new_n636));
  AOI22_X1  g450(.A1(new_n539), .A2(new_n540), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n608), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n430), .A2(new_n603), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G12));
  NOR2_X1   g456(.A1(new_n308), .A2(new_n495), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n600), .A2(new_n602), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n636), .A2(new_n633), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n541), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n644), .A2(new_n646), .A3(new_n552), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n548), .B1(new_n549), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n359), .A2(new_n627), .A3(new_n429), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n643), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  INV_X1    g467(.A(new_n308), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n649), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT40), .Z(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n644), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n661));
  INV_X1    g475(.A(new_n374), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n350), .A2(new_n352), .B1(new_n367), .B2(KEYINPUT89), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(new_n371), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n661), .B1(new_n664), .B2(new_n376), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n428), .B1(new_n665), .B2(new_n359), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n637), .A2(new_n666), .A3(new_n552), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n485), .A2(new_n486), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n309), .B1(new_n669), .B2(new_n461), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n456), .A2(new_n463), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n461), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n475), .A2(new_n479), .A3(new_n476), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n479), .B1(new_n475), .B2(new_n476), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT99), .Z(new_n678));
  NAND3_X1  g492(.A1(new_n658), .A2(new_n668), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NAND3_X1  g494(.A1(new_n618), .A2(new_n378), .A3(new_n650), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n643), .A2(new_n647), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  INV_X1    g498(.A(new_n188), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n190), .B1(new_n284), .B2(new_n299), .ZN(new_n686));
  INV_X1    g500(.A(G469), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(G469), .B1(new_n686), .B2(KEYINPUT101), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n490), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT29), .B1(new_n491), .B2(new_n492), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n693), .A2(new_n694), .A3(new_n190), .ZN(new_n695));
  INV_X1    g509(.A(G472), .ZN(new_n696));
  OAI22_X1  g510(.A1(new_n675), .A2(new_n676), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n692), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n644), .A2(new_n552), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n551), .A3(new_n619), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT41), .B(G113), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT102), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n703), .B(new_n705), .ZN(G15));
  AOI21_X1  g520(.A(new_n553), .B1(new_n600), .B2(new_n602), .ZN(new_n707));
  INV_X1    g521(.A(new_n551), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n707), .A2(new_n629), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n686), .A2(new_n687), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n188), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n291), .A2(new_n290), .A3(new_n195), .A4(new_n298), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n195), .B1(new_n303), .B2(new_n291), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n189), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n687), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n711), .B1(new_n689), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n709), .A2(new_n546), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NOR3_X1   g533(.A1(new_n378), .A2(new_n429), .A3(new_n551), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n697), .A2(new_n720), .A3(new_n646), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n717), .A3(new_n707), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  NAND2_X1  g537(.A1(new_n465), .A2(new_n474), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n461), .B1(new_n487), .B2(new_n488), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n476), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n607), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n545), .A2(new_n727), .A3(new_n551), .ZN(new_n728));
  INV_X1    g542(.A(new_n602), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n588), .A2(new_n309), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT86), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n588), .A2(new_n556), .A3(new_n309), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n554), .B1(new_n733), .B2(new_n601), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n666), .B(new_n552), .C1(new_n729), .C2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n717), .A2(new_n728), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR3_X1   g552(.A1(new_n681), .A2(new_n727), .A3(new_n637), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n717), .A2(new_n739), .A3(new_n707), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND3_X1  g555(.A1(new_n600), .A2(new_n552), .A3(new_n602), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n308), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n546), .A3(new_n682), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(new_n546), .A3(KEYINPUT42), .A4(new_n682), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  NAND3_X1  g563(.A1(new_n743), .A2(new_n546), .A3(new_n651), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  AOI21_X1  g565(.A(new_n378), .B1(new_n617), .B2(new_n615), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT43), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n646), .A2(new_n608), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n755), .A2(KEYINPUT103), .A3(KEYINPUT44), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT103), .B1(new_n755), .B2(KEYINPUT44), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n742), .B1(new_n755), .B2(KEYINPUT44), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n302), .A2(new_n304), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT45), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(G469), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n306), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n300), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n188), .A3(new_n656), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT104), .B(G137), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G39));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n188), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n767), .A2(new_n188), .A3(new_n773), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n697), .A2(new_n681), .A3(new_n742), .A4(new_n698), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT106), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NAND2_X1  g596(.A1(new_n775), .A2(new_n776), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n714), .A2(new_n715), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(G469), .A3(new_n689), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n685), .A3(new_n710), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n548), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n753), .A2(new_n545), .A3(new_n788), .A4(new_n727), .ZN(new_n789));
  INV_X1    g603(.A(new_n742), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT114), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n660), .A2(new_n553), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n717), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n799), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n800), .A2(new_n801), .B1(KEYINPUT115), .B2(KEYINPUT50), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n787), .A2(new_n804), .A3(new_n792), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n717), .A2(new_n548), .A3(new_n790), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n753), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT116), .Z(new_n808));
  NOR2_X1   g622(.A1(new_n727), .A2(new_n637), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n806), .A2(new_n678), .A3(new_n545), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n618), .A2(new_n378), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n794), .A2(new_n803), .A3(new_n805), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n803), .A2(KEYINPUT117), .A3(new_n815), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n802), .B2(new_n814), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n787), .B2(new_n792), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n811), .A2(new_n620), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n692), .A2(new_n701), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n547), .B1(new_n789), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n808), .A2(new_n546), .ZN(new_n827));
  XNOR2_X1  g641(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n824), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n818), .A2(new_n823), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n643), .B(new_n647), .C1(new_n651), .C2(new_n682), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n649), .B(KEYINPUT109), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n646), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n736), .A2(new_n654), .A3(new_n677), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n740), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n833), .A2(new_n740), .A3(new_n836), .A4(KEYINPUT52), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n839), .B1(KEYINPUT110), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT110), .B(KEYINPUT111), .Z(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n839), .B(new_n842), .C1(KEYINPUT110), .C2(new_n840), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n603), .A2(new_n620), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT107), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT107), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n603), .A2(new_n850), .A3(new_n620), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n851), .A3(new_n609), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n430), .B(new_n603), .C1(new_n546), .C2(new_n638), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n429), .A2(new_n665), .A3(new_n359), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n609), .A2(new_n603), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n703), .A2(new_n718), .A3(new_n722), .A4(new_n737), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n627), .A2(new_n359), .A3(new_n428), .A4(new_n650), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n742), .A2(new_n860), .A3(new_n637), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n643), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n739), .A2(new_n743), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n750), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT108), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n750), .A2(new_n862), .A3(new_n863), .A4(KEYINPUT108), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n866), .A2(new_n867), .B1(new_n746), .B2(new_n747), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n846), .A2(new_n847), .A3(new_n859), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n839), .A2(new_n840), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n859), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n722), .A2(new_n737), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n785), .A2(new_n697), .A3(new_n698), .A4(new_n688), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n603), .A2(new_n629), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n848), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT112), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n700), .B1(new_n702), .B2(new_n709), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT112), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n722), .A4(new_n737), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n748), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n879), .A2(new_n882), .A3(new_n748), .A4(KEYINPUT113), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n866), .A2(new_n867), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT53), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n846), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n871), .A2(new_n847), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n874), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n832), .A2(new_n896), .B1(G952), .B2(G953), .ZN(new_n897));
  INV_X1    g711(.A(new_n678), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n698), .A2(new_n752), .A3(new_n552), .A4(new_n188), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n660), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n785), .A2(new_n710), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT49), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n897), .B1(new_n900), .B2(new_n902), .ZN(G75));
  AOI21_X1  g717(.A(new_n189), .B1(new_n892), .B2(new_n894), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT56), .B1(new_n904), .B2(new_n555), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n595), .A2(new_n597), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(new_n598), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n909), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n191), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(KEYINPUT119), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n905), .B2(new_n909), .ZN(new_n916));
  AOI211_X1 g730(.A(KEYINPUT56), .B(new_n908), .C1(new_n904), .C2(new_n555), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n914), .A2(new_n918), .ZN(G51));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n189), .B(new_n763), .C1(new_n892), .C2(new_n894), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n306), .B(KEYINPUT57), .Z(new_n922));
  AOI21_X1  g736(.A(new_n890), .B1(new_n885), .B2(new_n886), .ZN(new_n923));
  AOI221_X4 g737(.A(KEYINPUT54), .B1(new_n871), .B2(new_n847), .C1(new_n923), .C2(new_n846), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n712), .A2(new_n713), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n921), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n920), .B1(new_n929), .B2(new_n912), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n858), .A2(KEYINPUT112), .B1(new_n746), .B2(new_n747), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT113), .B1(new_n931), .B2(new_n882), .ZN(new_n932));
  INV_X1    g746(.A(new_n886), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n891), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n844), .A2(new_n845), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n894), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT54), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n895), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n927), .B1(new_n938), .B2(new_n922), .ZN(new_n939));
  OAI211_X1 g753(.A(KEYINPUT120), .B(new_n913), .C1(new_n939), .C2(new_n921), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n930), .A2(new_n940), .ZN(G54));
  NAND4_X1  g755(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .A4(new_n372), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .ZN(new_n945));
  INV_X1    g759(.A(new_n372), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n912), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(G60));
  XOR2_X1   g762(.A(new_n613), .B(KEYINPUT122), .Z(new_n949));
  NAND2_X1  g763(.A1(G478), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT59), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n949), .B1(new_n896), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n938), .A2(new_n949), .A3(new_n951), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n912), .ZN(G63));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n936), .A2(new_n636), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n913), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n961));
  INV_X1    g775(.A(new_n936), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n542), .B1(new_n962), .B2(new_n956), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n960), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(G66));
  INV_X1    g780(.A(G224), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n550), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n859), .B2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n906), .B1(G898), .B2(new_n191), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  AOI21_X1  g785(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n443), .A2(new_n455), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(new_n360), .Z(new_n974));
  NAND2_X1  g788(.A1(G900), .A2(G953), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n769), .B1(new_n779), .B2(new_n780), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n748), .A2(new_n750), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT125), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n833), .A2(new_n740), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT124), .Z(new_n980));
  NOR3_X1   g794(.A1(new_n768), .A2(new_n699), .A3(new_n735), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n976), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n974), .B(new_n975), .C1(new_n983), .C2(G953), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n679), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n980), .A2(KEYINPUT62), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n790), .B1(new_n620), .B2(new_n855), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n657), .A2(new_n988), .A3(new_n699), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT62), .B1(new_n980), .B2(new_n986), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n976), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n974), .B1(new_n992), .B2(new_n191), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n972), .B1(new_n985), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n972), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n992), .A2(new_n191), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n984), .B(new_n995), .C1(new_n996), .C2(new_n974), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n994), .A2(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT126), .Z(new_n1001));
  INV_X1    g815(.A(new_n859), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n992), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n673), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1001), .B1(new_n983), .B2(new_n1002), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n492), .B(KEYINPUT127), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n873), .A2(new_n492), .A3(new_n672), .A4(new_n1000), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n913), .A2(new_n1004), .A3(new_n1007), .A4(new_n1008), .ZN(G57));
endmodule


