//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n189), .A2(KEYINPUT68), .A3(new_n196), .ZN(new_n197));
  OR3_X1    g011(.A1(new_n187), .A2(KEYINPUT68), .A3(new_n188), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G131), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n203), .A2(new_n205), .A3(new_n209), .A4(new_n206), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT65), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT65), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G143), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT65), .A2(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT65), .A2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT66), .A3(G143), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT64), .A2(G143), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT64), .A2(G143), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n218), .A2(new_n222), .A3(new_n223), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n224), .B2(new_n225), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n221), .B2(G143), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n213), .A2(new_n228), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n221), .B2(G143), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n231), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n218), .A2(new_n222), .A3(new_n227), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n204), .A2(G134), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n209), .B1(new_n243), .B2(new_n206), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n203), .A2(new_n206), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n209), .A4(new_n205), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n235), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT30), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n235), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n200), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n235), .A2(new_n250), .A3(new_n200), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G210), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n260), .B(KEYINPUT27), .Z(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT69), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n255), .A2(new_n257), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT31), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n251), .A2(new_n199), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(new_n256), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n256), .A2(new_n268), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n264), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n235), .A2(new_n250), .A3(new_n253), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n253), .B1(new_n235), .B2(new_n250), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n199), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n262), .B(new_n263), .Z(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT71), .B(KEYINPUT31), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n276), .A2(new_n256), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n256), .A3(new_n277), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT31), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n267), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G472), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OR3_X1    g106(.A1(new_n270), .A2(new_n272), .A3(new_n264), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT73), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n255), .A2(new_n257), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(new_n277), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n294), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n295), .A2(KEYINPUT73), .ZN(new_n301));
  OAI21_X1  g115(.A(G472), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n288), .A2(KEYINPUT72), .A3(new_n289), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n286), .A4(new_n287), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n292), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT74), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n306), .A3(G125), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT16), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G125), .B(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT74), .A2(KEYINPUT16), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n229), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n309), .B1(G125), .B2(new_n306), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n320), .A2(KEYINPUT74), .A3(G140), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n307), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n325), .A3(new_n229), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT75), .ZN(new_n327));
  OAI21_X1  g141(.A(G146), .B1(new_n311), .B2(new_n314), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n238), .A2(G119), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n238), .A2(KEYINPUT23), .A3(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n190), .A2(G128), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G110), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n334), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n329), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n312), .B(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n221), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n338), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT76), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n335), .A2(G110), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n328), .B(new_n341), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n339), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n351), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G217), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(G234), .B2(new_n287), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n287), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n359), .B2(KEYINPUT25), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n352), .B2(new_n353), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n358), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n305), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  OAI21_X1  g181(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT79), .Z(new_n369));
  XNOR2_X1  g183(.A(G110), .B(G140), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n259), .A2(G227), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g186(.A(new_n213), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n239), .A2(new_n241), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G104), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT83), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(G104), .B2(new_n375), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT80), .B(G107), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n377), .A2(new_n379), .B1(new_n380), .B2(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n375), .B2(G104), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n380), .A2(new_n384), .B1(new_n386), .B2(new_n376), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT81), .B(G101), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT82), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n376), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n375), .A2(KEYINPUT80), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AND4_X1   g208(.A1(KEYINPUT82), .A2(new_n390), .A3(new_n394), .A4(new_n388), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n382), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n374), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n387), .A2(KEYINPUT82), .A3(new_n388), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n390), .A2(new_n394), .A3(new_n388), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  AND4_X1   g216(.A1(new_n222), .A2(new_n218), .A3(new_n227), .A4(new_n240), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n238), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n216), .A2(new_n217), .B1(new_n226), .B2(G146), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n222), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n402), .B(new_n382), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n373), .B1(new_n397), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT12), .B1(new_n213), .B2(KEYINPUT84), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n408), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n406), .A2(new_n403), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n396), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n390), .A2(new_n394), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(G101), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n389), .B2(new_n395), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n415), .A3(G101), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n418), .A2(new_n228), .A3(new_n234), .A4(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n398), .A2(new_n401), .B1(G101), .B2(new_n381), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT10), .A3(new_n242), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n414), .A2(new_n420), .A3(new_n373), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n372), .B1(new_n411), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n372), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n414), .A2(new_n420), .A3(new_n422), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n213), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT85), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n429), .A3(new_n213), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n425), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n424), .A2(new_n431), .A3(KEYINPUT86), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n408), .A2(new_n410), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n408), .A2(new_n410), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n423), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n372), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n426), .A2(new_n429), .A3(new_n213), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n429), .B1(new_n426), .B2(new_n213), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n423), .B(new_n372), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n433), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n287), .B1(new_n432), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G469), .ZN(new_n444));
  INV_X1    g258(.A(new_n423), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(new_n428), .B2(new_n430), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT88), .B1(new_n446), .B2(new_n372), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n423), .B1(new_n439), .B2(new_n440), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n437), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n411), .A2(new_n423), .A3(new_n372), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT87), .B(G469), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n287), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n369), .B1(new_n444), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n192), .A2(G122), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT98), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n457), .A2(KEYINPUT14), .B1(G116), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(KEYINPUT14), .B2(new_n457), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G107), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(G116), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n380), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n226), .A2(G128), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n238), .A2(G143), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n202), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n202), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n461), .B(new_n464), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(KEYINPUT99), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n472), .B(new_n466), .C1(new_n471), .C2(new_n465), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT99), .B1(new_n465), .B2(new_n471), .ZN(new_n474));
  OAI21_X1  g288(.A(G134), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n463), .A2(new_n380), .ZN(new_n476));
  INV_X1    g290(.A(new_n464), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n467), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n367), .A2(new_n355), .A3(G953), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n470), .B2(new_n478), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n287), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n483), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G113), .B(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(new_n383), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n258), .A2(new_n259), .A3(G143), .A4(G214), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT64), .B(G143), .ZN(new_n491));
  INV_X1    g305(.A(G214), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n492), .A2(G237), .A3(G953), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n490), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G131), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n209), .B(new_n490), .C1(new_n491), .C2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n497), .A2(new_n328), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n340), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n312), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n504), .A3(new_n500), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT94), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n501), .B(new_n506), .C1(new_n500), .C2(new_n312), .ZN(new_n507));
  INV_X1    g321(.A(new_n221), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n498), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n494), .A2(KEYINPUT93), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n209), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT18), .B(G131), .C1(new_n494), .C2(KEYINPUT93), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n340), .A2(new_n221), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n312), .A2(new_n229), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n489), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n495), .A2(new_n518), .A3(new_n496), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n495), .A2(KEYINPUT95), .A3(new_n518), .A4(new_n496), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n494), .A2(KEYINPUT17), .A3(G131), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n489), .B(new_n516), .C1(new_n524), .C2(new_n329), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n328), .B1(new_n326), .B2(KEYINPUT75), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n316), .B1(new_n315), .B2(new_n229), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n530), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n531), .A2(KEYINPUT96), .A3(new_n489), .A4(new_n516), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n517), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(G475), .A2(G902), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT20), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT97), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(KEYINPUT20), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  OR3_X1    g352(.A1(new_n533), .A2(KEYINPUT20), .A3(new_n534), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n489), .B1(new_n531), .B2(new_n516), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n527), .B2(new_n532), .ZN(new_n542));
  OAI21_X1  g356(.A(G475), .B1(new_n542), .B2(G902), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n487), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n259), .A2(G952), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(G234), .B2(G237), .ZN(new_n546));
  NAND2_X1  g360(.A1(G234), .A2(G237), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(G902), .A3(G953), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT21), .B(G898), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G214), .B1(G237), .B2(G902), .ZN(new_n553));
  OAI21_X1  g367(.A(G210), .B1(G237), .B2(G902), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT90), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n418), .A2(new_n199), .A3(new_n419), .ZN(new_n557));
  OAI21_X1  g371(.A(G113), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(KEYINPUT5), .B2(new_n188), .ZN(new_n559));
  INV_X1    g373(.A(new_n189), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n421), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT89), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT89), .B1(new_n557), .B2(new_n562), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT6), .B(new_n556), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n556), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n557), .A2(new_n562), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT89), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT89), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n557), .A2(new_n562), .A3(new_n555), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT6), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n565), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n228), .A2(G125), .A3(new_n234), .ZN(new_n576));
  AOI21_X1  g390(.A(G125), .B1(new_n239), .B2(new_n241), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n259), .A2(G224), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n578), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT91), .B(KEYINPUT8), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n555), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n558), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n558), .A2(new_n586), .B1(new_n188), .B2(KEYINPUT5), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n560), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n421), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n421), .A2(new_n561), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n578), .B1(new_n593), .B2(new_n580), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT7), .B(new_n579), .C1(new_n576), .C2(new_n577), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n592), .A2(new_n594), .A3(new_n572), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n287), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n554), .B1(new_n582), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n554), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n600), .B(new_n597), .C1(new_n575), .C2(new_n581), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n553), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n455), .A2(new_n552), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n366), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n388), .B(KEYINPUT100), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G3));
  INV_X1    g421(.A(new_n288), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n364), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n455), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n540), .A2(new_n543), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n483), .A2(G478), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n470), .A2(new_n478), .ZN(new_n614));
  INV_X1    g428(.A(new_n479), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n480), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT33), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n619), .A3(new_n480), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n287), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n613), .B1(new_n622), .B2(G478), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n612), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n581), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n556), .B1(new_n563), .B2(new_n564), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n573), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n627), .B2(new_n565), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n600), .B1(new_n628), .B2(new_n597), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n582), .A2(new_n554), .A3(new_n598), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n551), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n553), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n611), .A2(new_n624), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND3_X1  g450(.A1(new_n540), .A2(new_n543), .A3(new_n486), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n611), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT35), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NAND2_X1  g454(.A1(new_n359), .A2(KEYINPUT25), .ZN(new_n641));
  INV_X1    g455(.A(new_n356), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n361), .B2(new_n362), .ZN(new_n643));
  INV_X1    g457(.A(new_n351), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n348), .B(new_n645), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n641), .A2(new_n643), .B1(new_n646), .B2(new_n357), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n608), .A2(new_n647), .A3(new_n609), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n455), .A2(new_n648), .A3(new_n552), .A4(new_n603), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  INV_X1    g465(.A(new_n369), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n452), .A2(new_n287), .A3(new_n453), .ZN(new_n653));
  INV_X1    g467(.A(G469), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT86), .B1(new_n424), .B2(new_n431), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n438), .A2(new_n441), .A3(new_n433), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n657), .B2(new_n287), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n652), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n546), .B(KEYINPUT102), .ZN(new_n660));
  NOR2_X1   g474(.A1(KEYINPUT101), .A2(G900), .ZN(new_n661));
  AND2_X1   g475(.A1(KEYINPUT101), .A2(G900), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n549), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n540), .A2(new_n543), .A3(new_n486), .A4(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n602), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n647), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT103), .B1(new_n665), .B2(new_n602), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n667), .A2(new_n305), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XNOR2_X1  g485(.A(new_n664), .B(KEYINPUT39), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n455), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n269), .A2(new_n256), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n265), .B1(new_n675), .B2(new_n264), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n676), .B2(G902), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n292), .A2(new_n303), .A3(new_n304), .A4(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n612), .A2(new_n486), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n631), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n553), .A3(new_n647), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n674), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n491), .B(KEYINPUT105), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G45));
  AOI211_X1 g501(.A(new_n602), .B(new_n369), .C1(new_n444), .C2(new_n454), .ZN(new_n688));
  INV_X1    g502(.A(new_n613), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n618), .B2(new_n620), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(new_n484), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n543), .B2(new_n540), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n664), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n688), .A2(new_n305), .A3(new_n668), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  NAND2_X1  g510(.A1(new_n452), .A2(new_n287), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G469), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n698), .A2(new_n652), .A3(new_n454), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n624), .A2(new_n633), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n305), .A2(new_n699), .A3(new_n365), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT106), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NOR2_X1   g518(.A1(new_n633), .A2(new_n637), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n305), .A2(new_n699), .A3(new_n365), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND4_X1  g521(.A1(new_n698), .A2(new_n603), .A3(new_n652), .A4(new_n454), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n305), .A3(new_n552), .A4(new_n668), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NOR2_X1   g525(.A1(new_n680), .A2(new_n602), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n282), .A2(KEYINPUT31), .ZN(new_n713));
  AOI211_X1 g527(.A(G472), .B(G902), .C1(new_n281), .C2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT107), .B(G472), .Z(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n285), .B2(new_n287), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n364), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n699), .A2(new_n632), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NOR2_X1   g533(.A1(new_n716), .A2(new_n714), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n668), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n708), .A2(new_n693), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n320), .ZN(G27));
  NOR2_X1   g537(.A1(new_n424), .A2(new_n431), .ZN(new_n724));
  OAI21_X1  g538(.A(G469), .B1(new_n724), .B2(G902), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n454), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n629), .A2(new_n630), .A3(new_n553), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n369), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n305), .A2(new_n729), .A3(new_n365), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n290), .A2(KEYINPUT108), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n288), .A2(new_n733), .A3(new_n289), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n302), .A3(new_n304), .A4(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n729), .A3(new_n694), .A4(new_n365), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n730), .A2(new_n731), .B1(new_n736), .B2(KEYINPUT42), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n665), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n730), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n305), .A3(new_n729), .A4(new_n365), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT110), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n612), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT43), .A3(new_n623), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n612), .B2(new_n691), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n668), .B1(new_n608), .B2(new_n609), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT112), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(new_n754), .A3(KEYINPUT44), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n657), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n654), .B1(new_n724), .B2(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n654), .A2(new_n287), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n454), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT46), .B1(new_n762), .B2(new_n764), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n652), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n672), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n727), .B(KEYINPUT113), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n757), .A2(new_n758), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  NOR4_X1   g587(.A1(new_n305), .A2(new_n365), .A3(new_n693), .A4(new_n727), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n768), .A2(KEYINPUT114), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n652), .C1(new_n766), .C2(new_n767), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n779), .A3(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n776), .A2(new_n778), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n775), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n306), .ZN(G42));
  NAND2_X1  g600(.A1(new_n748), .A2(new_n623), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n652), .A2(new_n553), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n787), .A2(new_n682), .A3(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n698), .A2(new_n454), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT49), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n789), .A2(new_n791), .A3(new_n365), .A4(new_n679), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n790), .A2(new_n546), .A3(new_n728), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n612), .A2(new_n623), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n365), .A3(new_n679), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT119), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n728), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n660), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT116), .B1(new_n752), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n801), .B(new_n660), .C1(new_n749), .C2(new_n751), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n798), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n796), .B1(new_n721), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n682), .A2(new_n553), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n699), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n717), .B(new_n806), .C1(new_n800), .C2(new_n802), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT50), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT50), .ZN(new_n811));
  INV_X1    g625(.A(new_n770), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n717), .B(new_n812), .C1(new_n800), .C2(new_n802), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n782), .A2(new_n784), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n790), .A2(new_n369), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT117), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n810), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  INV_X1    g634(.A(new_n811), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n804), .A3(new_n809), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n782), .A2(new_n784), .A3(new_n816), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n823), .B2(new_n814), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n819), .A2(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n693), .A2(new_n721), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n709), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n647), .A2(new_n652), .A3(new_n664), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n678), .A2(new_n712), .A3(new_n726), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n670), .A2(new_n695), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n288), .A2(KEYINPUT72), .A3(new_n289), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT72), .B1(new_n288), .B2(new_n289), .ZN(new_n836));
  INV_X1    g650(.A(new_n304), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n647), .B1(new_n838), .B2(new_n302), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n659), .A2(new_n693), .A3(new_n602), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n722), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n670), .A4(new_n831), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n701), .A2(new_n710), .A3(new_n718), .A4(new_n706), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n455), .B(new_n610), .C1(new_n700), .C2(new_n705), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n845), .B(new_n649), .C1(new_n366), .C2(new_n604), .ZN(new_n846));
  INV_X1    g660(.A(new_n664), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n544), .A2(new_n847), .A3(new_n727), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n305), .A2(new_n848), .A3(new_n455), .A4(new_n668), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n827), .A2(new_n729), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n745), .A2(new_n844), .A3(new_n852), .A4(new_n737), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n826), .B1(new_n843), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n745), .A2(new_n852), .A3(new_n737), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n834), .A2(new_n842), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT53), .A4(new_n844), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n858), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n709), .B(new_n717), .C1(new_n800), .C2(new_n802), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n793), .A2(new_n365), .A3(new_n679), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n545), .B1(new_n863), .B2(new_n692), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n735), .A2(new_n365), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n867), .B(new_n798), .C1(new_n800), .C2(new_n802), .ZN(new_n868));
  XNOR2_X1  g682(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n871), .A3(new_n864), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n869), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n866), .A2(new_n870), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT122), .ZN(new_n875));
  INV_X1    g689(.A(new_n869), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n868), .B(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n872), .A4(new_n866), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n825), .A2(new_n859), .A3(new_n861), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n792), .B1(new_n881), .B2(new_n882), .ZN(G75));
  AOI21_X1  g697(.A(new_n287), .B1(new_n854), .B2(new_n858), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(G210), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n575), .B(new_n625), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n885), .B2(new_n886), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n259), .A2(G952), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G51));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n859), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n854), .A2(new_n858), .A3(KEYINPUT123), .A4(new_n855), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n861), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n763), .B(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n452), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n884), .A2(new_n760), .A3(new_n761), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n891), .B1(new_n899), .B2(new_n900), .ZN(G54));
  INV_X1    g715(.A(new_n884), .ZN(new_n902));
  NAND2_X1  g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n533), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n891), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n902), .A2(new_n533), .A3(new_n903), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(G60));
  XOR2_X1   g722(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n909));
  NOR2_X1   g723(.A1(new_n484), .A2(new_n287), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n861), .B2(new_n859), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n905), .B1(new_n912), .B2(new_n621), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n618), .B2(new_n620), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n896), .B2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n860), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n352), .A3(new_n353), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n860), .A2(new_n646), .A3(new_n917), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n905), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(KEYINPUT61), .A3(new_n905), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G66));
  INV_X1    g739(.A(new_n846), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n844), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(G224), .A2(G953), .ZN(new_n928));
  OAI22_X1  g742(.A1(new_n927), .A2(G953), .B1(new_n550), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n627), .B(new_n565), .C1(G898), .C2(new_n259), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n929), .B(new_n930), .Z(G69));
  AOI21_X1  g745(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT126), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n252), .A2(new_n254), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n507), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n841), .A2(new_n670), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n685), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n685), .A3(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n815), .A2(new_n774), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n624), .A2(new_n637), .ZN(new_n944));
  NOR4_X1   g758(.A1(new_n366), .A2(new_n673), .A3(new_n727), .A4(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n942), .A2(new_n772), .A3(new_n943), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n936), .B1(new_n947), .B2(new_n259), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n935), .B1(G900), .B2(G953), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n867), .A2(new_n712), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n951), .A2(new_n769), .A3(new_n768), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n736), .A2(KEYINPUT42), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n730), .A2(new_n731), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(new_n745), .A3(new_n772), .A4(new_n937), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n785), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n950), .B1(new_n957), .B2(new_n259), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n933), .B1(new_n948), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n932), .A2(KEYINPUT126), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G72));
  INV_X1    g775(.A(new_n860), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n298), .B2(new_n265), .ZN(new_n965));
  INV_X1    g779(.A(new_n964), .ZN(new_n966));
  INV_X1    g780(.A(new_n927), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n957), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n297), .A2(new_n264), .ZN(new_n969));
  OAI221_X1 g783(.A(new_n905), .B1(new_n962), .B2(new_n965), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n964), .B1(new_n947), .B2(new_n927), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n264), .B(new_n297), .C1(new_n971), .C2(KEYINPUT127), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G57));
endmodule


