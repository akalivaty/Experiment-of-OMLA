//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n188));
  INV_X1    g002(.A(G210), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(G237), .A3(G953), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT26), .B(G101), .Z(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  AOI21_X1  g010(.A(G131), .B1(new_n195), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n197), .A3(new_n202), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(G128), .B(new_n206), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n211), .B(new_n212), .C1(KEYINPUT1), .C2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n195), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n198), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n204), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT65), .A2(G116), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT65), .A2(G116), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G119), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT2), .B(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n227), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n222), .A3(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n219), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n196), .B(new_n199), .C1(G134), .C2(new_n198), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n204), .A2(KEYINPUT66), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT66), .B1(new_n204), .B2(new_n235), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n211), .A2(new_n212), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G143), .B(G146), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G128), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n233), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n201), .A2(new_n203), .B1(G131), .B2(new_n234), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n219), .B1(new_n246), .B2(new_n243), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n247), .A2(new_n231), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT28), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n204), .A2(new_n235), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n244), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n210), .A2(new_n218), .A3(new_n214), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n203), .B2(new_n201), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(new_n231), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT28), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n193), .B1(new_n249), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(KEYINPUT30), .A3(new_n219), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n232), .B1(new_n247), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n254), .A2(new_n257), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n264), .A2(new_n193), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n187), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT70), .B(new_n187), .C1(new_n260), .C2(new_n266), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n232), .B1(new_n254), .B2(new_n219), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(KEYINPUT28), .C1(new_n272), .C2(new_n245), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n254), .A2(new_n219), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n231), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n276), .B2(new_n265), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n193), .A2(new_n187), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n270), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G472), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n247), .A2(new_n231), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n274), .B1(new_n265), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n193), .B1(new_n285), .B2(new_n258), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n193), .B1(new_n254), .B2(new_n257), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n219), .A2(KEYINPUT30), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n238), .B2(new_n244), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n243), .B1(new_n204), .B2(new_n235), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n262), .B1(new_n290), .B2(new_n256), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n231), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n287), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT31), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n264), .A2(new_n295), .A3(new_n287), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n298), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n297), .A2(KEYINPUT68), .A3(new_n298), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT69), .B(KEYINPUT32), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n283), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT9), .B(G234), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT74), .ZN(new_n308));
  OAI21_X1  g122(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G140), .ZN(new_n310));
  INV_X1    g124(.A(G953), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G227), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n310), .B(new_n312), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(KEYINPUT75), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g132(.A(G104), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n316), .A2(new_n318), .B1(new_n319), .B2(G107), .ZN(new_n320));
  INV_X1    g134(.A(G107), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G104), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n319), .A2(G107), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G101), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G101), .B1(new_n323), .B2(new_n322), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n210), .A2(new_n214), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT10), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT10), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n327), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n323), .A2(new_n324), .ZN(new_n336));
  INV_X1    g150(.A(new_n322), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n323), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G101), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT4), .A3(new_n327), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n326), .B1(new_n320), .B2(new_n325), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n243), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n314), .B1(new_n346), .B2(new_n238), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n331), .A2(new_n334), .B1(new_n341), .B2(new_n344), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n252), .A2(new_n253), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n313), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT77), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n327), .A2(new_n329), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n210), .A2(new_n214), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n354), .A2(new_n355), .B1(new_n332), .B2(new_n327), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n250), .A2(KEYINPUT12), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n357), .A2(KEYINPUT12), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n346), .A2(new_n238), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n350), .A2(new_n351), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n313), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI211_X1 g177(.A(G469), .B(G902), .C1(new_n360), .C2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n356), .A2(new_n358), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n327), .A2(new_n329), .ZN(new_n366));
  OAI22_X1  g180(.A1(new_n366), .A2(new_n215), .B1(new_n328), .B2(new_n330), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n252), .A3(new_n253), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT12), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n313), .B1(new_n370), .B2(new_n361), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n352), .A2(KEYINPUT76), .ZN(new_n372));
  OAI211_X1 g186(.A(KEYINPUT76), .B(new_n314), .C1(new_n346), .C2(new_n238), .ZN(new_n373));
  INV_X1    g187(.A(new_n362), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n371), .B(G469), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(G469), .A2(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n309), .B1(new_n364), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n309), .C1(new_n364), .C2(new_n378), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n222), .A2(KEYINPUT5), .A3(new_n225), .ZN(new_n385));
  INV_X1    g199(.A(G113), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT5), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n386), .B1(new_n224), .B2(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n385), .A2(KEYINPUT80), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT80), .B1(new_n385), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n327), .A2(new_n230), .A3(new_n329), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n342), .A2(new_n343), .B1(new_n228), .B2(new_n230), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n391), .A2(new_n392), .B1(new_n393), .B2(new_n341), .ZN(new_n394));
  XNOR2_X1  g208(.A(G110), .B(G122), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n384), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n395), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n392), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(new_n341), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n400), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n396), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n394), .A2(new_n398), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n384), .A4(new_n397), .ZN(new_n407));
  INV_X1    g221(.A(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n355), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n243), .A2(new_n410), .A3(G125), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n243), .A2(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT82), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n311), .A2(G224), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n415), .B(new_n416), .Z(new_n417));
  NAND3_X1  g231(.A1(new_n403), .A2(new_n407), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n385), .A2(new_n388), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n385), .A2(KEYINPUT80), .A3(new_n388), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n230), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n354), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n392), .A2(new_n419), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n395), .B(KEYINPUT8), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n416), .A2(KEYINPUT7), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n412), .A2(KEYINPUT83), .A3(new_n414), .A4(new_n431), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n431), .A2(KEYINPUT83), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n414), .A2(new_n409), .A3(new_n411), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(KEYINPUT83), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n437), .A3(KEYINPUT84), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n427), .B1(new_n424), .B2(new_n425), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n432), .A2(new_n436), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n394), .A2(new_n395), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G902), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n418), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n418), .A2(new_n444), .A3(new_n445), .A4(new_n447), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n452), .B(KEYINPUT79), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G475), .ZN(new_n456));
  INV_X1    g270(.A(G237), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n311), .A3(G214), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n205), .ZN(new_n459));
  INV_X1    g273(.A(G131), .ZN(new_n460));
  NOR2_X1   g274(.A1(G237), .A2(G953), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(G143), .A3(G214), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT17), .ZN(new_n465));
  INV_X1    g279(.A(new_n462), .ZN(new_n466));
  AOI21_X1  g280(.A(G143), .B1(new_n461), .B2(G214), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n459), .A2(new_n469), .A3(new_n460), .A4(new_n462), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n464), .A2(new_n465), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n408), .A2(KEYINPUT16), .A3(G140), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT72), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G140), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G125), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n408), .A2(G140), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT16), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n473), .B1(new_n479), .B2(new_n472), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n208), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n479), .A2(new_n472), .ZN(new_n482));
  OAI211_X1 g296(.A(G146), .B(new_n474), .C1(new_n482), .C2(new_n473), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n459), .A2(new_n462), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT17), .A3(G131), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n471), .A2(new_n481), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G125), .B(G140), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n487), .A2(new_n208), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n208), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT18), .A2(G131), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n488), .A2(new_n489), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n459), .A2(new_n462), .A3(new_n490), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n484), .A2(KEYINPUT85), .A3(new_n491), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G113), .B(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n319), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT88), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n486), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n486), .A2(new_n496), .A3(new_n502), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n486), .A2(new_n496), .ZN(new_n505));
  INV_X1    g319(.A(new_n498), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n456), .B1(new_n508), .B2(new_n445), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n487), .B(KEYINPUT19), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n208), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n464), .A2(new_n468), .A3(new_n470), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(KEYINPUT87), .A3(new_n208), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n483), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n498), .B1(new_n516), .B2(new_n496), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT90), .B1(new_n504), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n501), .B2(new_n503), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI22_X1  g336(.A1(new_n519), .A2(KEYINPUT20), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n504), .A2(new_n518), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(KEYINPUT90), .A3(new_n525), .A4(new_n521), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n509), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n445), .B(new_n311), .C1(G234), .C2(G237), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT21), .B(G898), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G952), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(G953), .ZN(new_n532));
  INV_X1    g346(.A(G234), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(new_n457), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n311), .A2(G217), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n308), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n213), .A2(G143), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n205), .A2(G128), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(G134), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n539), .A2(new_n541), .A3(new_n195), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n220), .A2(G122), .A3(new_n221), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n223), .A2(G122), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n321), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT14), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n546), .A2(new_n549), .A3(new_n547), .ZN(new_n550));
  OAI21_X1  g364(.A(G107), .B1(new_n546), .B2(new_n549), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n545), .B(new_n548), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n540), .A2(new_n542), .ZN(new_n553));
  OAI21_X1  g367(.A(G134), .B1(new_n541), .B2(KEYINPUT13), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n554), .A2(new_n539), .A3(new_n541), .ZN(new_n556));
  INV_X1    g370(.A(new_n548), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n321), .B1(new_n546), .B2(new_n547), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n538), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(new_n559), .A3(new_n538), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n536), .B1(new_n563), .B2(new_n445), .ZN(new_n564));
  INV_X1    g378(.A(new_n562), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n536), .B(new_n445), .C1(new_n565), .C2(new_n560), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n564), .A2(new_n567), .B1(KEYINPUT15), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT15), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n566), .A2(new_n570), .A3(G478), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n527), .A2(new_n535), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n455), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G217), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(G234), .B2(new_n445), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  INV_X1    g394(.A(G119), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(G128), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(new_n583), .C1(G119), .C2(new_n213), .ZN(new_n584));
  XNOR2_X1  g398(.A(G119), .B(G128), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT24), .B(G110), .Z(new_n586));
  OAI22_X1  g400(.A1(new_n584), .A2(G110), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n483), .A2(new_n587), .A3(new_n489), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(G110), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n585), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n483), .B2(new_n481), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT22), .B(G137), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n311), .A2(G221), .A3(G234), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(KEYINPUT73), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n588), .B2(new_n592), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n579), .B1(new_n600), .B2(G902), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n597), .A2(KEYINPUT25), .A3(new_n445), .A4(new_n599), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n578), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n600), .A2(G902), .A3(new_n577), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n306), .A2(new_n383), .A3(new_n575), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT92), .B(G101), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  NAND3_X1  g422(.A1(new_n563), .A2(new_n568), .A3(new_n445), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n568), .A2(new_n445), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n560), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n563), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n609), .B(new_n611), .C1(new_n615), .C2(new_n568), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n523), .A2(new_n526), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n508), .A2(new_n445), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G475), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n453), .B1(new_n449), .B2(new_n450), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n620), .A2(new_n621), .A3(new_n535), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n302), .A2(new_n303), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n297), .A2(new_n445), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(G472), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT93), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(KEYINPUT93), .A3(G472), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n622), .A2(new_n383), .A3(new_n629), .A4(new_n605), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  AND2_X1   g446(.A1(new_n621), .A2(new_n535), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n383), .A2(new_n629), .A3(new_n633), .A4(new_n605), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n520), .A2(new_n522), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n525), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n520), .A2(KEYINPUT20), .A3(new_n522), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n572), .B(new_n619), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT35), .B(G107), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NAND2_X1  g455(.A1(new_n601), .A2(new_n602), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n577), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n593), .B(new_n644), .Z(new_n645));
  NOR2_X1   g459(.A1(new_n577), .A2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n383), .A2(new_n575), .A3(new_n629), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  AND3_X1   g465(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n298), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n297), .A2(KEYINPUT68), .A3(new_n298), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT68), .B1(new_n297), .B2(new_n298), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n652), .B1(new_n655), .B2(new_n304), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n656), .A2(new_n283), .B1(new_n382), .B2(new_n380), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n451), .A2(new_n454), .A3(new_n648), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n528), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n534), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n658), .A2(new_n638), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XNOR2_X1  g479(.A(new_n661), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n383), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT97), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n667), .B(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n276), .A2(new_n193), .A3(new_n265), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n445), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n193), .B1(new_n264), .B2(new_n265), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n305), .A2(new_n299), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT95), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n305), .A2(KEYINPUT95), .A3(new_n299), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT96), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n451), .B(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n527), .A2(new_n648), .A3(new_n573), .A4(new_n453), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n674), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n205), .ZN(G45));
  INV_X1    g506(.A(KEYINPUT90), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n524), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n635), .B1(new_n694), .B2(new_n525), .ZN(new_n695));
  INV_X1    g509(.A(new_n526), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n619), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n616), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n661), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n658), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n306), .A3(new_n383), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT98), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n657), .A2(KEYINPUT98), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(G469), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT12), .B1(new_n238), .B2(new_n367), .ZN(new_n708));
  OAI22_X1  g522(.A1(new_n352), .A2(KEYINPUT77), .B1(new_n708), .B2(new_n365), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n347), .A2(new_n348), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n363), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n707), .B1(new_n711), .B2(new_n445), .ZN(new_n712));
  INV_X1    g526(.A(new_n309), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n364), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n306), .A2(new_n622), .A3(new_n605), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  INV_X1    g531(.A(new_n638), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n621), .A2(new_n718), .A3(new_n535), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n306), .A2(new_n719), .A3(new_n605), .A4(new_n714), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND2_X1  g535(.A1(new_n714), .A2(new_n621), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n648), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n574), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n306), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  INV_X1    g541(.A(new_n604), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n643), .A2(KEYINPUT99), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n603), .B2(new_n604), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n193), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n294), .A3(new_n296), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n298), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n625), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n527), .A2(new_n573), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n633), .A3(new_n738), .A4(new_n714), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  NAND3_X1  g554(.A1(new_n735), .A2(new_n625), .A3(new_n648), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n722), .A2(new_n699), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n408), .ZN(G27));
  NAND4_X1  g557(.A1(new_n449), .A2(new_n309), .A3(new_n454), .A4(new_n450), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT100), .B1(new_n375), .B2(new_n372), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT76), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n347), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT100), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n374), .A4(new_n373), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT101), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n751), .A3(G469), .A4(new_n371), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n711), .A2(new_n707), .A3(new_n445), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n752), .A2(new_n753), .A3(new_n377), .ZN(new_n754));
  INV_X1    g568(.A(new_n371), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n745), .B2(new_n749), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n751), .B1(new_n756), .B2(G469), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n744), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n699), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n306), .A3(new_n605), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT32), .B1(new_n297), .B2(new_n298), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT103), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n652), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT32), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n300), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT103), .B1(new_n767), .B2(new_n299), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n732), .B1(new_n769), .B2(new_n283), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n752), .A2(new_n753), .A3(new_n377), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n757), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n697), .A2(new_n698), .A3(KEYINPUT42), .A4(new_n661), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n744), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n761), .A2(new_n762), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n460), .ZN(G33));
  NOR2_X1   g590(.A1(new_n638), .A2(new_n662), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n759), .A2(new_n306), .A3(new_n605), .A4(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT104), .B(G134), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G36));
  NOR2_X1   g594(.A1(new_n629), .A2(new_n724), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT107), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n527), .B(KEYINPUT106), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT43), .A3(new_n698), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n697), .A2(new_n616), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(KEYINPUT43), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n782), .A2(KEYINPUT44), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT108), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n782), .A2(new_n789), .A3(KEYINPUT44), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT44), .B1(new_n782), .B2(new_n786), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n449), .A2(new_n454), .A3(new_n450), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n756), .A2(KEYINPUT45), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n375), .A2(new_n372), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n755), .ZN(new_n796));
  OAI21_X1  g610(.A(G469), .B1(new_n796), .B2(KEYINPUT45), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT105), .A3(KEYINPUT46), .A4(new_n377), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT105), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n377), .B1(new_n794), .B2(new_n797), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n364), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n309), .A3(new_n666), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n792), .A2(new_n793), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n791), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  NAND2_X1  g623(.A1(new_n805), .A2(new_n309), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT47), .ZN(new_n811));
  OR4_X1    g625(.A1(new_n306), .A2(new_n605), .A3(new_n699), .A4(new_n793), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n476), .ZN(G42));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n742), .B1(new_n657), .B2(new_n663), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n738), .A2(new_n621), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n724), .A2(new_n309), .A3(new_n661), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n772), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n683), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT98), .B1(new_n657), .B2(new_n700), .ZN(new_n822));
  AND4_X1   g636(.A1(KEYINPUT98), .A2(new_n700), .A3(new_n306), .A4(new_n383), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n817), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n705), .A2(new_n827), .A3(new_n817), .A4(new_n821), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n715), .A2(new_n720), .A3(new_n726), .A4(new_n739), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n775), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT109), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n606), .B2(new_n630), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n527), .A2(new_n572), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n649), .B1(new_n634), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n606), .A2(new_n630), .A3(new_n832), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n648), .A2(new_n573), .A3(new_n661), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n619), .B1(new_n636), .B2(new_n637), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n838), .A2(new_n793), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n657), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n741), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n759), .A2(new_n760), .A3(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n841), .A2(new_n778), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n831), .A2(new_n836), .A3(new_n837), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n816), .B1(new_n829), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n824), .A2(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n828), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n845), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n846), .A2(KEYINPUT111), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n853), .B(new_n816), .C1(new_n829), .C2(new_n845), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n815), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n850), .B1(new_n848), .B2(new_n845), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n836), .A2(new_n837), .A3(new_n844), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n775), .A2(new_n830), .A3(new_n816), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n828), .A3(new_n826), .A4(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n856), .A2(new_n815), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT113), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n846), .A2(KEYINPUT111), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n849), .A2(new_n851), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n854), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n856), .A2(new_n859), .A3(new_n815), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n687), .A2(new_n453), .A3(new_n714), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n869), .B(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n732), .A2(new_n736), .A3(new_n534), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n786), .A2(new_n873), .ZN(new_n874));
  OR3_X1    g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n872), .B1(new_n871), .B2(new_n874), .ZN(new_n876));
  INV_X1    g690(.A(new_n712), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n753), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n878), .A2(new_n793), .A3(new_n713), .A4(new_n534), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n786), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n875), .A2(new_n876), .B1(new_n842), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n309), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n882), .B2(new_n878), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n811), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n793), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n786), .A2(new_n886), .A3(new_n873), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT114), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n683), .B(KEYINPUT96), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n879), .A2(new_n605), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n527), .A3(new_n616), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n881), .B(new_n889), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n894), .A2(new_n895), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(KEYINPUT51), .A3(new_n889), .A4(new_n881), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n880), .A2(new_n770), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT48), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n874), .A2(new_n722), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT118), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n890), .A2(new_n620), .A3(new_n891), .ZN(new_n905));
  AND4_X1   g719(.A1(new_n532), .A2(new_n902), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n898), .A2(new_n900), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n861), .A2(new_n868), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n531), .A2(new_n311), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n732), .A2(new_n713), .A3(new_n453), .A4(new_n616), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n878), .A2(KEYINPUT49), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n878), .A2(KEYINPUT49), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n890), .A2(new_n687), .A3(new_n783), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n910), .A2(new_n915), .ZN(G75));
  AND2_X1   g730(.A1(new_n403), .A2(new_n407), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n417), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n856), .A2(new_n859), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n445), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G210), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g740(.A(KEYINPUT56), .B(new_n919), .C1(new_n923), .C2(G210), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n311), .A2(G952), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G51));
  INV_X1    g743(.A(new_n798), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n921), .A2(G902), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n921), .A2(new_n933), .A3(G902), .A4(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n711), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n867), .A2(KEYINPUT119), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n921), .A2(KEYINPUT54), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n856), .A2(new_n859), .A3(new_n939), .A4(new_n815), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n377), .B(KEYINPUT57), .Z(new_n942));
  AOI21_X1  g756(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n942), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n815), .B1(new_n856), .B2(new_n859), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n860), .B2(new_n939), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(new_n937), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT120), .B1(new_n949), .B2(new_n936), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n928), .B1(new_n945), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n520), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n520), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n928), .ZN(G60));
  XOR2_X1   g769(.A(new_n610), .B(KEYINPUT59), .Z(new_n956));
  NAND3_X1  g770(.A1(new_n941), .A2(new_n615), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n928), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n855), .A2(KEYINPUT113), .A3(new_n860), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n962), .B2(new_n614), .ZN(G63));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT60), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(KEYINPUT60), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n921), .A2(new_n645), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(new_n958), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n600), .B1(new_n922), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT61), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  AOI211_X1 g788(.A(KEYINPUT122), .B(new_n974), .C1(new_n968), .C2(new_n970), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n973), .A2(new_n975), .ZN(G66));
  INV_X1    g790(.A(G224), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n529), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT123), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n836), .A2(new_n837), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n830), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n982), .B2(new_n311), .ZN(new_n983));
  INV_X1    g797(.A(G898), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n917), .B1(new_n984), .B2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  AOI21_X1  g800(.A(new_n813), .B1(new_n791), .B2(new_n807), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n705), .A2(new_n817), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT62), .B1(new_n691), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n697), .A2(new_n698), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n793), .B1(new_n990), .B2(new_n834), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n671), .A2(new_n306), .A3(new_n605), .A4(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n993));
  INV_X1    g807(.A(new_n988), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n993), .B(new_n994), .C1(new_n674), .C2(new_n690), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n987), .A2(new_n989), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n311), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n261), .A2(new_n291), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n510), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT124), .Z(new_n1000));
  NAND3_X1  g814(.A1(new_n770), .A2(new_n621), .A3(new_n738), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n806), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n778), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n1002), .A2(new_n988), .A3(new_n775), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n987), .A2(new_n311), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n999), .B1(G900), .B2(G953), .ZN(new_n1006));
  AOI22_X1  g820(.A1(new_n997), .A2(new_n1000), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n311), .B1(G227), .B2(G900), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(KEYINPUT125), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1007), .B(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n996), .B2(new_n982), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n677), .ZN(new_n1015));
  INV_X1    g829(.A(new_n266), .ZN(new_n1016));
  INV_X1    g830(.A(new_n677), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n1017), .A3(new_n1013), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT126), .Z(new_n1019));
  NAND2_X1  g833(.A1(new_n864), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n987), .A2(new_n981), .A3(new_n1004), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n1013), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n928), .B1(new_n1022), .B2(new_n266), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1015), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(KEYINPUT127), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1015), .A2(new_n1023), .A3(new_n1026), .A4(new_n1020), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1025), .A2(new_n1027), .ZN(G57));
endmodule


