//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994;
  AND2_X1   g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n208), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n213), .A3(KEYINPUT71), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(new_n204), .C1(new_n207), .C2(new_n208), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G226gat), .A2(G233gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G169gat), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT23), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n221), .B1(new_n229), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n232), .A2(new_n238), .A3(new_n235), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n232), .B2(new_n235), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n230), .A2(new_n231), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n221), .B1(new_n242), .B2(new_n233), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n227), .B(new_n228), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n222), .A2(new_n245), .A3(new_n223), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n237), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n235), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n242), .B2(KEYINPUT26), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n242), .A2(KEYINPUT68), .A3(KEYINPUT26), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  NOR2_X1   g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n251), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT27), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G183gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n260), .A3(new_n226), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n261), .A2(new_n262), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n257), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n220), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n219), .B1(new_n249), .B2(new_n265), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n218), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n220), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT29), .B1(new_n249), .B2(new_n265), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n271), .B(new_n217), .C1(new_n220), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT72), .ZN(new_n276));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT73), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n281), .B(new_n278), .C1(new_n270), .C2(new_n273), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n278), .B1(new_n270), .B2(new_n273), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT30), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n274), .B2(new_n279), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT83), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n279), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n281), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(KEYINPUT73), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n283), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT83), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n274), .A2(new_n279), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(KEYINPUT30), .B2(new_n286), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G1gat), .B(G29gat), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT0), .ZN(new_n299));
  XNOR2_X1  g098(.A(G57gat), .B(G85gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303));
  AND2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(G155gat), .B2(G162gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G141gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(G148gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G141gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G155gat), .B(G162gat), .ZN(new_n316));
  INV_X1    g115(.A(G155gat), .ZN(new_n317));
  INV_X1    g116(.A(G162gat), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT2), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n329), .B(new_n330), .C1(new_n331), .C2(KEYINPUT69), .ZN(new_n332));
  INV_X1    g131(.A(G127gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G134gat), .ZN(new_n334));
  INV_X1    g133(.A(G134gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G127gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n338));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(KEYINPUT1), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n310), .A2(new_n320), .A3(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n321), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n332), .A2(new_n340), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n310), .A2(new_n320), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT4), .B1(new_n341), .B2(new_n321), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n303), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT39), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n302), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n341), .B(new_n321), .ZN(new_n356));
  INV_X1    g155(.A(new_n303), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT39), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n303), .A3(new_n352), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n356), .B2(new_n357), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n346), .A2(new_n352), .A3(new_n364), .A4(new_n303), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n301), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n361), .A2(new_n362), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n289), .A2(new_n297), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371));
  INV_X1    g170(.A(G50gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n214), .A2(new_n267), .A3(new_n321), .A4(new_n216), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n322), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n343), .A2(new_n267), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n343), .A2(KEYINPUT80), .A3(new_n267), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n217), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G228gat), .ZN(new_n385));
  INV_X1    g184(.A(G233gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n377), .A2(new_n388), .A3(new_n322), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n379), .A2(new_n384), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n217), .A2(new_n380), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n210), .B1(new_n212), .B2(new_n211), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n209), .A2(new_n213), .A3(KEYINPUT78), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n396), .B2(new_n349), .ZN(new_n397));
  INV_X1    g196(.A(new_n387), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G22gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n376), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n377), .A2(new_n388), .A3(new_n322), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n388), .B1(new_n377), .B2(new_n322), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n380), .A2(new_n381), .B1(new_n216), .B2(new_n214), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n398), .B1(new_n406), .B2(new_n383), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n405), .A2(new_n407), .B1(new_n398), .B2(new_n397), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G22gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n375), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n390), .B2(new_n399), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT82), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n399), .A3(new_n411), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n376), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n417), .A2(new_n418), .A3(new_n413), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n410), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n270), .A2(KEYINPUT37), .A3(new_n273), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n421), .A2(new_n278), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT37), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n274), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g224(.A(KEYINPUT85), .B(KEYINPUT37), .C1(new_n270), .C2(new_n273), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n366), .A2(new_n367), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n302), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n368), .A2(KEYINPUT76), .A3(KEYINPUT6), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n368), .A2(KEYINPUT6), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n366), .A2(new_n301), .A3(new_n367), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n280), .A2(new_n282), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n422), .B(new_n438), .C1(new_n425), .C2(new_n426), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n428), .A2(new_n436), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n370), .A2(new_n420), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n429), .A2(new_n302), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n435), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n368), .A2(KEYINPUT76), .A3(KEYINPUT6), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT76), .B1(new_n368), .B2(KEYINPUT6), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n293), .A3(new_n296), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n412), .A2(KEYINPUT82), .A3(new_n414), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n418), .B1(new_n417), .B2(new_n413), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n449), .A2(new_n450), .B1(new_n409), .B2(new_n402), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n234), .A2(KEYINPUT25), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n227), .A2(new_n228), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n245), .B1(new_n222), .B2(new_n223), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n247), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n240), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n232), .A2(new_n238), .A3(new_n235), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(new_n234), .A3(new_n235), .A4(new_n232), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n457), .A2(new_n460), .B1(new_n221), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n257), .A2(new_n263), .A3(new_n264), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n341), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n466), .B(KEYINPUT64), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n249), .A2(new_n347), .A3(new_n265), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT34), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n465), .A2(new_n472), .A3(new_n468), .A4(new_n469), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G15gat), .B(G43gat), .Z(new_n475));
  XNOR2_X1  g274(.A(G71gat), .B(G99gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n469), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n347), .B1(new_n249), .B2(new_n265), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n467), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n468), .B1(new_n465), .B2(new_n469), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n477), .B1(new_n485), .B2(KEYINPUT33), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n471), .A3(new_n473), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(KEYINPUT32), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n484), .B2(new_n487), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT36), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n490), .A2(new_n491), .B1(KEYINPUT70), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n486), .B1(new_n471), .B2(new_n473), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n474), .A2(new_n483), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n488), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n448), .A2(new_n451), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n289), .A2(new_n297), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n497), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n451), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n420), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT35), .B1(new_n508), .B2(new_n448), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n441), .A2(new_n501), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT87), .ZN(new_n511));
  INV_X1    g310(.A(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n512), .A3(new_n513), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n514), .A2(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G43gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n372), .ZN(new_n521));
  NAND2_X1  g320(.A1(G43gat), .A2(G50gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(new_n528), .C1(new_n524), .C2(new_n519), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n519), .A2(KEYINPUT88), .A3(new_n524), .A4(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(G1gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT16), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(G1gat), .B2(new_n533), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G8gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n529), .A2(new_n530), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n532), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n538), .A2(new_n529), .A3(new_n530), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n544), .B(KEYINPUT13), .Z(new_n547));
  NOR2_X1   g346(.A1(new_n539), .A2(new_n531), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n538), .B1(new_n529), .B2(new_n530), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G169gat), .B(G197gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT12), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n546), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(KEYINPUT90), .A3(new_n561), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n550), .A3(new_n546), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n556), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n510), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G57gat), .B(G64gat), .Z(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(KEYINPUT92), .A3(new_n573), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G71gat), .B(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n582), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(KEYINPUT93), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G231gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n386), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT20), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n594), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n591), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n590), .B2(new_n591), .ZN(new_n602));
  AOI211_X1 g401(.A(KEYINPUT21), .B(new_n594), .C1(new_n588), .C2(new_n589), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT95), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT21), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n539), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n608), .A3(new_n539), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n612), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n613), .B1(new_n616), .B2(new_n610), .ZN(new_n617));
  INV_X1    g416(.A(new_n606), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n604), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n607), .A2(new_n615), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n615), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n601), .A2(new_n604), .A3(new_n618), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n618), .B1(new_n601), .B2(new_n604), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT7), .ZN(new_n628));
  XOR2_X1   g427(.A(G99gat), .B(G106gat), .Z(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  INV_X1    g430(.A(G92gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(KEYINPUT8), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n629), .B1(new_n628), .B2(new_n633), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n626), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(KEYINPUT98), .A3(new_n634), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n532), .A2(new_n542), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n637), .A2(new_n639), .A3(new_n529), .A4(new_n530), .ZN(new_n642));
  NAND3_X1  g441(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n642), .A2(KEYINPUT99), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT99), .B1(new_n642), .B2(new_n643), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n641), .B(new_n649), .C1(new_n644), .C2(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT96), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT97), .ZN(new_n654));
  XNOR2_X1  g453(.A(G190gat), .B(G218gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n654), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n648), .A2(new_n650), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n625), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n635), .A2(new_n636), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n588), .B2(new_n589), .ZN(new_n667));
  INV_X1    g466(.A(new_n586), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n628), .A2(new_n633), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  INV_X1    g469(.A(new_n629), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n664), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(KEYINPUT102), .B(new_n664), .C1(new_n667), .C2(new_n673), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n590), .A2(new_n665), .ZN(new_n685));
  INV_X1    g484(.A(new_n673), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT10), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n590), .A2(new_n687), .A3(new_n640), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n684), .B1(new_n690), .B2(new_n663), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n676), .A2(KEYINPUT103), .A3(new_n677), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n680), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n663), .B(KEYINPUT104), .Z(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n688), .B2(new_n689), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n684), .B1(new_n678), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n662), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n570), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n447), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n534), .ZN(G1324gat));
  INV_X1    g500(.A(new_n502), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n570), .A2(new_n702), .A3(new_n698), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(G8gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT16), .B(G8gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT42), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT42), .B2(new_n706), .ZN(G1325gat));
  INV_X1    g507(.A(G15gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n493), .A2(new_n500), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n699), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n699), .B2(new_n503), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(G1326gat));
  NAND3_X1  g515(.A1(new_n570), .A2(new_n451), .A3(new_n698), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT106), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  NOR2_X1   g519(.A1(new_n510), .A2(new_n661), .ZN(new_n721));
  INV_X1    g520(.A(new_n625), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n693), .A2(new_n696), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n569), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n721), .A2(new_n512), .A3(new_n436), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT44), .B1(new_n510), .B2(new_n661), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n289), .A2(new_n297), .A3(new_n369), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n432), .A2(new_n433), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n439), .A2(new_n731), .A3(new_n444), .A4(new_n437), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n420), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n501), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n506), .A2(new_n509), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n661), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n729), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n725), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n512), .B1(new_n742), .B2(new_n436), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT108), .B1(new_n728), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n742), .A2(new_n436), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n745), .B(new_n727), .C1(new_n746), .C2(new_n512), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1328gat));
  AND2_X1   g547(.A1(new_n721), .A2(new_n725), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n513), .A3(new_n702), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT46), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n750), .A2(new_n754), .A3(KEYINPUT46), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n750), .B2(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n702), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G36gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n753), .A2(new_n757), .A3(new_n759), .ZN(G1329gat));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  INV_X1    g560(.A(new_n710), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n741), .A2(new_n762), .A3(new_n725), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(new_n520), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n520), .A3(new_n507), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n763), .B2(new_n520), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI221_X1 g567(.A(new_n765), .B1(new_n761), .B2(KEYINPUT47), .C1(new_n763), .C2(new_n520), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(G1330gat));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n737), .B2(new_n738), .ZN(new_n773));
  INV_X1    g572(.A(new_n739), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n661), .B(new_n774), .C1(new_n735), .C2(new_n736), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n451), .B(new_n725), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(G50gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n738), .A2(new_n372), .A3(new_n451), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n510), .A2(new_n569), .A3(new_n724), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n771), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n771), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n372), .B1(new_n776), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n741), .A2(KEYINPUT112), .A3(new_n451), .A4(new_n725), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT113), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n776), .A2(new_n783), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(G50gat), .A3(new_n785), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n789), .B2(new_n781), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n780), .B1(new_n786), .B2(new_n790), .ZN(G1331gat));
  INV_X1    g590(.A(new_n569), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n662), .A2(new_n792), .A3(new_n723), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n737), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n436), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g596(.A1(new_n794), .A2(new_n502), .ZN(new_n798));
  NOR2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  AND2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n798), .B2(new_n799), .ZN(G1333gat));
  NAND3_X1  g601(.A1(new_n795), .A2(G71gat), .A3(new_n762), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT114), .B1(new_n794), .B2(new_n503), .ZN(new_n804));
  INV_X1    g603(.A(G71gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n794), .A2(KEYINPUT114), .A3(new_n503), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n808), .B(new_n809), .Z(G1334gat));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n451), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g611(.A1(new_n792), .A2(new_n625), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n697), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n729), .B2(new_n740), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n436), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n721), .A2(KEYINPUT51), .A3(new_n813), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n721), .B2(new_n813), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n697), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n436), .A2(new_n631), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n631), .A2(new_n816), .B1(new_n819), .B2(new_n820), .ZN(G1336gat));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n702), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G92gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n502), .A2(G92gat), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n697), .B(new_n825), .C1(new_n817), .C2(new_n818), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g627(.A(G99gat), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n815), .A2(new_n762), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(KEYINPUT117), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(KEYINPUT117), .B2(new_n830), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n507), .A2(new_n829), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n819), .B2(new_n833), .ZN(G1338gat));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  INV_X1    g634(.A(G106gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n697), .A2(new_n836), .A3(new_n451), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT119), .Z(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n817), .B2(new_n818), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n815), .A2(new_n451), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT120), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G106gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n840), .A2(KEYINPUT120), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n835), .B(new_n839), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n836), .B1(new_n815), .B2(new_n451), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(KEYINPUT118), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n839), .B1(new_n845), .B2(KEYINPUT118), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT53), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(G1339gat));
  AND4_X1   g648(.A1(new_n569), .A2(new_n723), .A3(new_n625), .A4(new_n661), .ZN(new_n850));
  INV_X1    g649(.A(new_n565), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT90), .B1(new_n560), .B2(new_n561), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n558), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n548), .A2(new_n549), .ZN(new_n854));
  INV_X1    g653(.A(new_n547), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT121), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857));
  NOR4_X1   g656(.A1(new_n548), .A2(new_n549), .A3(new_n857), .A4(new_n547), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n543), .A2(new_n545), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(G229gat), .A3(G233gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n555), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n697), .A2(new_n863), .A3(new_n661), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n660), .B(new_n659), .C1(new_n853), .C2(new_n862), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n648), .A2(new_n650), .A3(new_n657), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n657), .B1(new_n648), .B2(new_n650), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n566), .B(new_n568), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n693), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n683), .B1(new_n695), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n667), .A2(new_n673), .A3(KEYINPUT10), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n590), .A2(new_n687), .A3(new_n640), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n663), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT54), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT55), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n871), .B2(new_n876), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n864), .B1(new_n869), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n850), .B1(new_n882), .B2(new_n722), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n451), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n702), .A2(new_n447), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n507), .A3(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(new_n327), .A3(new_n569), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n883), .A2(new_n447), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n502), .A3(new_n504), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n792), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n891), .B2(new_n327), .ZN(G1340gat));
  NOR3_X1   g691(.A1(new_n886), .A2(new_n325), .A3(new_n723), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n697), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n325), .ZN(G1341gat));
  OAI21_X1  g694(.A(G127gat), .B1(new_n886), .B2(new_n722), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n625), .A2(new_n333), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n889), .B2(new_n897), .ZN(G1342gat));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n335), .A3(new_n738), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n900));
  OAI21_X1  g699(.A(G134gat), .B1(new_n886), .B2(new_n661), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G1343gat));
  XOR2_X1   g702(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n883), .B2(new_n420), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n871), .A2(new_n876), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT55), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n878), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n910), .A2(new_n693), .A3(new_n865), .A4(new_n868), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n625), .B1(new_n911), .B2(new_n864), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n907), .B(new_n451), .C1(new_n912), .C2(new_n850), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n762), .A2(new_n702), .A3(new_n447), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n906), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G141gat), .B1(new_n915), .B2(new_n569), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n702), .A2(new_n762), .A3(new_n420), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n888), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n792), .A2(new_n311), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g720(.A(new_n918), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n313), .A3(new_n697), .ZN(new_n923));
  XOR2_X1   g722(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n924));
  NAND2_X1  g723(.A1(new_n914), .A2(new_n697), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n907), .B1(new_n883), .B2(new_n420), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n451), .B(new_n905), .C1(new_n912), .C2(new_n850), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n928), .B2(new_n313), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  INV_X1    g729(.A(new_n915), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT59), .B(new_n313), .C1(new_n931), .C2(new_n697), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n923), .B1(new_n930), .B2(new_n932), .ZN(G1345gat));
  NAND3_X1  g732(.A1(new_n922), .A2(KEYINPUT125), .A3(new_n625), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n918), .B2(new_n722), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n317), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(G155gat), .A3(new_n625), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(G1346gat));
  AOI21_X1  g738(.A(G162gat), .B1(new_n922), .B2(new_n738), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n915), .A2(new_n318), .A3(new_n661), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(G1347gat));
  NAND2_X1  g741(.A1(new_n702), .A2(new_n447), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n883), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n504), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(G169gat), .B1(new_n946), .B2(new_n792), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n943), .B(KEYINPUT126), .Z(new_n948));
  AND3_X1   g747(.A1(new_n884), .A2(new_n948), .A3(new_n507), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n569), .A2(new_n230), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1348gat));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n231), .A3(new_n697), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n949), .A2(new_n697), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n231), .ZN(G1349gat));
  AOI21_X1  g753(.A(new_n225), .B1(new_n949), .B2(new_n625), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n258), .A2(new_n260), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n946), .A2(new_n958), .A3(new_n625), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT60), .A4(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n962));
  INV_X1    g761(.A(new_n959), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n961), .B(new_n962), .C1(new_n963), .C2(new_n955), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n960), .A2(new_n964), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n946), .A2(new_n226), .A3(new_n738), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n738), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G190gat), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NOR2_X1   g770(.A1(new_n762), .A2(new_n420), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n944), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974), .B2(new_n792), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n948), .A2(new_n710), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n976), .B1(new_n927), .B2(new_n926), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n792), .A2(G197gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NOR2_X1   g778(.A1(new_n723), .A2(G204gat), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT62), .B1(new_n973), .B2(new_n981), .ZN(new_n982));
  OR3_X1    g781(.A1(new_n973), .A2(KEYINPUT62), .A3(new_n981), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n977), .A2(new_n697), .ZN(new_n984));
  INV_X1    g783(.A(G204gat), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n985), .ZN(G1353gat));
  OR3_X1    g785(.A1(new_n973), .A2(G211gat), .A3(new_n722), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n977), .A2(new_n625), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  INV_X1    g790(.A(G218gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n992), .A3(new_n738), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n977), .A2(new_n738), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n994), .B2(new_n992), .ZN(G1355gat));
endmodule


