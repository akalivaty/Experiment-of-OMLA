

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836;

  XNOR2_X1 U380 ( .A(n629), .B(n628), .ZN(n763) );
  XNOR2_X1 U381 ( .A(n452), .B(n621), .ZN(n833) );
  AND2_X1 U382 ( .A1(n417), .A2(n366), .ZN(n360) );
  INV_X1 U383 ( .A(G953), .ZN(n409) );
  INV_X2 U384 ( .A(G953), .ZN(n567) );
  XNOR2_X2 U385 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n512) );
  AND2_X2 U386 ( .A1(n494), .A2(n491), .ZN(n441) );
  XNOR2_X2 U387 ( .A(n613), .B(KEYINPUT94), .ZN(n644) );
  NAND2_X2 U388 ( .A1(n510), .A2(n411), .ZN(n509) );
  AND2_X1 U389 ( .A1(n398), .A2(n396), .ZN(n395) );
  NAND2_X1 U390 ( .A1(n384), .A2(n383), .ZN(n498) );
  NOR2_X1 U391 ( .A1(n388), .A2(n386), .ZN(n496) );
  NOR2_X1 U392 ( .A1(n388), .A2(n387), .ZN(n825) );
  NAND2_X1 U393 ( .A1(n487), .A2(n485), .ZN(n388) );
  NAND2_X1 U394 ( .A1(n483), .A2(KEYINPUT48), .ZN(n484) );
  AND2_X1 U395 ( .A1(n486), .A2(n697), .ZN(n485) );
  XNOR2_X1 U396 ( .A(n669), .B(KEYINPUT40), .ZN(n834) );
  AND2_X1 U397 ( .A1(n689), .A2(n756), .ZN(n669) );
  NOR2_X1 U398 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U399 ( .A1(n367), .A2(n375), .ZN(n374) );
  NAND2_X1 U400 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U401 ( .A(n474), .B(n495), .ZN(n615) );
  NAND2_X1 U402 ( .A1(n441), .A2(n492), .ZN(n474) );
  NAND2_X1 U403 ( .A1(n791), .A2(n502), .ZN(n381) );
  XNOR2_X1 U404 ( .A(n660), .B(n503), .ZN(n791) );
  NAND2_X1 U405 ( .A1(n670), .A2(n382), .ZN(n375) );
  AND2_X1 U406 ( .A1(n792), .A2(KEYINPUT41), .ZN(n376) );
  AND2_X1 U407 ( .A1(n634), .A2(n635), .ZN(n756) );
  NAND2_X1 U408 ( .A1(n422), .A2(n421), .ZN(n406) );
  NAND2_X1 U409 ( .A1(n422), .A2(n361), .ZN(n403) );
  NAND2_X1 U410 ( .A1(n361), .A2(KEYINPUT87), .ZN(n405) );
  INV_X1 U411 ( .A(n421), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n553), .B(KEYINPUT4), .ZN(n565) );
  INV_X1 U413 ( .A(KEYINPUT41), .ZN(n382) );
  NAND2_X1 U414 ( .A1(n395), .A2(n393), .ZN(n400) );
  NAND2_X1 U415 ( .A1(n392), .A2(n394), .ZN(n393) );
  NAND2_X1 U416 ( .A1(n464), .A2(n414), .ZN(n463) );
  NAND2_X1 U417 ( .A1(n498), .A2(n496), .ZN(n443) );
  NAND2_X1 U418 ( .A1(n385), .A2(n404), .ZN(n384) );
  INV_X1 U419 ( .A(n509), .ZN(n385) );
  NAND2_X1 U420 ( .A1(n484), .A2(n497), .ZN(n386) );
  INV_X1 U421 ( .A(n484), .ZN(n387) );
  AND2_X1 U422 ( .A1(n472), .A2(n640), .ZN(n641) );
  AND2_X1 U423 ( .A1(n485), .A2(KEYINPUT2), .ZN(n458) );
  NOR2_X1 U424 ( .A1(n834), .A2(n835), .ZN(n674) );
  AND2_X1 U425 ( .A1(n688), .A2(n419), .ZN(n501) );
  NAND2_X1 U426 ( .A1(n446), .A2(n444), .ZN(n452) );
  AND2_X1 U427 ( .A1(n450), .A2(n447), .ZN(n446) );
  NAND2_X1 U428 ( .A1(n372), .A2(n369), .ZN(n802) );
  XNOR2_X1 U429 ( .A(n365), .B(KEYINPUT39), .ZN(n689) );
  NAND2_X1 U430 ( .A1(n482), .A2(n360), .ZN(n365) );
  AND2_X1 U431 ( .A1(n657), .A2(n424), .ZN(n757) );
  NAND2_X1 U432 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U433 ( .A1(n379), .A2(n376), .ZN(n367) );
  NAND2_X1 U434 ( .A1(n615), .A2(n561), .ZN(n563) );
  NAND2_X1 U435 ( .A1(n445), .A2(n617), .ZN(n444) );
  NOR2_X1 U436 ( .A1(n692), .A2(n679), .ZN(n680) );
  INV_X1 U437 ( .A(n377), .ZN(n370) );
  INV_X1 U438 ( .A(n508), .ZN(n507) );
  XNOR2_X1 U439 ( .A(n457), .B(KEYINPUT30), .ZN(n482) );
  NOR2_X1 U440 ( .A1(n775), .A2(n774), .ZN(n504) );
  NOR2_X1 U441 ( .A1(n662), .A2(n790), .ZN(n457) );
  AND2_X1 U442 ( .A1(n397), .A2(n742), .ZN(n396) );
  XNOR2_X1 U443 ( .A(n630), .B(n577), .ZN(n775) );
  OR2_X1 U444 ( .A1(n724), .A2(G472), .ZN(n397) );
  INV_X1 U445 ( .A(n724), .ZN(n394) );
  NOR2_X1 U446 ( .A1(n652), .A2(n663), .ZN(n653) );
  XNOR2_X1 U447 ( .A(n576), .B(G469), .ZN(n630) );
  XNOR2_X1 U448 ( .A(n456), .B(n587), .ZN(n723) );
  XNOR2_X1 U449 ( .A(n436), .B(n556), .ZN(n702) );
  NAND2_X1 U450 ( .A1(n690), .A2(KEYINPUT114), .ZN(n378) );
  XNOR2_X1 U451 ( .A(n551), .B(n552), .ZN(n436) );
  NAND2_X1 U452 ( .A1(n406), .A2(n405), .ZN(n404) );
  NAND2_X1 U453 ( .A1(n790), .A2(n502), .ZN(n380) );
  NAND2_X1 U454 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U455 ( .A1(n421), .A2(KEYINPUT87), .ZN(n402) );
  XNOR2_X1 U456 ( .A(n511), .B(n809), .ZN(n572) );
  XNOR2_X1 U457 ( .A(G110), .B(G128), .ZN(n593) );
  XNOR2_X1 U458 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n522) );
  XNOR2_X1 U459 ( .A(G146), .B(G125), .ZN(n543) );
  XNOR2_X1 U460 ( .A(G137), .B(G116), .ZN(n583) );
  XNOR2_X1 U461 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n511) );
  NAND2_X1 U462 ( .A1(n427), .A2(n468), .ZN(n390) );
  XNOR2_X2 U463 ( .A(n824), .B(G146), .ZN(n456) );
  XNOR2_X2 U464 ( .A(n362), .B(n565), .ZN(n824) );
  NAND2_X1 U465 ( .A1(n364), .A2(n363), .ZN(n362) );
  NAND2_X1 U466 ( .A1(n566), .A2(n564), .ZN(n363) );
  NAND2_X1 U467 ( .A1(n429), .A2(G134), .ZN(n364) );
  NAND2_X1 U468 ( .A1(n482), .A2(n417), .ZN(n668) );
  INV_X1 U469 ( .A(n791), .ZN(n366) );
  NAND2_X1 U470 ( .A1(n370), .A2(n368), .ZN(n788) );
  INV_X1 U471 ( .A(n379), .ZN(n368) );
  NOR2_X1 U472 ( .A1(n379), .A2(KEYINPUT41), .ZN(n371) );
  AND2_X1 U473 ( .A1(n377), .A2(n376), .ZN(n373) );
  NOR2_X1 U474 ( .A1(n791), .A2(n378), .ZN(n377) );
  NAND2_X1 U475 ( .A1(n509), .A2(n401), .ZN(n383) );
  NAND2_X1 U476 ( .A1(n701), .A2(n389), .ZN(n391) );
  INV_X1 U477 ( .A(n390), .ZN(n389) );
  AND2_X1 U478 ( .A1(n701), .A2(n427), .ZN(n407) );
  XNOR2_X2 U479 ( .A(n460), .B(KEYINPUT89), .ZN(n701) );
  NAND2_X1 U480 ( .A1(n467), .A2(n391), .ZN(n466) );
  XNOR2_X2 U481 ( .A(n509), .B(n361), .ZN(n427) );
  INV_X1 U482 ( .A(n431), .ZN(n392) );
  NAND2_X1 U483 ( .A1(n431), .A2(n399), .ZN(n398) );
  AND2_X1 U484 ( .A1(n724), .A2(G472), .ZN(n399) );
  XNOR2_X1 U485 ( .A(n400), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U486 ( .A1(n644), .A2(KEYINPUT44), .ZN(n614) );
  XNOR2_X1 U487 ( .A(n462), .B(n413), .ZN(n408) );
  XNOR2_X1 U488 ( .A(n462), .B(n413), .ZN(n659) );
  NAND2_X1 U489 ( .A1(n465), .A2(n463), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U491 ( .A1(n723), .A2(n602), .ZN(n589) );
  XNOR2_X1 U492 ( .A(G902), .B(KEYINPUT15), .ZN(n646) );
  NOR2_X1 U493 ( .A1(G953), .A2(G237), .ZN(n579) );
  XOR2_X1 U494 ( .A(G137), .B(G140), .Z(n591) );
  NOR2_X1 U495 ( .A1(G237), .A2(G902), .ZN(n527) );
  INV_X1 U496 ( .A(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U497 ( .A1(n449), .A2(n617), .ZN(n448) );
  XNOR2_X1 U498 ( .A(n440), .B(KEYINPUT33), .ZN(n616) );
  NOR2_X1 U499 ( .A1(n651), .A2(n650), .ZN(n663) );
  XNOR2_X1 U500 ( .A(n648), .B(KEYINPUT112), .ZN(n439) );
  INV_X1 U501 ( .A(G902), .ZN(n602) );
  XNOR2_X1 U502 ( .A(G119), .B(KEYINPUT99), .ZN(n594) );
  INV_X1 U503 ( .A(KEYINPUT82), .ZN(n455) );
  XNOR2_X1 U504 ( .A(n674), .B(n673), .ZN(n489) );
  XNOR2_X1 U505 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n673) );
  NAND2_X1 U506 ( .A1(n646), .A2(n499), .ZN(n497) );
  AND2_X1 U507 ( .A1(n412), .A2(n493), .ZN(n491) );
  INV_X1 U508 ( .A(KEYINPUT65), .ZN(n468) );
  XNOR2_X1 U509 ( .A(KEYINPUT7), .B(KEYINPUT108), .ZN(n548) );
  XOR2_X1 U510 ( .A(KEYINPUT107), .B(KEYINPUT9), .Z(n549) );
  XOR2_X1 U511 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n540) );
  XNOR2_X1 U512 ( .A(G140), .B(KEYINPUT106), .ZN(n539) );
  XNOR2_X1 U513 ( .A(G122), .B(G104), .ZN(n537) );
  XOR2_X1 U514 ( .A(G143), .B(G113), .Z(n538) );
  INV_X1 U515 ( .A(KEYINPUT97), .ZN(n479) );
  XNOR2_X1 U516 ( .A(n532), .B(KEYINPUT14), .ZN(n535) );
  NAND2_X1 U517 ( .A1(G237), .A2(G234), .ZN(n532) );
  INV_X1 U518 ( .A(KEYINPUT114), .ZN(n502) );
  INV_X1 U519 ( .A(G210), .ZN(n528) );
  XOR2_X1 U520 ( .A(KEYINPUT5), .B(KEYINPUT102), .Z(n580) );
  INV_X1 U521 ( .A(KEYINPUT103), .ZN(n582) );
  AND2_X1 U522 ( .A1(n448), .A2(n620), .ZN(n447) );
  INV_X1 U523 ( .A(n663), .ZN(n481) );
  XNOR2_X1 U524 ( .A(n557), .B(G478), .ZN(n636) );
  BUF_X1 U525 ( .A(n630), .Z(n656) );
  NAND2_X1 U526 ( .A1(n790), .A2(n531), .ZN(n493) );
  XNOR2_X1 U527 ( .A(n823), .B(n601), .ZN(n725) );
  XOR2_X1 U528 ( .A(n702), .B(KEYINPUT121), .Z(n703) );
  XNOR2_X1 U529 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U530 ( .A(n738), .B(n739), .ZN(n740) );
  NAND2_X1 U531 ( .A1(n705), .A2(G953), .ZN(n742) );
  NOR2_X1 U532 ( .A1(n507), .A2(n681), .ZN(n765) );
  INV_X1 U533 ( .A(KEYINPUT36), .ZN(n438) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT32), .ZN(n718) );
  AND2_X1 U535 ( .A1(n610), .A2(n507), .ZN(n506) );
  AND2_X1 U536 ( .A1(n507), .A2(n623), .ZN(n475) );
  AND2_X1 U537 ( .A1(n494), .A2(n418), .ZN(n410) );
  OR2_X1 U538 ( .A1(n645), .A2(n644), .ZN(n411) );
  OR2_X1 U539 ( .A1(n536), .A2(n651), .ZN(n412) );
  INV_X1 U540 ( .A(n775), .ZN(n508) );
  OR2_X1 U541 ( .A1(n530), .A2(n528), .ZN(n413) );
  AND2_X1 U542 ( .A1(n772), .A2(n468), .ZN(n414) );
  AND2_X1 U543 ( .A1(n579), .A2(G214), .ZN(n415) );
  NOR2_X1 U544 ( .A1(n790), .A2(n531), .ZN(n416) );
  AND2_X1 U545 ( .A1(n664), .A2(n481), .ZN(n417) );
  AND2_X1 U546 ( .A1(n492), .A2(n493), .ZN(n418) );
  AND2_X1 U547 ( .A1(n667), .A2(n717), .ZN(n419) );
  INV_X1 U548 ( .A(G134), .ZN(n564) );
  XNOR2_X1 U549 ( .A(n562), .B(KEYINPUT22), .ZN(n420) );
  XOR2_X1 U550 ( .A(KEYINPUT88), .B(KEYINPUT45), .Z(n421) );
  NAND2_X1 U551 ( .A1(n698), .A2(KEYINPUT87), .ZN(n422) );
  OR2_X1 U552 ( .A1(n700), .A2(KEYINPUT65), .ZN(n423) );
  INV_X1 U553 ( .A(KEYINPUT48), .ZN(n500) );
  INV_X1 U554 ( .A(KEYINPUT87), .ZN(n499) );
  XNOR2_X1 U555 ( .A(n626), .B(KEYINPUT109), .ZN(n662) );
  AND2_X1 U556 ( .A1(n656), .A2(n410), .ZN(n424) );
  NAND2_X1 U557 ( .A1(n498), .A2(n496), .ZN(n425) );
  XNOR2_X1 U558 ( .A(n611), .B(KEYINPUT110), .ZN(n720) );
  INV_X1 U559 ( .A(n407), .ZN(n426) );
  XNOR2_X1 U560 ( .A(n425), .B(KEYINPUT86), .ZN(n428) );
  XNOR2_X1 U561 ( .A(n443), .B(KEYINPUT86), .ZN(n471) );
  INV_X1 U562 ( .A(n566), .ZN(n429) );
  XNOR2_X1 U563 ( .A(n723), .B(n722), .ZN(n724) );
  BUF_X1 U564 ( .A(n615), .Z(n633) );
  NAND2_X1 U565 ( .A1(n465), .A2(n463), .ZN(n431) );
  NAND2_X1 U566 ( .A1(n516), .A2(n543), .ZN(n434) );
  NAND2_X1 U567 ( .A1(n432), .A2(n433), .ZN(n435) );
  NAND2_X1 U568 ( .A1(n435), .A2(n434), .ZN(n517) );
  INV_X1 U569 ( .A(n516), .ZN(n432) );
  INV_X1 U570 ( .A(n543), .ZN(n433) );
  NAND2_X1 U571 ( .A1(n465), .A2(n463), .ZN(n736) );
  NAND2_X1 U572 ( .A1(n437), .A2(n682), .ZN(n442) );
  XNOR2_X1 U573 ( .A(n765), .B(KEYINPUT91), .ZN(n437) );
  XNOR2_X1 U574 ( .A(n680), .B(n438), .ZN(n681) );
  NOR2_X1 U575 ( .A1(n439), .A2(G900), .ZN(n649) );
  OR2_X1 U576 ( .A1(n501), .A2(n500), .ZN(n486) );
  NAND2_X1 U577 ( .A1(n459), .A2(n484), .ZN(n460) );
  XNOR2_X1 U578 ( .A(n678), .B(n455), .ZN(n454) );
  AND2_X1 U579 ( .A1(n454), .A2(n453), .ZN(n505) );
  NAND2_X1 U580 ( .A1(n504), .A2(n678), .ZN(n440) );
  NAND2_X1 U581 ( .A1(n616), .A2(n451), .ZN(n450) );
  NAND2_X1 U582 ( .A1(n490), .A2(n505), .ZN(n477) );
  XNOR2_X2 U583 ( .A(n563), .B(n420), .ZN(n490) );
  NOR2_X1 U584 ( .A1(n442), .A2(n687), .ZN(n688) );
  INV_X1 U585 ( .A(n408), .ZN(n461) );
  NAND2_X1 U586 ( .A1(n471), .A2(n470), .ZN(n469) );
  INV_X1 U587 ( .A(n616), .ZN(n445) );
  INV_X1 U588 ( .A(n633), .ZN(n449) );
  AND2_X1 U589 ( .A1(n633), .A2(n618), .ZN(n451) );
  NOR2_X1 U590 ( .A1(n775), .A2(n777), .ZN(n453) );
  XNOR2_X2 U591 ( .A(n626), .B(n612), .ZN(n678) );
  XNOR2_X1 U592 ( .A(n456), .B(n575), .ZN(n729) );
  XNOR2_X2 U593 ( .A(n589), .B(n588), .ZN(n626) );
  AND2_X1 U594 ( .A1(n458), .A2(n487), .ZN(n459) );
  NAND2_X1 U595 ( .A1(n461), .A2(n416), .ZN(n492) );
  NAND2_X1 U596 ( .A1(n737), .A2(n646), .ZN(n462) );
  INV_X1 U597 ( .A(n428), .ZN(n464) );
  AND2_X2 U598 ( .A1(n469), .A2(n466), .ZN(n465) );
  NAND2_X1 U599 ( .A1(n772), .A2(n423), .ZN(n467) );
  AND2_X1 U600 ( .A1(n700), .A2(KEYINPUT65), .ZN(n470) );
  NAND2_X1 U601 ( .A1(n622), .A2(KEYINPUT44), .ZN(n472) );
  NAND2_X1 U602 ( .A1(n718), .A2(n720), .ZN(n613) );
  XNOR2_X1 U603 ( .A(n473), .B(n590), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n566), .B(n415), .ZN(n473) );
  XNOR2_X1 U605 ( .A(n569), .B(n479), .ZN(n478) );
  XNOR2_X1 U606 ( .A(n478), .B(n570), .ZN(n574) );
  NAND2_X1 U607 ( .A1(n490), .A2(n475), .ZN(n624) );
  XNOR2_X1 U608 ( .A(n476), .B(KEYINPUT93), .ZN(n510) );
  NAND2_X1 U609 ( .A1(n642), .A2(n641), .ZN(n476) );
  XNOR2_X1 U610 ( .A(n518), .B(n519), .ZN(n526) );
  NAND2_X1 U611 ( .A1(n729), .A2(n602), .ZN(n576) );
  XNOR2_X2 U612 ( .A(n480), .B(KEYINPUT70), .ZN(n566) );
  XNOR2_X2 U613 ( .A(G131), .B(KEYINPUT71), .ZN(n480) );
  INV_X1 U614 ( .A(n489), .ZN(n483) );
  NAND2_X1 U615 ( .A1(n489), .A2(n488), .ZN(n487) );
  AND2_X1 U616 ( .A1(n501), .A2(n500), .ZN(n488) );
  NAND2_X1 U617 ( .A1(n490), .A2(n506), .ZN(n611) );
  OR2_X1 U618 ( .A1(n660), .A2(n790), .ZN(n679) );
  NAND2_X1 U619 ( .A1(n659), .A2(n531), .ZN(n494) );
  INV_X1 U620 ( .A(KEYINPUT0), .ZN(n495) );
  INV_X1 U621 ( .A(n833), .ZN(n622) );
  NAND2_X1 U622 ( .A1(n504), .A2(n781), .ZN(n784) );
  XNOR2_X2 U623 ( .A(G143), .B(G128), .ZN(n553) );
  XNOR2_X1 U624 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U625 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U626 ( .A(n572), .B(n571), .ZN(n573) );
  INV_X1 U627 ( .A(n665), .ZN(n620) );
  INV_X1 U628 ( .A(KEYINPUT122), .ZN(n707) );
  INV_X1 U629 ( .A(G101), .ZN(n809) );
  XNOR2_X1 U630 ( .A(G119), .B(G113), .ZN(n513) );
  XNOR2_X1 U631 ( .A(n513), .B(n512), .ZN(n810) );
  XNOR2_X1 U632 ( .A(n810), .B(n572), .ZN(n578) );
  INV_X1 U633 ( .A(n578), .ZN(n519) );
  XNOR2_X2 U634 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n515) );
  NAND2_X1 U635 ( .A1(n567), .A2(G224), .ZN(n514) );
  XNOR2_X1 U636 ( .A(n517), .B(n565), .ZN(n518) );
  XNOR2_X1 U637 ( .A(G122), .B(G116), .ZN(n521) );
  INV_X1 U638 ( .A(G107), .ZN(n520) );
  XNOR2_X1 U639 ( .A(n521), .B(n520), .ZN(n555) );
  INV_X1 U640 ( .A(n555), .ZN(n523) );
  XNOR2_X1 U641 ( .A(n523), .B(n522), .ZN(n525) );
  XNOR2_X1 U642 ( .A(KEYINPUT77), .B(G110), .ZN(n524) );
  XNOR2_X1 U643 ( .A(n524), .B(G104), .ZN(n569) );
  XNOR2_X1 U644 ( .A(n525), .B(n569), .ZN(n812) );
  XNOR2_X1 U645 ( .A(n526), .B(n812), .ZN(n737) );
  XNOR2_X1 U646 ( .A(n527), .B(KEYINPUT76), .ZN(n530) );
  INV_X1 U647 ( .A(G214), .ZN(n529) );
  OR2_X1 U648 ( .A1(n530), .A2(n529), .ZN(n690) );
  INV_X1 U649 ( .A(n690), .ZN(n790) );
  INV_X1 U650 ( .A(KEYINPUT19), .ZN(n531) );
  NAND2_X1 U651 ( .A1(G902), .A2(n535), .ZN(n533) );
  XNOR2_X1 U652 ( .A(KEYINPUT96), .B(n533), .ZN(n647) );
  NOR2_X1 U653 ( .A1(G898), .A2(n409), .ZN(n534) );
  XNOR2_X1 U654 ( .A(KEYINPUT95), .B(n534), .ZN(n813) );
  NOR2_X1 U655 ( .A1(n647), .A2(n813), .ZN(n536) );
  NAND2_X1 U656 ( .A1(G952), .A2(n535), .ZN(n801) );
  NOR2_X1 U657 ( .A1(n801), .A2(G953), .ZN(n651) );
  XNOR2_X1 U658 ( .A(n538), .B(n537), .ZN(n542) );
  XNOR2_X1 U659 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U660 ( .A(n542), .B(n541), .ZN(n545) );
  XNOR2_X1 U661 ( .A(n543), .B(KEYINPUT10), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n545), .B(n544), .ZN(n710) );
  NAND2_X1 U663 ( .A1(n710), .A2(n602), .ZN(n547) );
  XOR2_X1 U664 ( .A(KEYINPUT13), .B(G475), .Z(n546) );
  XNOR2_X1 U665 ( .A(n547), .B(n546), .ZN(n635) );
  XNOR2_X1 U666 ( .A(n549), .B(n548), .ZN(n552) );
  NAND2_X1 U667 ( .A1(G234), .A2(n409), .ZN(n550) );
  XOR2_X1 U668 ( .A(KEYINPUT8), .B(n550), .Z(n598) );
  NAND2_X1 U669 ( .A1(G217), .A2(n598), .ZN(n551) );
  XNOR2_X1 U670 ( .A(n553), .B(G134), .ZN(n554) );
  XNOR2_X1 U671 ( .A(n555), .B(n554), .ZN(n556) );
  NAND2_X1 U672 ( .A1(n702), .A2(n602), .ZN(n557) );
  OR2_X1 U673 ( .A1(n635), .A2(n636), .ZN(n670) );
  NAND2_X1 U674 ( .A1(n646), .A2(G234), .ZN(n558) );
  XNOR2_X1 U675 ( .A(n558), .B(KEYINPUT20), .ZN(n603) );
  AND2_X1 U676 ( .A1(n603), .A2(G221), .ZN(n560) );
  INV_X1 U677 ( .A(KEYINPUT21), .ZN(n559) );
  XNOR2_X1 U678 ( .A(n560), .B(n559), .ZN(n652) );
  NOR2_X1 U679 ( .A1(n670), .A2(n652), .ZN(n561) );
  INV_X1 U680 ( .A(KEYINPUT74), .ZN(n562) );
  NAND2_X1 U681 ( .A1(G227), .A2(n567), .ZN(n568) );
  XOR2_X1 U682 ( .A(n568), .B(KEYINPUT79), .Z(n570) );
  XNOR2_X1 U683 ( .A(n591), .B(G107), .ZN(n571) );
  XNOR2_X1 U684 ( .A(n574), .B(n573), .ZN(n575) );
  INV_X1 U685 ( .A(KEYINPUT1), .ZN(n577) );
  NAND2_X1 U686 ( .A1(n579), .A2(G210), .ZN(n581) );
  XNOR2_X1 U687 ( .A(n581), .B(n580), .ZN(n585) );
  XNOR2_X1 U688 ( .A(n578), .B(n586), .ZN(n587) );
  XOR2_X1 U689 ( .A(KEYINPUT73), .B(G472), .Z(n588) );
  INV_X1 U690 ( .A(n590), .ZN(n592) );
  XNOR2_X1 U691 ( .A(n592), .B(n591), .ZN(n823) );
  XNOR2_X1 U692 ( .A(n593), .B(KEYINPUT23), .ZN(n597) );
  XOR2_X1 U693 ( .A(KEYINPUT24), .B(KEYINPUT98), .Z(n595) );
  XNOR2_X1 U694 ( .A(n595), .B(n594), .ZN(n596) );
  XOR2_X1 U695 ( .A(n597), .B(n596), .Z(n600) );
  NAND2_X1 U696 ( .A1(G221), .A2(n598), .ZN(n599) );
  XNOR2_X1 U697 ( .A(n600), .B(n599), .ZN(n601) );
  NAND2_X1 U698 ( .A1(n725), .A2(n602), .ZN(n609) );
  XNOR2_X1 U699 ( .A(KEYINPUT100), .B(KEYINPUT78), .ZN(n605) );
  NAND2_X1 U700 ( .A1(G217), .A2(n603), .ZN(n604) );
  XNOR2_X1 U701 ( .A(n605), .B(n604), .ZN(n607) );
  XOR2_X1 U702 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n606) );
  XNOR2_X1 U703 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U704 ( .A(n609), .B(n608), .ZN(n654) );
  AND2_X1 U705 ( .A1(n662), .A2(n654), .ZN(n610) );
  INV_X1 U706 ( .A(KEYINPUT6), .ZN(n612) );
  INV_X1 U707 ( .A(n654), .ZN(n777) );
  XNOR2_X1 U708 ( .A(n614), .B(KEYINPUT66), .ZN(n642) );
  INV_X1 U709 ( .A(n652), .ZN(n778) );
  NAND2_X1 U710 ( .A1(n777), .A2(n778), .ZN(n774) );
  XOR2_X1 U711 ( .A(KEYINPUT34), .B(KEYINPUT81), .Z(n617) );
  INV_X1 U712 ( .A(n617), .ZN(n618) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n619) );
  XOR2_X1 U714 ( .A(KEYINPUT111), .B(n619), .Z(n665) );
  XOR2_X1 U715 ( .A(KEYINPUT80), .B(KEYINPUT35), .Z(n621) );
  INV_X1 U716 ( .A(n678), .ZN(n623) );
  XNOR2_X1 U717 ( .A(n624), .B(KEYINPUT92), .ZN(n625) );
  OR2_X1 U718 ( .A1(n625), .A2(n654), .ZN(n746) );
  BUF_X1 U719 ( .A(n626), .Z(n781) );
  OR2_X1 U720 ( .A1(n784), .A2(n449), .ZN(n629) );
  XNOR2_X1 U721 ( .A(KEYINPUT105), .B(KEYINPUT31), .ZN(n627) );
  XNOR2_X1 U722 ( .A(n627), .B(KEYINPUT104), .ZN(n628) );
  INV_X1 U723 ( .A(n774), .ZN(n631) );
  NAND2_X1 U724 ( .A1(n631), .A2(n656), .ZN(n661) );
  NOR2_X1 U725 ( .A1(n661), .A2(n781), .ZN(n632) );
  NAND2_X1 U726 ( .A1(n633), .A2(n632), .ZN(n749) );
  NAND2_X1 U727 ( .A1(n763), .A2(n749), .ZN(n638) );
  INV_X1 U728 ( .A(n636), .ZN(n634) );
  INV_X1 U729 ( .A(n635), .ZN(n637) );
  AND2_X1 U730 ( .A1(n637), .A2(n636), .ZN(n753) );
  NOR2_X1 U731 ( .A1(n756), .A2(n753), .ZN(n684) );
  INV_X1 U732 ( .A(n684), .ZN(n789) );
  NAND2_X1 U733 ( .A1(n638), .A2(n789), .ZN(n639) );
  AND2_X1 U734 ( .A1(n639), .A2(n746), .ZN(n640) );
  INV_X1 U735 ( .A(KEYINPUT44), .ZN(n643) );
  NAND2_X1 U736 ( .A1(n833), .A2(n643), .ZN(n645) );
  INV_X1 U737 ( .A(n646), .ZN(n698) );
  OR2_X1 U738 ( .A1(n409), .A2(n647), .ZN(n648) );
  XOR2_X1 U739 ( .A(KEYINPUT113), .B(n649), .Z(n650) );
  NAND2_X1 U740 ( .A1(n654), .A2(n653), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n662), .A2(n676), .ZN(n655) );
  XNOR2_X1 U742 ( .A(KEYINPUT28), .B(n655), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n671) );
  NOR2_X1 U744 ( .A1(KEYINPUT47), .A2(n684), .ZN(n658) );
  NAND2_X1 U745 ( .A1(n757), .A2(n658), .ZN(n667) );
  BUF_X1 U746 ( .A(n408), .Z(n660) );
  INV_X1 U747 ( .A(n660), .ZN(n694) );
  INV_X1 U748 ( .A(n661), .ZN(n664) );
  NOR2_X1 U749 ( .A1(n665), .A2(n668), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n694), .A2(n666), .ZN(n717) );
  INV_X1 U751 ( .A(n670), .ZN(n792) );
  NOR2_X1 U752 ( .A1(n671), .A2(n802), .ZN(n672) );
  XNOR2_X1 U753 ( .A(n672), .B(KEYINPUT42), .ZN(n835) );
  INV_X1 U754 ( .A(KEYINPUT47), .ZN(n685) );
  OR2_X1 U755 ( .A1(n757), .A2(n685), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n675), .A2(KEYINPUT85), .ZN(n682) );
  INV_X1 U757 ( .A(n756), .ZN(n760) );
  NOR2_X1 U758 ( .A1(n760), .A2(n676), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n692) );
  NOR2_X1 U760 ( .A1(n757), .A2(KEYINPUT85), .ZN(n683) );
  NOR2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n686) );
  NOR2_X1 U762 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U763 ( .A1(n753), .A2(n689), .ZN(n767) );
  INV_X1 U764 ( .A(n767), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n507), .A2(n690), .ZN(n691) );
  NOR2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U767 ( .A(n693), .B(KEYINPUT43), .ZN(n695) );
  NOR2_X1 U768 ( .A1(n695), .A2(n694), .ZN(n716) );
  NOR2_X1 U769 ( .A1(n696), .A2(n716), .ZN(n697) );
  NAND2_X1 U770 ( .A1(n698), .A2(KEYINPUT2), .ZN(n699) );
  XOR2_X1 U771 ( .A(KEYINPUT67), .B(n699), .Z(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n427), .ZN(n772) );
  NAND2_X1 U773 ( .A1(n430), .A2(G478), .ZN(n704) );
  XNOR2_X1 U774 ( .A(n704), .B(n703), .ZN(n706) );
  INV_X1 U775 ( .A(G952), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n706), .A2(n742), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n708), .B(n707), .ZN(G63) );
  NAND2_X1 U778 ( .A1(n736), .A2(G475), .ZN(n712) );
  XOR2_X1 U779 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n709) );
  XNOR2_X1 U780 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n713), .A2(n742), .ZN(n715) );
  INV_X1 U782 ( .A(KEYINPUT60), .ZN(n714) );
  XNOR2_X1 U783 ( .A(n715), .B(n714), .ZN(G60) );
  XOR2_X1 U784 ( .A(G140), .B(n716), .Z(G42) );
  XNOR2_X1 U785 ( .A(n717), .B(G143), .ZN(G45) );
  BUF_X1 U786 ( .A(n718), .Z(n719) );
  XNOR2_X1 U787 ( .A(n719), .B(G119), .ZN(G21) );
  BUF_X1 U788 ( .A(n720), .Z(n721) );
  XNOR2_X1 U789 ( .A(n721), .B(G110), .ZN(G12) );
  XOR2_X1 U790 ( .A(KEYINPUT115), .B(KEYINPUT62), .Z(n722) );
  NAND2_X1 U791 ( .A1(n430), .A2(G217), .ZN(n726) );
  XNOR2_X1 U792 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U793 ( .A1(n727), .A2(n742), .ZN(n728) );
  XNOR2_X1 U794 ( .A(n728), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U795 ( .A1(n431), .A2(G469), .ZN(n733) );
  XOR2_X1 U796 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n730) );
  XNOR2_X1 U797 ( .A(n730), .B(KEYINPUT58), .ZN(n731) );
  XNOR2_X1 U798 ( .A(n729), .B(n731), .ZN(n732) );
  XNOR2_X1 U799 ( .A(n733), .B(n732), .ZN(n735) );
  INV_X1 U800 ( .A(n742), .ZN(n734) );
  NOR2_X1 U801 ( .A1(n735), .A2(n734), .ZN(G54) );
  NAND2_X1 U802 ( .A1(n736), .A2(G210), .ZN(n741) );
  BUF_X1 U803 ( .A(n737), .Z(n738) );
  XOR2_X1 U804 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n739) );
  XNOR2_X1 U805 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U806 ( .A1(n743), .A2(n742), .ZN(n745) );
  XOR2_X1 U807 ( .A(KEYINPUT90), .B(KEYINPUT56), .Z(n744) );
  XNOR2_X1 U808 ( .A(n745), .B(n744), .ZN(G51) );
  XNOR2_X1 U809 ( .A(G101), .B(n746), .ZN(G3) );
  NOR2_X1 U810 ( .A1(n749), .A2(n760), .ZN(n747) );
  XOR2_X1 U811 ( .A(KEYINPUT116), .B(n747), .Z(n748) );
  XNOR2_X1 U812 ( .A(G104), .B(n748), .ZN(G6) );
  INV_X1 U813 ( .A(n753), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n749), .A2(n762), .ZN(n751) );
  XNOR2_X1 U815 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n750) );
  XNOR2_X1 U816 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U817 ( .A(G107), .B(n752), .ZN(G9) );
  XOR2_X1 U818 ( .A(G128), .B(KEYINPUT29), .Z(n755) );
  NAND2_X1 U819 ( .A1(n757), .A2(n753), .ZN(n754) );
  XNOR2_X1 U820 ( .A(n755), .B(n754), .ZN(G30) );
  XOR2_X1 U821 ( .A(G146), .B(KEYINPUT117), .Z(n759) );
  NAND2_X1 U822 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U823 ( .A(n759), .B(n758), .ZN(G48) );
  NOR2_X1 U824 ( .A1(n763), .A2(n760), .ZN(n761) );
  XOR2_X1 U825 ( .A(G113), .B(n761), .Z(G15) );
  NOR2_X1 U826 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U827 ( .A(G116), .B(n764), .Z(G18) );
  XNOR2_X1 U828 ( .A(G125), .B(n765), .ZN(n766) );
  XNOR2_X1 U829 ( .A(n766), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U830 ( .A(G134), .B(KEYINPUT118), .ZN(n768) );
  XNOR2_X1 U831 ( .A(n768), .B(n767), .ZN(G36) );
  NAND2_X1 U832 ( .A1(n825), .A2(n427), .ZN(n770) );
  XOR2_X1 U833 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n769) );
  NAND2_X1 U834 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U835 ( .A(KEYINPUT83), .B(n771), .Z(n773) );
  NAND2_X1 U836 ( .A1(n773), .A2(n426), .ZN(n806) );
  NAND2_X1 U837 ( .A1(n507), .A2(n774), .ZN(n776) );
  XNOR2_X1 U838 ( .A(n776), .B(KEYINPUT50), .ZN(n783) );
  NOR2_X1 U839 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U840 ( .A(KEYINPUT49), .B(n779), .Z(n780) );
  NOR2_X1 U841 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U842 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U843 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U844 ( .A(KEYINPUT51), .B(n786), .ZN(n787) );
  NOR2_X1 U845 ( .A1(n802), .A2(n787), .ZN(n798) );
  NAND2_X1 U846 ( .A1(n789), .A2(n788), .ZN(n795) );
  NAND2_X1 U847 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U848 ( .A1(n793), .A2(n792), .ZN(n794) );
  AND2_X1 U849 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U850 ( .A1(n796), .A2(n445), .ZN(n797) );
  NOR2_X1 U851 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U852 ( .A(n799), .B(KEYINPUT52), .ZN(n800) );
  NOR2_X1 U853 ( .A1(n801), .A2(n800), .ZN(n804) );
  NOR2_X1 U854 ( .A1(n802), .A2(n445), .ZN(n803) );
  NOR2_X1 U855 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U856 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U857 ( .A1(n807), .A2(G953), .ZN(n808) );
  XNOR2_X1 U858 ( .A(n808), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U859 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U860 ( .A(n812), .B(n811), .ZN(n814) );
  NAND2_X1 U861 ( .A1(n814), .A2(n813), .ZN(n821) );
  NAND2_X1 U862 ( .A1(n427), .A2(n409), .ZN(n819) );
  NAND2_X1 U863 ( .A1(G224), .A2(G953), .ZN(n815) );
  XNOR2_X1 U864 ( .A(n815), .B(KEYINPUT61), .ZN(n816) );
  XNOR2_X1 U865 ( .A(KEYINPUT124), .B(n816), .ZN(n817) );
  NAND2_X1 U866 ( .A1(G898), .A2(n817), .ZN(n818) );
  NAND2_X1 U867 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U868 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U869 ( .A(KEYINPUT125), .B(n822), .ZN(G69) );
  XOR2_X1 U870 ( .A(n824), .B(n823), .Z(n827) );
  XOR2_X1 U871 ( .A(n825), .B(n827), .Z(n826) );
  NAND2_X1 U872 ( .A1(n826), .A2(n409), .ZN(n832) );
  XNOR2_X1 U873 ( .A(G227), .B(n827), .ZN(n828) );
  NAND2_X1 U874 ( .A1(n828), .A2(G900), .ZN(n829) );
  XNOR2_X1 U875 ( .A(KEYINPUT126), .B(n829), .ZN(n830) );
  NAND2_X1 U876 ( .A1(G953), .A2(n830), .ZN(n831) );
  NAND2_X1 U877 ( .A1(n832), .A2(n831), .ZN(G72) );
  XNOR2_X1 U878 ( .A(n833), .B(G122), .ZN(G24) );
  XOR2_X1 U879 ( .A(G131), .B(n834), .Z(G33) );
  XNOR2_X1 U880 ( .A(G137), .B(KEYINPUT127), .ZN(n836) );
  XNOR2_X1 U881 ( .A(n836), .B(n835), .ZN(G39) );
endmodule

