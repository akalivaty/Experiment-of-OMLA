

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  XNOR2_X1 U324 ( .A(n304), .B(n303), .ZN(n309) );
  XNOR2_X1 U325 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U326 ( .A(n475), .B(KEYINPUT122), .ZN(n476) );
  NOR2_X1 U327 ( .A1(n518), .A2(n488), .ZN(n444) );
  XOR2_X1 U328 ( .A(n314), .B(n313), .Z(n548) );
  XOR2_X1 U329 ( .A(n318), .B(KEYINPUT4), .Z(n292) );
  XOR2_X1 U330 ( .A(n342), .B(n341), .Z(n293) );
  XOR2_X1 U331 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n294) );
  XNOR2_X1 U332 ( .A(n470), .B(n469), .ZN(n530) );
  INV_X1 U333 ( .A(KEYINPUT95), .ZN(n361) );
  XNOR2_X1 U334 ( .A(n547), .B(n361), .ZN(n365) );
  XNOR2_X1 U335 ( .A(n414), .B(n413), .ZN(n415) );
  NAND2_X1 U336 ( .A1(n365), .A2(n364), .ZN(n366) );
  XNOR2_X1 U337 ( .A(n468), .B(KEYINPUT116), .ZN(n469) );
  XNOR2_X1 U338 ( .A(n416), .B(n415), .ZN(n419) );
  NOR2_X1 U339 ( .A1(n531), .A2(n371), .ZN(n372) );
  INV_X1 U340 ( .A(KEYINPUT55), .ZN(n475) );
  XNOR2_X1 U341 ( .A(n348), .B(n347), .ZN(n571) );
  XNOR2_X1 U342 ( .A(n302), .B(n301), .ZN(n303) );
  INV_X1 U343 ( .A(n571), .ZN(n572) );
  XNOR2_X1 U344 ( .A(n427), .B(n426), .ZN(n454) );
  XNOR2_X1 U345 ( .A(n343), .B(n293), .ZN(n344) );
  XNOR2_X1 U346 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U347 ( .A(n345), .B(n344), .ZN(n346) );
  INV_X1 U348 ( .A(G43GAT), .ZN(n450) );
  INV_X1 U349 ( .A(G29GAT), .ZN(n446) );
  XNOR2_X1 U350 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U351 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U352 ( .A(n482), .B(n481), .ZN(G1349GAT) );
  XNOR2_X1 U353 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT86), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n294), .B(n295), .ZN(n318) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U357 ( .A(n292), .B(n296), .ZN(n304) );
  XOR2_X1 U358 ( .A(G155GAT), .B(G148GAT), .Z(n298) );
  XNOR2_X1 U359 ( .A(G1GAT), .B(G127GAT), .ZN(n297) );
  XNOR2_X1 U360 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U361 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n300) );
  XNOR2_X1 U362 ( .A(G57GAT), .B(KEYINPUT90), .ZN(n299) );
  XNOR2_X1 U363 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U364 ( .A(G85GAT), .B(G162GAT), .Z(n307) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n305), .B(G120GAT), .ZN(n336) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(n336), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U369 ( .A(n309), .B(n308), .Z(n314) );
  XOR2_X1 U370 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n311) );
  XNOR2_X1 U371 ( .A(KEYINPUT1), .B(KEYINPUT88), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U373 ( .A(G134GAT), .B(n312), .ZN(n313) );
  INV_X1 U374 ( .A(n548), .ZN(n569) );
  XOR2_X1 U375 ( .A(G50GAT), .B(G162GAT), .Z(n394) );
  XOR2_X1 U376 ( .A(G148GAT), .B(KEYINPUT72), .Z(n316) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n412) );
  XNOR2_X1 U379 ( .A(n394), .B(n412), .ZN(n317) );
  XOR2_X1 U380 ( .A(G22GAT), .B(G155GAT), .Z(n379) );
  XNOR2_X1 U381 ( .A(n317), .B(n379), .ZN(n322) );
  XOR2_X1 U382 ( .A(n318), .B(G204GAT), .Z(n320) );
  NAND2_X1 U383 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U385 ( .A(n322), .B(n321), .Z(n331) );
  XNOR2_X1 U386 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n323), .B(KEYINPUT85), .ZN(n324) );
  XOR2_X1 U388 ( .A(n324), .B(KEYINPUT84), .Z(n326) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n349) );
  XOR2_X1 U391 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n328) );
  XNOR2_X1 U392 ( .A(G78GAT), .B(KEYINPUT23), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n349), .B(n329), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n473) );
  XNOR2_X1 U396 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n332), .B(KEYINPUT17), .ZN(n333) );
  XOR2_X1 U398 ( .A(n333), .B(KEYINPUT82), .Z(n335) );
  XNOR2_X1 U399 ( .A(G169GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n335), .B(n334), .ZN(n350) );
  XOR2_X1 U401 ( .A(G43GAT), .B(G134GAT), .Z(n404) );
  XNOR2_X1 U402 ( .A(n336), .B(n404), .ZN(n337) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G127GAT), .Z(n386) );
  XNOR2_X1 U404 ( .A(n337), .B(n386), .ZN(n345) );
  XOR2_X1 U405 ( .A(G71GAT), .B(KEYINPUT81), .Z(n339) );
  XNOR2_X1 U406 ( .A(G190GAT), .B(G99GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n340), .B(KEYINPUT20), .ZN(n343) );
  XOR2_X1 U409 ( .A(KEYINPUT80), .B(G176GAT), .Z(n342) );
  NAND2_X1 U410 ( .A1(G227GAT), .A2(G233GAT), .ZN(n341) );
  XOR2_X1 U411 ( .A(n350), .B(n346), .Z(n523) );
  NAND2_X1 U412 ( .A1(n473), .A2(n523), .ZN(n348) );
  XOR2_X1 U413 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n347) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n352) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .Z(n353) );
  XOR2_X1 U419 ( .A(KEYINPUT76), .B(n353), .Z(n393) );
  XOR2_X1 U420 ( .A(n354), .B(n393), .Z(n358) );
  XOR2_X1 U421 ( .A(G64GAT), .B(G92GAT), .Z(n356) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G204GAT), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n421) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(n421), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U426 ( .A(n360), .B(n359), .Z(n508) );
  XNOR2_X1 U427 ( .A(n508), .B(KEYINPUT27), .ZN(n370) );
  NAND2_X1 U428 ( .A1(n571), .A2(n370), .ZN(n547) );
  INV_X1 U429 ( .A(n508), .ZN(n521) );
  NOR2_X1 U430 ( .A1(n523), .A2(n521), .ZN(n362) );
  NOR2_X1 U431 ( .A1(n473), .A2(n362), .ZN(n363) );
  XNOR2_X1 U432 ( .A(KEYINPUT25), .B(n363), .ZN(n364) );
  NAND2_X1 U433 ( .A1(n366), .A2(n569), .ZN(n367) );
  XOR2_X1 U434 ( .A(KEYINPUT96), .B(n367), .Z(n374) );
  XNOR2_X1 U435 ( .A(n473), .B(KEYINPUT66), .ZN(n368) );
  XOR2_X1 U436 ( .A(n368), .B(KEYINPUT28), .Z(n526) );
  INV_X1 U437 ( .A(n526), .ZN(n512) );
  NOR2_X1 U438 ( .A1(n569), .A2(n512), .ZN(n369) );
  NAND2_X1 U439 ( .A1(n370), .A2(n369), .ZN(n531) );
  INV_X1 U440 ( .A(n523), .ZN(n533) );
  XOR2_X1 U441 ( .A(KEYINPUT83), .B(n533), .Z(n371) );
  XOR2_X1 U442 ( .A(KEYINPUT93), .B(n372), .Z(n373) );
  NOR2_X1 U443 ( .A1(n374), .A2(n373), .ZN(n487) );
  XOR2_X1 U444 ( .A(KEYINPUT14), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U445 ( .A(G183GAT), .B(G211GAT), .ZN(n375) );
  XOR2_X1 U446 ( .A(n376), .B(n375), .Z(n390) );
  XOR2_X1 U447 ( .A(KEYINPUT13), .B(G57GAT), .Z(n378) );
  XNOR2_X1 U448 ( .A(G71GAT), .B(G78GAT), .ZN(n377) );
  XNOR2_X1 U449 ( .A(n378), .B(n377), .ZN(n420) );
  XOR2_X1 U450 ( .A(n420), .B(n379), .Z(n381) );
  NAND2_X1 U451 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U453 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n383) );
  XNOR2_X1 U454 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n382) );
  XNOR2_X1 U455 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U456 ( .A(n385), .B(n384), .Z(n388) );
  XOR2_X1 U457 ( .A(G8GAT), .B(G1GAT), .Z(n428) );
  XNOR2_X1 U458 ( .A(n428), .B(n386), .ZN(n387) );
  XNOR2_X1 U459 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U460 ( .A(n390), .B(n389), .ZN(n582) );
  INV_X1 U461 ( .A(n582), .ZN(n483) );
  NOR2_X1 U462 ( .A1(n487), .A2(n483), .ZN(n410) );
  XOR2_X1 U463 ( .A(G29GAT), .B(KEYINPUT7), .Z(n392) );
  XNOR2_X1 U464 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n391) );
  XNOR2_X1 U465 ( .A(n392), .B(n391), .ZN(n429) );
  XOR2_X1 U466 ( .A(n429), .B(n393), .Z(n408) );
  XOR2_X1 U467 ( .A(G99GAT), .B(G85GAT), .Z(n417) );
  XOR2_X1 U468 ( .A(n417), .B(n394), .Z(n396) );
  NAND2_X1 U469 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U470 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U471 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n398) );
  XNOR2_X1 U472 ( .A(G106GAT), .B(G92GAT), .ZN(n397) );
  XOR2_X1 U473 ( .A(n398), .B(n397), .Z(n399) );
  XNOR2_X1 U474 ( .A(n400), .B(n399), .ZN(n406) );
  XOR2_X1 U475 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n402) );
  XNOR2_X1 U476 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n401) );
  XNOR2_X1 U477 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U479 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U480 ( .A(n408), .B(n407), .Z(n559) );
  INV_X1 U481 ( .A(n559), .ZN(n566) );
  XOR2_X1 U482 ( .A(n566), .B(KEYINPUT101), .Z(n409) );
  XNOR2_X1 U483 ( .A(n409), .B(KEYINPUT36), .ZN(n585) );
  NAND2_X1 U484 ( .A1(n410), .A2(n585), .ZN(n411) );
  XOR2_X1 U485 ( .A(KEYINPUT37), .B(n411), .Z(n518) );
  XNOR2_X1 U486 ( .A(n412), .B(KEYINPUT73), .ZN(n416) );
  AND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n414) );
  INV_X1 U488 ( .A(KEYINPUT33), .ZN(n413) );
  XNOR2_X1 U489 ( .A(G120GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U490 ( .A(n419), .B(n418), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U492 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n423) );
  XNOR2_X1 U493 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n422) );
  XOR2_X1 U494 ( .A(n423), .B(n422), .Z(n424) );
  XOR2_X1 U495 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U496 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U498 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n433) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(KEYINPUT29), .ZN(n432) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U501 ( .A(n435), .B(n434), .Z(n443) );
  XOR2_X1 U502 ( .A(G141GAT), .B(G43GAT), .Z(n437) );
  XNOR2_X1 U503 ( .A(G36GAT), .B(G50GAT), .ZN(n436) );
  XNOR2_X1 U504 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U505 ( .A(G15GAT), .B(G113GAT), .Z(n439) );
  XNOR2_X1 U506 ( .A(G22GAT), .B(G197GAT), .ZN(n438) );
  XNOR2_X1 U507 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U508 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U509 ( .A(n443), .B(n442), .Z(n535) );
  NAND2_X1 U510 ( .A1(n454), .A2(n535), .ZN(n488) );
  XOR2_X1 U511 ( .A(KEYINPUT102), .B(n444), .Z(n445) );
  XNOR2_X1 U512 ( .A(KEYINPUT38), .B(n445), .ZN(n501) );
  NOR2_X1 U513 ( .A1(n569), .A2(n501), .ZN(n449) );
  XNOR2_X1 U514 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n447) );
  XNOR2_X1 U515 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U516 ( .A(n449), .B(n448), .ZN(G1328GAT) );
  NOR2_X1 U517 ( .A1(n523), .A2(n501), .ZN(n453) );
  XNOR2_X1 U518 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n451) );
  INV_X1 U519 ( .A(n535), .ZN(n574) );
  XOR2_X1 U520 ( .A(n454), .B(KEYINPUT41), .Z(n553) );
  NOR2_X1 U521 ( .A1(n574), .A2(n553), .ZN(n456) );
  XOR2_X1 U522 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n455) );
  XNOR2_X1 U523 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U524 ( .A(KEYINPUT112), .B(n582), .Z(n563) );
  NOR2_X1 U525 ( .A1(n457), .A2(n563), .ZN(n458) );
  XOR2_X1 U526 ( .A(KEYINPUT114), .B(n458), .Z(n459) );
  NOR2_X1 U527 ( .A1(n566), .A2(n459), .ZN(n460) );
  XNOR2_X1 U528 ( .A(KEYINPUT47), .B(n460), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n483), .A2(n585), .ZN(n461) );
  XNOR2_X1 U530 ( .A(n461), .B(KEYINPUT45), .ZN(n462) );
  XNOR2_X1 U531 ( .A(KEYINPUT65), .B(n462), .ZN(n463) );
  NAND2_X1 U532 ( .A1(n463), .A2(n454), .ZN(n464) );
  XNOR2_X1 U533 ( .A(KEYINPUT115), .B(n464), .ZN(n465) );
  NAND2_X1 U534 ( .A1(n465), .A2(n574), .ZN(n466) );
  NAND2_X1 U535 ( .A1(n467), .A2(n466), .ZN(n470) );
  XOR2_X1 U536 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n468) );
  XNOR2_X1 U537 ( .A(KEYINPUT121), .B(n508), .ZN(n471) );
  NOR2_X1 U538 ( .A1(n530), .A2(n471), .ZN(n472) );
  XNOR2_X1 U539 ( .A(KEYINPUT54), .B(n472), .ZN(n570) );
  NOR2_X1 U540 ( .A1(n473), .A2(n548), .ZN(n474) );
  AND2_X1 U541 ( .A1(n570), .A2(n474), .ZN(n477) );
  NAND2_X1 U542 ( .A1(n478), .A2(n533), .ZN(n562) );
  XOR2_X1 U543 ( .A(n553), .B(KEYINPUT105), .Z(n538) );
  NOR2_X1 U544 ( .A1(n562), .A2(n538), .ZN(n482) );
  XOR2_X1 U545 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n480) );
  XNOR2_X1 U546 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n479) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n490) );
  XOR2_X1 U548 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n485) );
  NAND2_X1 U549 ( .A1(n559), .A2(n483), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(n486) );
  OR2_X1 U551 ( .A1(n487), .A2(n486), .ZN(n503) );
  NOR2_X1 U552 ( .A1(n488), .A2(n503), .ZN(n496) );
  NAND2_X1 U553 ( .A1(n496), .A2(n548), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  XOR2_X1 U555 ( .A(G8GAT), .B(KEYINPUT97), .Z(n492) );
  NAND2_X1 U556 ( .A1(n496), .A2(n508), .ZN(n491) );
  XNOR2_X1 U557 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n494) );
  NAND2_X1 U559 ( .A1(n496), .A2(n533), .ZN(n493) );
  XNOR2_X1 U560 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n498) );
  NAND2_X1 U563 ( .A1(n496), .A2(n512), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n499), .ZN(G1327GAT) );
  NOR2_X1 U566 ( .A1(n521), .A2(n501), .ZN(n500) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  NOR2_X1 U568 ( .A1(n526), .A2(n501), .ZN(n502) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  OR2_X1 U570 ( .A1(n538), .A2(n535), .ZN(n517) );
  NOR2_X1 U571 ( .A1(n517), .A2(n503), .ZN(n513) );
  NAND2_X1 U572 ( .A1(n548), .A2(n513), .ZN(n507) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n505) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n504) );
  XNOR2_X1 U575 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U577 ( .A1(n508), .A2(n513), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n509), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n533), .A2(n513), .ZN(n511) );
  XNOR2_X1 U581 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U585 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  OR2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n569), .A2(n525), .ZN(n519) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n519), .Z(n520) );
  XNOR2_X1 U589 ( .A(KEYINPUT110), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n523), .A2(n525), .ZN(n524) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U595 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n530), .A2(n531), .ZN(n532) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(n534), .B(KEYINPUT117), .Z(n537) );
  INV_X1 U601 ( .A(n537), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n535), .A2(n544), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  NOR2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n544), .A2(n563), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n566), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n530), .A2(n547), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n574), .A2(n558), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n558), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n582), .A2(n558), .ZN(n557) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NOR2_X1 U628 ( .A1(n574), .A2(n562), .ZN(n561) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  INV_X1 U630 ( .A(n562), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n573) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n586) );
  INV_X1 U638 ( .A(n586), .ZN(n581) );
  NOR2_X1 U639 ( .A1(n574), .A2(n581), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n454), .A2(n581), .ZN(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(G218GAT), .B(n589), .Z(G1355GAT) );
endmodule

