

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(n706), .A2(n705), .ZN(n707) );
  OR2_X1 U555 ( .A1(n801), .A2(n800), .ZN(n815) );
  XNOR2_X1 U556 ( .A(n743), .B(KEYINPUT92), .ZN(n523) );
  XNOR2_X1 U557 ( .A(n743), .B(KEYINPUT92), .ZN(n758) );
  AND2_X1 U558 ( .A1(n921), .A2(n812), .ZN(n524) );
  AND2_X1 U559 ( .A1(n689), .A2(G1996), .ZN(n690) );
  INV_X1 U560 ( .A(G2105), .ZN(n527) );
  OR2_X1 U561 ( .A1(n799), .A2(n524), .ZN(n800) );
  NOR2_X1 U562 ( .A1(n628), .A2(G651), .ZN(n651) );
  XOR2_X1 U563 ( .A(KEYINPUT17), .B(n532), .Z(n868) );
  INV_X1 U564 ( .A(KEYINPUT64), .ZN(n535) );
  NOR2_X1 U565 ( .A1(n543), .A2(n542), .ZN(G164) );
  NOR2_X2 U566 ( .A1(G2104), .A2(n527), .ZN(n872) );
  NAND2_X1 U567 ( .A1(G125), .A2(n872), .ZN(n526) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n873) );
  NAND2_X1 U569 ( .A1(G113), .A2(n873), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U571 ( .A1(n527), .A2(G2104), .ZN(n528) );
  XNOR2_X2 U572 ( .A(n528), .B(KEYINPUT65), .ZN(n869) );
  NAND2_X1 U573 ( .A1(G101), .A2(n869), .ZN(n529) );
  XNOR2_X1 U574 ( .A(n529), .B(KEYINPUT23), .ZN(n530) );
  NOR2_X1 U575 ( .A1(n531), .A2(n530), .ZN(n534) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  NAND2_X1 U577 ( .A1(n868), .A2(G137), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X2 U579 ( .A(n536), .B(n535), .ZN(G160) );
  NAND2_X1 U580 ( .A1(n872), .A2(G126), .ZN(n537) );
  XNOR2_X1 U581 ( .A(n537), .B(KEYINPUT82), .ZN(n539) );
  NAND2_X1 U582 ( .A1(G138), .A2(n868), .ZN(n538) );
  NAND2_X1 U583 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U584 ( .A1(G102), .A2(n869), .ZN(n541) );
  NAND2_X1 U585 ( .A1(G114), .A2(n873), .ZN(n540) );
  NAND2_X1 U586 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n628) );
  NAND2_X1 U588 ( .A1(G53), .A2(n651), .ZN(n546) );
  INV_X1 U589 ( .A(G651), .ZN(n547) );
  NOR2_X1 U590 ( .A1(G543), .A2(n547), .ZN(n544) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n544), .Z(n652) );
  NAND2_X1 U592 ( .A1(G65), .A2(n652), .ZN(n545) );
  NAND2_X1 U593 ( .A1(n546), .A2(n545), .ZN(n551) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n647) );
  NAND2_X1 U595 ( .A1(G91), .A2(n647), .ZN(n549) );
  NOR2_X1 U596 ( .A1(n628), .A2(n547), .ZN(n648) );
  NAND2_X1 U597 ( .A1(G78), .A2(n648), .ZN(n548) );
  NAND2_X1 U598 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U599 ( .A1(n551), .A2(n550), .ZN(G299) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  NAND2_X1 U604 ( .A1(G52), .A2(n651), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G64), .A2(n652), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U607 ( .A1(G90), .A2(n647), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G77), .A2(n648), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U611 ( .A1(n558), .A2(n557), .ZN(G171) );
  NAND2_X1 U612 ( .A1(n647), .A2(G89), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G76), .A2(n648), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U616 ( .A(KEYINPUT5), .B(n562), .ZN(n569) );
  XNOR2_X1 U617 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n567) );
  NAND2_X1 U618 ( .A1(G51), .A2(n651), .ZN(n564) );
  NAND2_X1 U619 ( .A1(G63), .A2(n652), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U621 ( .A(n565), .B(KEYINPUT6), .ZN(n566) );
  XNOR2_X1 U622 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U624 ( .A(KEYINPUT7), .B(n570), .ZN(G168) );
  XOR2_X1 U625 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U627 ( .A(n571), .B(KEYINPUT10), .ZN(n572) );
  XNOR2_X1 U628 ( .A(KEYINPUT68), .B(n572), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n817) );
  NAND2_X1 U630 ( .A1(n817), .A2(G567), .ZN(n573) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  INV_X1 U632 ( .A(G860), .ZN(n617) );
  NAND2_X1 U633 ( .A1(n651), .A2(G43), .ZN(n574) );
  XNOR2_X1 U634 ( .A(KEYINPUT70), .B(n574), .ZN(n584) );
  NAND2_X1 U635 ( .A1(n652), .A2(G56), .ZN(n575) );
  XNOR2_X1 U636 ( .A(KEYINPUT14), .B(n575), .ZN(n581) );
  NAND2_X1 U637 ( .A1(n647), .A2(G81), .ZN(n576) );
  XNOR2_X1 U638 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G68), .A2(n648), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(n579), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U643 ( .A(KEYINPUT69), .B(n582), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n930) );
  NOR2_X1 U645 ( .A1(n617), .A2(n930), .ZN(n585) );
  XNOR2_X1 U646 ( .A(n585), .B(KEYINPUT71), .ZN(G153) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U649 ( .A1(G54), .A2(n651), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G79), .A2(n648), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n593) );
  NAND2_X1 U652 ( .A1(n652), .A2(G66), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT72), .ZN(n590) );
  NAND2_X1 U654 ( .A1(G92), .A2(n647), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(KEYINPUT73), .B(n591), .Z(n592) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(KEYINPUT15), .B(n594), .ZN(n931) );
  INV_X1 U659 ( .A(G868), .ZN(n666) );
  NAND2_X1 U660 ( .A1(n931), .A2(n666), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(G284) );
  NOR2_X1 U662 ( .A1(G286), .A2(n666), .ZN(n598) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U664 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n617), .A2(G559), .ZN(n599) );
  INV_X1 U666 ( .A(n931), .ZN(n893) );
  NAND2_X1 U667 ( .A1(n599), .A2(n893), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n930), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G868), .A2(n893), .ZN(n601) );
  NOR2_X1 U671 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U672 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G135), .A2(n868), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n604), .B(KEYINPUT76), .ZN(n612) );
  NAND2_X1 U675 ( .A1(n872), .A2(G123), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G111), .A2(n873), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G99), .A2(n869), .ZN(n608) );
  XNOR2_X1 U680 ( .A(KEYINPUT77), .B(n608), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n978) );
  XOR2_X1 U683 ( .A(G2096), .B(KEYINPUT78), .Z(n613) );
  XNOR2_X1 U684 ( .A(n978), .B(n613), .ZN(n615) );
  INV_X1 U685 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G559), .A2(n893), .ZN(n616) );
  XOR2_X1 U688 ( .A(n930), .B(n616), .Z(n663) );
  NAND2_X1 U689 ( .A1(n617), .A2(n663), .ZN(n624) );
  NAND2_X1 U690 ( .A1(G55), .A2(n651), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G67), .A2(n652), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G93), .A2(n647), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G80), .A2(n648), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n665) );
  XOR2_X1 U697 ( .A(n624), .B(n665), .Z(G145) );
  NAND2_X1 U698 ( .A1(G49), .A2(n651), .ZN(n626) );
  NAND2_X1 U699 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n652), .A2(n627), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U704 ( .A1(G73), .A2(n648), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n631), .B(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U706 ( .A1(G86), .A2(n647), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G48), .A2(n651), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G61), .A2(n652), .ZN(n634) );
  XNOR2_X1 U710 ( .A(KEYINPUT79), .B(n634), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U713 ( .A1(n648), .A2(G72), .ZN(n645) );
  NAND2_X1 U714 ( .A1(G47), .A2(n651), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G60), .A2(n652), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G85), .A2(n647), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT66), .B(n641), .Z(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U721 ( .A(KEYINPUT67), .B(n646), .Z(G290) );
  NAND2_X1 U722 ( .A1(G88), .A2(n647), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G75), .A2(n648), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n656) );
  NAND2_X1 U725 ( .A1(G50), .A2(n651), .ZN(n654) );
  NAND2_X1 U726 ( .A1(G62), .A2(n652), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(KEYINPUT80), .ZN(G166) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(G288), .ZN(n662) );
  XOR2_X1 U731 ( .A(G290), .B(G166), .Z(n658) );
  XNOR2_X1 U732 ( .A(G305), .B(n658), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n665), .B(n659), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(G299), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(n894) );
  XOR2_X1 U736 ( .A(n894), .B(n663), .Z(n664) );
  NOR2_X1 U737 ( .A1(n666), .A2(n664), .ZN(n668) );
  AND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U739 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n669), .B(KEYINPUT81), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n670), .B(KEYINPUT20), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U749 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U750 ( .A1(G96), .A2(n676), .ZN(n823) );
  NAND2_X1 U751 ( .A1(n823), .A2(G2106), .ZN(n680) );
  NAND2_X1 U752 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U753 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U754 ( .A1(G108), .A2(n678), .ZN(n824) );
  NAND2_X1 U755 ( .A1(n824), .A2(G567), .ZN(n679) );
  NAND2_X1 U756 ( .A1(n680), .A2(n679), .ZN(n825) );
  NAND2_X1 U757 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U758 ( .A1(n825), .A2(n681), .ZN(n822) );
  NAND2_X1 U759 ( .A1(n822), .A2(G36), .ZN(G176) );
  XNOR2_X1 U760 ( .A(KEYINPUT83), .B(G166), .ZN(G303) );
  NOR2_X1 U761 ( .A1(G164), .A2(G1384), .ZN(n765) );
  AND2_X1 U762 ( .A1(G40), .A2(n765), .ZN(n682) );
  NAND2_X2 U763 ( .A1(n682), .A2(G160), .ZN(n724) );
  NAND2_X1 U764 ( .A1(G8), .A2(n724), .ZN(n759) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n683) );
  XOR2_X1 U766 ( .A(n683), .B(KEYINPUT24), .Z(n684) );
  NOR2_X1 U767 ( .A1(n759), .A2(n684), .ZN(n764) );
  INV_X1 U768 ( .A(n724), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n708), .A2(G2072), .ZN(n685) );
  XOR2_X1 U770 ( .A(KEYINPUT27), .B(n685), .Z(n687) );
  NAND2_X1 U771 ( .A1(G1956), .A2(n724), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n701) );
  NAND2_X1 U773 ( .A1(G299), .A2(n701), .ZN(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT28), .B(n688), .Z(n706) );
  INV_X1 U775 ( .A(n724), .ZN(n689) );
  XOR2_X1 U776 ( .A(n690), .B(KEYINPUT26), .Z(n693) );
  AND2_X1 U777 ( .A1(n724), .A2(G1341), .ZN(n691) );
  NOR2_X1 U778 ( .A1(n691), .A2(n930), .ZN(n692) );
  AND2_X1 U779 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n724), .ZN(n695) );
  NAND2_X1 U781 ( .A1(G2067), .A2(n708), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n698) );
  NOR2_X1 U783 ( .A1(n931), .A2(n698), .ZN(n696) );
  NOR2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n700) );
  AND2_X1 U785 ( .A1(n931), .A2(n698), .ZN(n699) );
  NOR2_X1 U786 ( .A1(n700), .A2(n699), .ZN(n703) );
  NOR2_X1 U787 ( .A1(G299), .A2(n701), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U789 ( .A(n704), .B(KEYINPUT90), .ZN(n705) );
  XNOR2_X1 U790 ( .A(n707), .B(KEYINPUT29), .ZN(n712) );
  XOR2_X1 U791 ( .A(KEYINPUT25), .B(G2078), .Z(n939) );
  NOR2_X1 U792 ( .A1(n939), .A2(n724), .ZN(n710) );
  NOR2_X1 U793 ( .A1(n708), .A2(G1961), .ZN(n709) );
  NOR2_X1 U794 ( .A1(n710), .A2(n709), .ZN(n717) );
  OR2_X1 U795 ( .A1(n717), .A2(G301), .ZN(n711) );
  NAND2_X1 U796 ( .A1(n712), .A2(n711), .ZN(n722) );
  NOR2_X1 U797 ( .A1(G1966), .A2(n759), .ZN(n736) );
  NOR2_X1 U798 ( .A1(G2084), .A2(n724), .ZN(n737) );
  NOR2_X1 U799 ( .A1(n736), .A2(n737), .ZN(n713) );
  NAND2_X1 U800 ( .A1(G8), .A2(n713), .ZN(n714) );
  XNOR2_X1 U801 ( .A(KEYINPUT30), .B(n714), .ZN(n715) );
  NOR2_X1 U802 ( .A1(G168), .A2(n715), .ZN(n716) );
  XNOR2_X1 U803 ( .A(n716), .B(KEYINPUT91), .ZN(n719) );
  NAND2_X1 U804 ( .A1(n717), .A2(G301), .ZN(n718) );
  NAND2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U806 ( .A(n720), .B(KEYINPUT31), .ZN(n721) );
  NAND2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n734) );
  AND2_X1 U808 ( .A1(G286), .A2(G8), .ZN(n723) );
  NAND2_X1 U809 ( .A1(n734), .A2(n723), .ZN(n731) );
  INV_X1 U810 ( .A(G8), .ZN(n729) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n759), .ZN(n726) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U814 ( .A1(G303), .A2(n727), .ZN(n728) );
  OR2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n731), .A2(n730), .ZN(n733) );
  INV_X1 U817 ( .A(KEYINPUT32), .ZN(n732) );
  XNOR2_X1 U818 ( .A(n733), .B(n732), .ZN(n742) );
  INV_X1 U819 ( .A(n734), .ZN(n735) );
  NOR2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n740) );
  NAND2_X1 U821 ( .A1(G8), .A2(n737), .ZN(n738) );
  XOR2_X1 U822 ( .A(KEYINPUT89), .B(n738), .Z(n739) );
  NAND2_X1 U823 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U824 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n919) );
  NOR2_X1 U826 ( .A1(G303), .A2(G1971), .ZN(n744) );
  XOR2_X1 U827 ( .A(n744), .B(KEYINPUT93), .Z(n745) );
  NOR2_X1 U828 ( .A1(n919), .A2(n745), .ZN(n746) );
  XNOR2_X1 U829 ( .A(n746), .B(KEYINPUT94), .ZN(n747) );
  NAND2_X1 U830 ( .A1(n758), .A2(n747), .ZN(n750) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n916) );
  INV_X1 U832 ( .A(n916), .ZN(n748) );
  NOR2_X1 U833 ( .A1(n759), .A2(n748), .ZN(n749) );
  AND2_X1 U834 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n751), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n919), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U837 ( .A1(n752), .A2(n759), .ZN(n753) );
  NOR2_X1 U838 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n926) );
  NAND2_X1 U840 ( .A1(n755), .A2(n926), .ZN(n762) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n523), .A2(n757), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U845 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U846 ( .A1(n764), .A2(n763), .ZN(n801) );
  NAND2_X1 U847 ( .A1(G40), .A2(G160), .ZN(n766) );
  NOR2_X1 U848 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U849 ( .A(n767), .B(KEYINPUT84), .ZN(n812) );
  INV_X1 U850 ( .A(n812), .ZN(n798) );
  XNOR2_X1 U851 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NAND2_X1 U852 ( .A1(n869), .A2(G104), .ZN(n768) );
  XNOR2_X1 U853 ( .A(KEYINPUT85), .B(n768), .ZN(n771) );
  NAND2_X1 U854 ( .A1(n868), .A2(G140), .ZN(n769) );
  XOR2_X1 U855 ( .A(KEYINPUT86), .B(n769), .Z(n770) );
  NOR2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U857 ( .A(n772), .B(KEYINPUT34), .ZN(n777) );
  NAND2_X1 U858 ( .A1(G128), .A2(n872), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G116), .A2(n873), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U861 ( .A(KEYINPUT35), .B(n775), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U863 ( .A(n778), .B(KEYINPUT36), .Z(n890) );
  OR2_X1 U864 ( .A1(n810), .A2(n890), .ZN(n980) );
  NOR2_X1 U865 ( .A1(n798), .A2(n980), .ZN(n779) );
  XOR2_X1 U866 ( .A(KEYINPUT87), .B(n779), .Z(n808) );
  INV_X1 U867 ( .A(G1991), .ZN(n788) );
  NAND2_X1 U868 ( .A1(G119), .A2(n872), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G131), .A2(n868), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G95), .A2(n869), .ZN(n783) );
  NAND2_X1 U872 ( .A1(G107), .A2(n873), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U875 ( .A(KEYINPUT88), .B(n786), .Z(n867) );
  INV_X1 U876 ( .A(n867), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n797) );
  NAND2_X1 U878 ( .A1(G129), .A2(n872), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G117), .A2(n873), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n869), .A2(G105), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n868), .A2(G141), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n885) );
  AND2_X1 U886 ( .A1(n885), .A2(G1996), .ZN(n796) );
  NOR2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n973) );
  NOR2_X1 U888 ( .A1(n798), .A2(n973), .ZN(n804) );
  OR2_X1 U889 ( .A1(n808), .A2(n804), .ZN(n799) );
  XNOR2_X1 U890 ( .A(G1986), .B(G290), .ZN(n921) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n885), .ZN(n970) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U893 ( .A1(G1991), .A2(n867), .ZN(n976) );
  NOR2_X1 U894 ( .A1(n802), .A2(n976), .ZN(n803) );
  NOR2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U896 ( .A1(n970), .A2(n805), .ZN(n806) );
  XOR2_X1 U897 ( .A(KEYINPUT39), .B(n806), .Z(n807) );
  NOR2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U899 ( .A(n809), .B(KEYINPUT95), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n810), .A2(n890), .ZN(n987) );
  NAND2_X1 U901 ( .A1(n811), .A2(n987), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U904 ( .A(n816), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U905 ( .A1(n817), .A2(G2106), .ZN(n818) );
  XNOR2_X1 U906 ( .A(n818), .B(KEYINPUT96), .ZN(G217) );
  NAND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n819) );
  XNOR2_X1 U908 ( .A(KEYINPUT97), .B(n819), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n820), .A2(G661), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U911 ( .A1(n822), .A2(n821), .ZN(G188) );
  INV_X1 U913 ( .A(G120), .ZN(G236) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  INV_X1 U915 ( .A(G69), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n824), .A2(n823), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  INV_X1 U918 ( .A(n825), .ZN(G319) );
  XOR2_X1 U919 ( .A(G1976), .B(G1971), .Z(n827) );
  XNOR2_X1 U920 ( .A(G1986), .B(G1966), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n827), .B(n826), .ZN(n837) );
  XOR2_X1 U922 ( .A(KEYINPUT99), .B(KEYINPUT41), .Z(n829) );
  XNOR2_X1 U923 ( .A(G1991), .B(G2474), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U925 ( .A(G1981), .B(G1956), .Z(n831) );
  XNOR2_X1 U926 ( .A(G1996), .B(G1961), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U928 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U929 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U931 ( .A(n837), .B(n836), .Z(G229) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U933 ( .A(G2090), .B(G2678), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U935 ( .A(n840), .B(G2100), .Z(n842) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT98), .Z(n844) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U941 ( .A(n846), .B(n845), .ZN(G227) );
  NAND2_X1 U942 ( .A1(n872), .A2(G124), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U944 ( .A1(G136), .A2(n868), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U946 ( .A(KEYINPUT102), .B(n850), .ZN(n855) );
  NAND2_X1 U947 ( .A1(G100), .A2(n869), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G112), .A2(n873), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U950 ( .A(KEYINPUT103), .B(n853), .Z(n854) );
  NOR2_X1 U951 ( .A1(n855), .A2(n854), .ZN(G162) );
  NAND2_X1 U952 ( .A1(n868), .A2(G142), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT105), .B(n856), .Z(n858) );
  NAND2_X1 U954 ( .A1(n869), .A2(G106), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n859), .B(KEYINPUT45), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G118), .A2(n873), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U959 ( .A1(n872), .A2(G130), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT104), .B(n862), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n865), .B(n978), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n889) );
  NAND2_X1 U964 ( .A1(G139), .A2(n868), .ZN(n871) );
  NAND2_X1 U965 ( .A1(G103), .A2(n869), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n878) );
  NAND2_X1 U967 ( .A1(G127), .A2(n872), .ZN(n875) );
  NAND2_X1 U968 ( .A1(G115), .A2(n873), .ZN(n874) );
  NAND2_X1 U969 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U971 ( .A1(n878), .A2(n877), .ZN(n963) );
  XOR2_X1 U972 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n880) );
  XNOR2_X1 U973 ( .A(G162), .B(KEYINPUT107), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U975 ( .A(n881), .B(KEYINPUT106), .Z(n883) );
  XNOR2_X1 U976 ( .A(G164), .B(KEYINPUT48), .ZN(n882) );
  XNOR2_X1 U977 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U978 ( .A(n963), .B(n884), .ZN(n887) );
  XOR2_X1 U979 ( .A(G160), .B(n885), .Z(n886) );
  XNOR2_X1 U980 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U981 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U982 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U983 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U984 ( .A(n893), .B(G286), .ZN(n895) );
  XNOR2_X1 U985 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U986 ( .A(n930), .B(G171), .Z(n896) );
  XNOR2_X1 U987 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U988 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U989 ( .A(G2451), .B(G2430), .Z(n900) );
  XNOR2_X1 U990 ( .A(G2438), .B(G2443), .ZN(n899) );
  XNOR2_X1 U991 ( .A(n900), .B(n899), .ZN(n906) );
  XOR2_X1 U992 ( .A(G2435), .B(G2454), .Z(n902) );
  XNOR2_X1 U993 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U995 ( .A(G2446), .B(G2427), .Z(n903) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U997 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U998 ( .A1(G14), .A2(n907), .ZN(n913) );
  NAND2_X1 U999 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1002 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G108), .ZN(G238) );
  INV_X1 U1007 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1008 ( .A(G301), .B(G1961), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(G299), .B(G1956), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(n923) );
  XNOR2_X1 U1013 ( .A(G1971), .B(G303), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n929) );
  XNOR2_X1 U1016 ( .A(G1966), .B(G168), .ZN(n924) );
  XNOR2_X1 U1017 ( .A(n924), .B(KEYINPUT120), .ZN(n925) );
  NAND2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1019 ( .A(KEYINPUT57), .B(n927), .Z(n928) );
  NOR2_X1 U1020 ( .A1(n929), .A2(n928), .ZN(n935) );
  XNOR2_X1 U1021 ( .A(n930), .B(G1341), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(n931), .B(G1348), .ZN(n932) );
  NOR2_X1 U1023 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1024 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1025 ( .A(G16), .B(KEYINPUT56), .Z(n936) );
  XNOR2_X1 U1026 ( .A(KEYINPUT119), .B(n936), .ZN(n937) );
  NAND2_X1 U1027 ( .A1(n938), .A2(n937), .ZN(n1027) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n992) );
  XOR2_X1 U1029 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n953) );
  XNOR2_X1 U1030 ( .A(G1991), .B(G25), .ZN(n950) );
  XOR2_X1 U1031 ( .A(n939), .B(G27), .Z(n942) );
  XOR2_X1 U1032 ( .A(KEYINPUT116), .B(G32), .Z(n940) );
  XNOR2_X1 U1033 ( .A(G1996), .B(n940), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(G2072), .B(G33), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(n945), .B(KEYINPUT115), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(n948), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(n953), .B(n952), .ZN(n955) );
  XNOR2_X1 U1044 ( .A(G35), .B(G2090), .ZN(n954) );
  NOR2_X1 U1045 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1046 ( .A(G2084), .B(KEYINPUT54), .Z(n956) );
  XNOR2_X1 U1047 ( .A(G34), .B(n956), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(n992), .B(n959), .ZN(n961) );
  INV_X1 U1050 ( .A(G29), .ZN(n960) );
  NAND2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n962), .ZN(n1025) );
  XOR2_X1 U1053 ( .A(KEYINPUT52), .B(KEYINPUT114), .Z(n990) );
  XNOR2_X1 U1054 ( .A(G2072), .B(n963), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G164), .B(G2078), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n964), .B(KEYINPUT112), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(n967), .B(KEYINPUT113), .ZN(n968) );
  XOR2_X1 U1059 ( .A(KEYINPUT50), .B(n968), .Z(n986) );
  XOR2_X1 U1060 ( .A(G2090), .B(G162), .Z(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1062 ( .A(KEYINPUT51), .B(n971), .Z(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT110), .B(n972), .ZN(n974) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n983) );
  XOR2_X1 U1065 ( .A(G2084), .B(G160), .Z(n975) );
  NOR2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(n979), .B(KEYINPUT109), .ZN(n981) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(KEYINPUT111), .B(n984), .ZN(n985) );
  NOR2_X1 U1072 ( .A1(n986), .A2(n985), .ZN(n988) );
  NAND2_X1 U1073 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(n990), .B(n989), .ZN(n991) );
  NAND2_X1 U1075 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1076 ( .A1(n993), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1077 ( .A(KEYINPUT121), .B(G16), .ZN(n1021) );
  XOR2_X1 U1078 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n1004) );
  XNOR2_X1 U1079 ( .A(KEYINPUT59), .B(G1348), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(n994), .B(G4), .ZN(n1002) );
  XNOR2_X1 U1081 ( .A(G1956), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1082 ( .A(G1981), .B(G6), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n995), .B(KEYINPUT122), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G19), .B(G1341), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT123), .B(n998), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(n1004), .B(n1003), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G1961), .B(G5), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1018) );
  XOR2_X1 U1094 ( .A(G1986), .B(G24), .Z(n1014) );
  XOR2_X1 U1095 ( .A(G1976), .B(KEYINPUT125), .Z(n1009) );
  XNOR2_X1 U1096 ( .A(G23), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G22), .B(G1971), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(n1012), .B(KEYINPUT126), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(KEYINPUT127), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1108 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

