//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n585, new_n586, new_n589, new_n590,
    new_n592, new_n593, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1100,
    new_n1101;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n453), .B2(G2106), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(new_n464), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT69), .Z(new_n476));
  INV_X1    g051(.A(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n465), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n465), .A2(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n464), .A2(KEYINPUT71), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  AND4_X1   g073(.A1(KEYINPUT72), .A2(new_n490), .A3(new_n492), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n493), .A2(new_n497), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT71), .B1(new_n464), .B2(new_n488), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT72), .B1(new_n502), .B2(new_n490), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n499), .A2(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n511), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  XOR2_X1   g091(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n507), .A2(new_n522), .B1(new_n509), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(G168));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n507), .A2(new_n526), .B1(new_n509), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n513), .ZN(new_n530));
  OR3_X1    g105(.A1(new_n528), .A2(new_n530), .A3(KEYINPUT74), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT74), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n513), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT75), .B(G81), .Z(new_n536));
  NOR2_X1   g111(.A1(new_n507), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n509), .ZN(new_n538));
  AOI211_X1 g113(.A(new_n535), .B(new_n537), .C1(G43), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  NAND2_X1  g119(.A1(G78), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n506), .ZN(new_n546));
  INV_X1    g121(.A(G65), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n513), .B1(new_n548), .B2(KEYINPUT76), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n549), .B1(KEYINPUT76), .B2(new_n548), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OR3_X1    g126(.A1(new_n509), .A2(KEYINPUT9), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n509), .B2(new_n551), .ZN(new_n553));
  INV_X1    g128(.A(new_n507), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n552), .A2(new_n553), .B1(G91), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  INV_X1    g132(.A(G168), .ZN(G286));
  OAI21_X1  g133(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n559));
  INV_X1    g134(.A(G49), .ZN(new_n560));
  INV_X1    g135(.A(G87), .ZN(new_n561));
  OAI221_X1 g136(.A(new_n559), .B1(new_n509), .B2(new_n560), .C1(new_n561), .C2(new_n507), .ZN(G288));
  NAND2_X1  g137(.A1(G73), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G61), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n546), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n538), .B2(G48), .ZN(new_n566));
  INV_X1    g141(.A(G86), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(new_n507), .ZN(G305));
  XOR2_X1   g143(.A(KEYINPUT77), .B(G85), .Z(new_n569));
  INV_X1    g144(.A(G47), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n507), .A2(new_n569), .B1(new_n509), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n513), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(new_n554), .A2(G92), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT10), .Z(new_n577));
  NAND2_X1  g152(.A1(G79), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G66), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n546), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n538), .B2(G54), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  MUX2_X1   g157(.A(new_n582), .B(G301), .S(G868), .Z(G321));
  XOR2_X1   g158(.A(G321), .B(KEYINPUT78), .Z(G284));
  NAND2_X1  g159(.A1(G286), .A2(G868), .ZN(new_n585));
  INV_X1    g160(.A(G299), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(G868), .ZN(G297));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(G868), .ZN(G280));
  INV_X1    g163(.A(new_n582), .ZN(new_n589));
  INV_X1    g164(.A(G559), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(G860), .ZN(G148));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G868), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G868), .B2(new_n539), .ZN(G323));
  XNOR2_X1  g169(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n595));
  XNOR2_X1  g170(.A(G323), .B(new_n595), .ZN(G282));
  NAND2_X1  g171(.A1(new_n477), .A2(G135), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n474), .A2(G123), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n465), .A2(G111), .ZN(new_n599));
  OAI21_X1  g174(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT81), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(G2096), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(G2096), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n464), .A2(new_n462), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT80), .B(G2100), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n607), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n604), .A2(new_n605), .A3(new_n610), .ZN(G156));
  XNOR2_X1  g186(.A(G2427), .B(G2438), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2430), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT15), .B(G2435), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(KEYINPUT14), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(G1341), .B(G1348), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2443), .B(G2446), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n617), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(G2451), .B(G2454), .Z(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G14), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n621), .A2(new_n624), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(G401));
  XOR2_X1   g203(.A(G2072), .B(G2078), .Z(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT83), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT17), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2067), .B(G2678), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT84), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n635), .B(new_n637), .C1(new_n634), .C2(new_n630), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n632), .A3(new_n636), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT18), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n633), .A2(new_n636), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n640), .C1(new_n631), .C2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT85), .ZN(new_n643));
  XOR2_X1   g218(.A(G2096), .B(G2100), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(G227));
  XOR2_X1   g220(.A(G1971), .B(G1976), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT19), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1956), .B(G2474), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1961), .B(G1966), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT87), .Z(new_n652));
  NOR2_X1   g227(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  NOR3_X1   g231(.A1(new_n647), .A2(new_n650), .A3(new_n653), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n652), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1981), .B(G1986), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G229));
  INV_X1    g239(.A(G16), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G24), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n574), .B2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT89), .B(G1986), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n667), .B(new_n668), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n477), .A2(G131), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n474), .A2(G119), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n465), .A2(G107), .ZN(new_n672));
  OAI21_X1  g247(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n671), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  MUX2_X1   g249(.A(G25), .B(new_n674), .S(G29), .Z(new_n675));
  XOR2_X1   g250(.A(KEYINPUT35), .B(G1991), .Z(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT88), .Z(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(new_n677), .Z(new_n678));
  NAND2_X1  g253(.A1(G303), .A2(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n665), .A2(G22), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G1971), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n665), .A2(G6), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G305), .B2(G16), .ZN(new_n688));
  AOI211_X1 g263(.A(new_n683), .B(new_n684), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  OR2_X1    g265(.A1(G288), .A2(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g266(.A1(G288), .A2(KEYINPUT90), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n693), .B2(G16), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n689), .B(new_n696), .C1(new_n686), .C2(new_n688), .ZN(new_n697));
  AOI211_X1 g272(.A(new_n669), .B(new_n678), .C1(new_n697), .C2(KEYINPUT34), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(KEYINPUT34), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n698), .A2(new_n699), .B1(KEYINPUT91), .B2(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n701), .A2(KEYINPUT91), .A3(new_n700), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(KEYINPUT91), .B2(new_n700), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n539), .A2(new_n665), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n665), .B2(G19), .ZN(new_n705));
  INV_X1    g280(.A(G1341), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  OAI22_X1  g282(.A1(new_n705), .A2(new_n706), .B1(new_n603), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT30), .B(G28), .ZN(new_n710));
  OR2_X1    g285(.A1(KEYINPUT31), .A2(G11), .ZN(new_n711));
  NAND2_X1  g286(.A1(KEYINPUT31), .A2(G11), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n710), .A2(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n474), .A2(G129), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT94), .Z(new_n715));
  AND2_X1   g290(.A1(new_n462), .A2(G105), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT26), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n716), .B(new_n718), .C1(new_n477), .C2(G141), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(new_n707), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n707), .B2(G32), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n709), .B(new_n713), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n707), .B1(KEYINPUT24), .B2(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(KEYINPUT24), .B2(G34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n468), .A2(new_n471), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G29), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n708), .B(new_n725), .C1(new_n726), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n707), .A2(G26), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n474), .A2(G128), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n477), .A2(G140), .ZN(new_n735));
  OR2_X1    g310(.A1(G104), .A2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n736), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n733), .B1(new_n738), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2067), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n589), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G4), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1348), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n723), .B2(new_n724), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G162), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT29), .B(G2090), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n731), .A2(new_n745), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G286), .A2(new_n665), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT95), .B1(G16), .B2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT96), .B(G1966), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n757), .B(new_n758), .Z(new_n759));
  NOR2_X1   g334(.A1(new_n730), .A2(new_n726), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G5), .A2(G16), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G171), .B2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT97), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G1961), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G139), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n466), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(KEYINPUT92), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(KEYINPUT92), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n773), .A2(new_n774), .B1(new_n465), .B2(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G33), .B(new_n776), .S(G29), .Z(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G2072), .Z(new_n778));
  NAND4_X1  g353(.A1(new_n762), .A2(new_n766), .A3(new_n767), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n665), .A2(G20), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT23), .Z(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G299), .B2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1956), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n707), .A2(G27), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G164), .B2(new_n707), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2078), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n752), .A2(new_n779), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n702), .A2(new_n703), .A3(new_n787), .ZN(G150));
  INV_X1    g363(.A(G150), .ZN(G311));
  NAND2_X1  g364(.A1(new_n589), .A2(G559), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT38), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT98), .B(G93), .Z(new_n792));
  NOR2_X1   g367(.A1(new_n507), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(new_n513), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n793), .B(new_n795), .C1(G55), .C2(new_n538), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n539), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n539), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n791), .B(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT39), .ZN(new_n802));
  INV_X1    g377(.A(G860), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(KEYINPUT39), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n796), .A2(new_n803), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT37), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n807), .ZN(G145));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n776), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT99), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(new_n738), .ZN(new_n812));
  AOI22_X1  g387(.A1(G130), .A2(new_n474), .B1(new_n477), .B2(G142), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n465), .A2(G118), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n461), .B1(new_n814), .B2(KEYINPUT101), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT101), .B1(G106), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n815), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n607), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n812), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n502), .A2(new_n490), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n720), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n674), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n821), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n602), .B(G160), .ZN(new_n826));
  XNOR2_X1  g401(.A(G162), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT102), .B(G37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(G395));
  XOR2_X1   g407(.A(new_n592), .B(new_n799), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n589), .A2(G299), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n582), .A2(new_n586), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(KEYINPUT104), .A3(new_n835), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n582), .A2(new_n586), .A3(KEYINPUT104), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT41), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n834), .A2(new_n835), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n839), .B1(new_n844), .B2(new_n833), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n693), .B(G305), .ZN(new_n848));
  XNOR2_X1  g423(.A(G303), .B(new_n574), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n847), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G868), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(G868), .B2(new_n796), .ZN(G295));
  OAI21_X1  g429(.A(new_n853), .B1(G868), .B2(new_n796), .ZN(G331));
  OR2_X1    g430(.A1(new_n841), .A2(new_n842), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n836), .A2(new_n837), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n842), .ZN(new_n858));
  XNOR2_X1  g433(.A(G171), .B(G168), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n800), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n799), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n856), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT108), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n856), .A2(new_n858), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT107), .B1(new_n860), .B2(new_n800), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n863), .B2(KEYINPUT107), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n865), .B(new_n867), .C1(new_n857), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n851), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n838), .A2(new_n861), .A3(new_n862), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n850), .B(new_n873), .C1(new_n844), .C2(new_n869), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n874), .A2(new_n829), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT43), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n840), .A3(new_n843), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n850), .B1(new_n878), .B2(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n884), .A3(KEYINPUT44), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n872), .A2(new_n875), .A3(new_n882), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n879), .B2(new_n881), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n888), .A2(KEYINPUT109), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT109), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT110), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(KEYINPUT110), .B(new_n885), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(G397));
  NAND2_X1  g471(.A1(G160), .A2(G40), .ZN(new_n897));
  AOI21_X1  g472(.A(G1384), .B1(new_n502), .B2(new_n490), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT45), .ZN(new_n899));
  INV_X1    g474(.A(G1996), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n720), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n738), .B(new_n740), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n676), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n674), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n899), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(G290), .A2(G1986), .ZN(new_n907));
  NOR2_X1   g482(.A1(G290), .A2(G1986), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT111), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT54), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT53), .ZN(new_n913));
  INV_X1    g488(.A(G1384), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n499), .B2(new_n503), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n498), .A2(new_n492), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(new_n916), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(new_n897), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n913), .B1(new_n923), .B2(G2078), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(KEYINPUT50), .ZN(new_n925));
  XNOR2_X1  g500(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n897), .B1(new_n898), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G1961), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n468), .B(KEYINPUT122), .ZN(new_n930));
  INV_X1    g505(.A(G2078), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(KEYINPUT53), .A3(G40), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n930), .A2(new_n471), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n898), .A2(KEYINPUT45), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n933), .A2(new_n921), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n924), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n912), .B1(new_n936), .B2(G171), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT121), .ZN(new_n938));
  OAI211_X1 g513(.A(KEYINPUT45), .B(new_n914), .C1(new_n499), .C2(new_n503), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n897), .B1(new_n916), .B2(new_n920), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n931), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n913), .B1(new_n941), .B2(KEYINPUT120), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT120), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n939), .A2(new_n940), .A3(new_n943), .A4(new_n931), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n938), .B(new_n928), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(KEYINPUT53), .A3(new_n944), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT121), .B1(new_n947), .B2(new_n929), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n924), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n937), .B1(new_n949), .B2(G171), .ZN(new_n950));
  INV_X1    g525(.A(G8), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n939), .A2(new_n940), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n758), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n925), .A2(new_n726), .A3(new_n927), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT51), .B1(new_n955), .B2(KEYINPUT119), .ZN(new_n956));
  NAND2_X1  g531(.A1(G286), .A2(G8), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT118), .Z(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n955), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(KEYINPUT119), .A3(KEYINPUT51), .A4(new_n958), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n953), .A2(new_n954), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n963), .A2(new_n958), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT114), .B(G86), .Z(new_n966));
  OAI21_X1  g541(.A(new_n566), .B1(new_n507), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(G1981), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT113), .B(G1981), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n566), .B(new_n969), .C1(new_n567), .C2(new_n507), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT115), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI211_X1 g548(.A(KEYINPUT115), .B(KEYINPUT49), .C1(new_n968), .C2(new_n970), .ZN(new_n974));
  INV_X1    g549(.A(new_n897), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n898), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G8), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n973), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n977), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n691), .A2(G1976), .A3(new_n692), .ZN(new_n980));
  INV_X1    g555(.A(G1976), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(G288), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n979), .B2(new_n980), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n978), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n923), .A2(new_n682), .ZN(new_n987));
  INV_X1    g562(.A(G2090), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n925), .A2(new_n988), .A3(new_n927), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n951), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(G303), .A2(G8), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT55), .Z(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n915), .A2(KEYINPUT50), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n975), .B1(new_n898), .B2(new_n926), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n988), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n987), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n992), .B1(new_n999), .B2(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n994), .A2(new_n1000), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n950), .A2(new_n965), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n936), .A2(G171), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n924), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n947), .A2(new_n929), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n938), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n947), .A2(KEYINPUT121), .A3(new_n929), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1004), .B1(new_n1009), .B2(G301), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT123), .B1(new_n1010), .B2(new_n912), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1003), .B1(new_n949), .B2(G171), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT123), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT54), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1002), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT124), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT124), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(new_n1002), .C1(new_n1011), .C2(new_n1014), .ZN(new_n1018));
  INV_X1    g593(.A(new_n976), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT58), .B(G1341), .ZN(new_n1020));
  OAI22_X1  g595(.A1(new_n923), .A2(G1996), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n539), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT117), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT59), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n997), .A2(G1956), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n917), .A2(new_n922), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(G299), .B(KEYINPUT57), .Z(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT61), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1030), .B2(new_n1028), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1028), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(KEYINPUT61), .A3(new_n1029), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n925), .A2(new_n927), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n744), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1019), .A2(new_n740), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OR3_X1    g614(.A1(new_n1039), .A2(KEYINPUT60), .A3(new_n582), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n589), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n582), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT60), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1024), .A2(new_n1035), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1029), .B(KEYINPUT116), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1042), .B1(new_n1045), .B2(new_n1028), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1016), .A2(new_n1018), .A3(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n978), .A2(G1976), .A3(G288), .ZN(new_n1051));
  INV_X1    g626(.A(new_n970), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n979), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n986), .A2(new_n992), .A3(new_n990), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT63), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n994), .A2(new_n1000), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n955), .A2(G168), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n990), .A2(new_n992), .ZN(new_n1060));
  OR4_X1    g635(.A1(new_n1056), .A2(new_n994), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1055), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1009), .A2(G301), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1065), .B(new_n1001), .C1(KEYINPUT62), .C2(new_n965), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1063), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n911), .B1(new_n1050), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n899), .A2(new_n908), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT48), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1073), .A2(KEYINPUT48), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n906), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n674), .A2(new_n904), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n903), .A2(new_n1077), .B1(G2067), .B2(new_n738), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n899), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT47), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n899), .A2(new_n900), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1081), .A2(KEYINPUT46), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(KEYINPUT46), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n721), .A2(new_n902), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n899), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1076), .B(new_n1079), .C1(new_n1080), .C2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1086), .A2(new_n1080), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT126), .B1(new_n1072), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT126), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1070), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1062), .B1(new_n1093), .B2(new_n1068), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1015), .A2(KEYINPUT124), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(new_n1018), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1092), .B(new_n1089), .C1(new_n1096), .C2(new_n911), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1091), .A2(new_n1097), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g673(.A(G319), .B1(new_n626), .B2(new_n627), .ZN(new_n1100));
  NOR3_X1   g674(.A1(G229), .A2(G227), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g675(.A1(new_n830), .A2(new_n888), .A3(new_n1101), .ZN(G225));
  INV_X1    g676(.A(G225), .ZN(G308));
endmodule


