//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT77), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT77), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n188), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(G101), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n188), .A2(new_n191), .A3(new_n198), .A4(new_n192), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n199), .A2(KEYINPUT4), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n210), .A2(KEYINPUT64), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n211), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n203), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n194), .A2(G101), .A3(new_n196), .A4(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n201), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n221));
  OAI21_X1  g035(.A(G128), .B1(new_n221), .B2(KEYINPUT66), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n210), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n227), .A2(new_n207), .A3(new_n209), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n187), .A2(G107), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n190), .A2(G104), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n199), .A2(new_n233), .A3(KEYINPUT10), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n221), .A2(G128), .B1(new_n207), .B2(new_n209), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n199), .B(new_n233), .C1(new_n235), .C2(new_n228), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n237));
  AOI22_X1  g051(.A1(new_n230), .A2(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n243), .A3(new_n247), .A4(new_n244), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n220), .A2(new_n238), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G110), .B(G140), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(G227), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n251), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n220), .A2(new_n238), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n246), .A2(new_n248), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT80), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT80), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n260), .B(new_n249), .C1(new_n220), .C2(new_n238), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n199), .A2(new_n233), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n225), .A2(new_n229), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n249), .B1(new_n264), .B2(new_n236), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n250), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n254), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT81), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n262), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(G469), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G469), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n257), .A2(new_n258), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n260), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n257), .A2(KEYINPUT80), .A3(new_n258), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n255), .B1(new_n280), .B2(new_n250), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n250), .A2(new_n255), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n267), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n275), .B(new_n276), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n275), .A2(new_n276), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n274), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G214), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G113), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT2), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G113), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G116), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT68), .B(G119), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(G116), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(KEYINPUT68), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n303), .A3(G116), .ZN(new_n304));
  INV_X1    g118(.A(new_n296), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n294), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(KEYINPUT67), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n201), .A2(new_n309), .A3(new_n219), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n301), .A2(new_n303), .A3(new_n311), .A4(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G113), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n304), .A2(KEYINPUT5), .A3(new_n305), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n314), .A2(new_n315), .B1(new_n298), .B2(new_n294), .ZN(new_n316));
  INV_X1    g130(.A(new_n263), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G122), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n310), .A2(new_n320), .A3(new_n318), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n322), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n216), .A2(G125), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(G125), .B2(new_n230), .ZN(new_n328));
  INV_X1    g142(.A(G224), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G953), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT7), .B1(new_n329), .B2(G953), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n333), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n327), .B(new_n335), .C1(G125), .C2(new_n230), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n323), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n298), .A2(new_n294), .ZN(new_n339));
  INV_X1    g153(.A(new_n315), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n313), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n341), .B2(new_n263), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n317), .B1(new_n316), .B2(KEYINPUT83), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n339), .B(KEYINPUT83), .C1(new_n340), .C2(new_n313), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n263), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n338), .A3(new_n344), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n320), .B(KEYINPUT8), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(G902), .B1(new_n337), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n332), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G210), .B1(G237), .B2(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n332), .A2(new_n352), .A3(new_n354), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n289), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT9), .B(G234), .ZN(new_n359));
  OAI21_X1  g173(.A(G221), .B1(new_n359), .B2(G902), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n287), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  AOI211_X1 g176(.A(KEYINPUT85), .B(G143), .C1(new_n362), .C2(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(G214), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT85), .A2(G143), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT17), .B(G131), .C1(new_n363), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G125), .ZN(new_n369));
  INV_X1    g183(.A(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G140), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n371), .A3(KEYINPUT16), .ZN(new_n372));
  OR3_X1    g186(.A1(new_n370), .A2(KEYINPUT16), .A3(G140), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G146), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT75), .A4(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n373), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n206), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n367), .A2(new_n376), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G146), .B1(new_n372), .B2(new_n373), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n375), .B2(new_n374), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n384), .A2(KEYINPUT87), .A3(new_n377), .A4(new_n367), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n363), .A2(new_n366), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n247), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n364), .B(new_n365), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G131), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n382), .A2(new_n385), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n187), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n386), .B1(new_n395), .B2(new_n247), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(KEYINPUT18), .A3(G131), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n206), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n392), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n387), .A2(new_n389), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n369), .A2(new_n371), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT19), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n398), .A2(KEYINPUT19), .ZN(new_n407));
  AOI21_X1  g221(.A(G146), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n374), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n408), .A2(new_n409), .A3(new_n403), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n400), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n394), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(G475), .A2(G902), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n417), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n401), .B2(new_n415), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT88), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(KEYINPUT20), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT88), .B1(new_n416), .B2(new_n417), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n392), .A2(new_n394), .A3(new_n400), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n394), .B1(new_n392), .B2(new_n400), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n276), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n425), .A2(new_n426), .B1(new_n429), .B2(G475), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G217), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n359), .A2(new_n432), .A3(G953), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G116), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G122), .ZN(new_n436));
  AND2_X1   g250(.A1(KEYINPUT89), .A2(G122), .ZN(new_n437));
  NOR2_X1   g251(.A1(KEYINPUT89), .A2(G122), .ZN(new_n438));
  OAI21_X1  g252(.A(G116), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n439), .A2(KEYINPUT90), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n441), .B(G116), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n190), .B(new_n436), .C1(new_n440), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n208), .A2(G128), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n226), .A2(G143), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G134), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n446), .A3(new_n240), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n436), .B(KEYINPUT14), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n439), .A2(KEYINPUT90), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n442), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n452), .B1(new_n455), .B2(new_n190), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n436), .B(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n440), .B2(new_n443), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT92), .A3(G107), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n451), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G134), .B1(new_n445), .B2(KEYINPUT13), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT13), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(KEYINPUT91), .C1(new_n464), .C2(new_n447), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n447), .A2(new_n464), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n462), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n468), .A3(new_n449), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n454), .A2(new_n442), .B1(new_n435), .B2(G122), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n470), .A2(new_n190), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n471), .B2(new_n444), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n434), .B1(new_n461), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n444), .A2(new_n450), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n455), .A2(new_n452), .A3(new_n190), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT92), .B1(new_n459), .B2(G107), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n468), .A2(new_n449), .ZN(new_n478));
  INV_X1    g292(.A(new_n444), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n470), .A2(new_n190), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n465), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n481), .A3(new_n433), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n276), .ZN(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(G902), .B1(new_n473), .B2(new_n482), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(KEYINPUT15), .B2(new_n485), .ZN(new_n489));
  INV_X1    g303(.A(G952), .ZN(new_n490));
  AOI211_X1 g304(.A(G953), .B(new_n490), .C1(G234), .C2(G237), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n276), .B(new_n252), .C1(G234), .C2(G237), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT21), .B(G898), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT93), .B1(new_n431), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n424), .A4(new_n430), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n249), .B2(new_n216), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n504), .A2(new_n202), .B1(new_n203), .B2(new_n214), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n505), .A2(new_n258), .A3(KEYINPUT69), .A4(new_n213), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n242), .A2(KEYINPUT65), .A3(G134), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT65), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n240), .B2(G137), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n242), .A2(G134), .ZN(new_n511));
  OAI211_X1 g325(.A(G131), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n248), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n225), .B2(new_n229), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n299), .B(new_n294), .C1(new_n304), .C2(new_n305), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n307), .B1(new_n306), .B2(KEYINPUT67), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n300), .A2(KEYINPUT70), .A3(new_n308), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n507), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n521), .B1(new_n507), .B2(new_n515), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT28), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n525));
  INV_X1    g339(.A(new_n521), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n217), .A2(new_n258), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n515), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n525), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n514), .B1(new_n258), .B2(new_n217), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT28), .B1(new_n532), .B2(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n362), .A2(G210), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n535), .B(KEYINPUT27), .Z(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT26), .B(G101), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n524), .A2(new_n531), .A3(new_n534), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT72), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n533), .B(new_n530), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT72), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n524), .A4(new_n540), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n276), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n527), .A2(new_n515), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n514), .B1(new_n503), .B2(new_n506), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(new_n547), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n309), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n507), .A2(new_n521), .A3(new_n515), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n538), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n528), .A2(new_n309), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT28), .ZN(new_n557));
  INV_X1    g371(.A(new_n538), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n557), .A2(new_n531), .A3(new_n534), .A4(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n554), .A2(new_n539), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G472), .B1(new_n546), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT32), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n551), .A2(new_n552), .A3(new_n558), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n522), .B1(new_n550), .B2(new_n309), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(KEYINPUT31), .A3(new_n558), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n557), .A2(new_n531), .A3(new_n534), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n565), .A2(new_n567), .B1(new_n568), .B2(new_n538), .ZN(new_n569));
  NOR2_X1   g383(.A1(G472), .A2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n562), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n538), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n563), .A2(new_n564), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT31), .B1(new_n566), .B2(new_n558), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(KEYINPUT32), .A3(new_n570), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n561), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n432), .B1(G234), .B2(new_n276), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n579), .B(KEYINPUT73), .Z(new_n580));
  INV_X1    g394(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n297), .B2(G128), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n295), .A2(new_n226), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n297), .B2(new_n226), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n584), .B2(new_n581), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT76), .B(G110), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT24), .B(G110), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT74), .ZN(new_n588));
  OAI22_X1  g402(.A1(new_n585), .A2(new_n586), .B1(new_n588), .B2(new_n584), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n589), .B(new_n374), .C1(G146), .C2(new_n404), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n585), .A2(G110), .B1(new_n588), .B2(new_n584), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n384), .A2(new_n377), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n590), .A2(new_n593), .A3(new_n597), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n599), .A2(new_n276), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT25), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n580), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n276), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT25), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n599), .A2(new_n600), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n580), .A2(new_n276), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n361), .A2(new_n501), .A3(new_n578), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n576), .B2(new_n276), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n565), .A2(new_n567), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n571), .B1(new_n616), .B2(new_n573), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n606), .A2(new_n610), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n287), .A2(new_n360), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n483), .A2(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n473), .A2(new_n482), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(G478), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n485), .A2(new_n276), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n488), .B2(new_n485), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n431), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n357), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n354), .B1(new_n332), .B2(new_n352), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n495), .B(new_n288), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n619), .A2(new_n620), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n487), .A2(new_n489), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n424), .A2(new_n430), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n619), .A2(new_n620), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n615), .A2(new_n617), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n594), .A2(KEYINPUT94), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT94), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n590), .B2(new_n593), .ZN(new_n648));
  OR3_X1    g462(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n646), .B1(new_n644), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n609), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n606), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n361), .A2(new_n501), .A3(new_n643), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  AND3_X1   g470(.A1(new_n424), .A2(new_n430), .A3(new_n637), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n492), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n491), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n657), .A2(new_n658), .A3(new_n358), .A4(new_n662), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n578), .A2(new_n620), .A3(new_n663), .A4(new_n653), .ZN(new_n664));
  INV_X1    g478(.A(new_n662), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n638), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n358), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT95), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XNOR2_X1  g484(.A(new_n662), .B(KEYINPUT39), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n620), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n522), .A2(new_n523), .A3(new_n558), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(G902), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n566), .A2(new_n538), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n572), .A2(new_n577), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n356), .A2(new_n357), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n431), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n637), .A2(new_n288), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n682), .A2(new_n683), .A3(new_n653), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n673), .A2(new_n674), .A3(new_n679), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  AND3_X1   g501(.A1(new_n578), .A2(new_n620), .A3(new_n653), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n627), .B1(new_n424), .B2(new_n430), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n662), .ZN(new_n690));
  INV_X1    g504(.A(new_n358), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT96), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT97), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT96), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n689), .A2(new_n694), .A3(new_n358), .A4(new_n662), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n688), .A2(new_n692), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n578), .A2(new_n620), .A3(new_n695), .A4(new_n653), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n629), .A2(new_n665), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n694), .B1(new_n698), .B2(new_n358), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT97), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NAND3_X1  g516(.A1(new_n554), .A2(new_n559), .A3(new_n539), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n276), .A3(new_n545), .A4(new_n542), .ZN(new_n704));
  AOI22_X1  g518(.A1(KEYINPUT32), .A2(new_n617), .B1(new_n704), .B2(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n618), .B1(new_n705), .B2(new_n572), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n250), .B1(new_n259), .B2(new_n261), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n283), .B1(new_n707), .B2(new_n254), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n708), .B2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n284), .A2(new_n709), .A3(new_n360), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT98), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT98), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n284), .A2(new_n709), .A3(new_n712), .A4(new_n360), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(KEYINPUT99), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT99), .B1(new_n711), .B2(new_n713), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n706), .B(new_n633), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  OAI211_X1 g533(.A(new_n706), .B(new_n639), .C1(new_n715), .C2(new_n716), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND3_X1  g535(.A1(new_n711), .A2(new_n358), .A3(new_n713), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT100), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT100), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n711), .A2(new_n724), .A3(new_n358), .A4(new_n713), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n501), .A2(new_n578), .A3(new_n653), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  OAI21_X1  g543(.A(G472), .B1(new_n569), .B2(G902), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n570), .B(KEYINPUT101), .Z(new_n731));
  NOR2_X1   g545(.A1(new_n574), .A2(new_n575), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n558), .B1(new_n543), .B2(new_n524), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n611), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n358), .A2(new_n431), .A3(new_n637), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n494), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n715), .B2(new_n716), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NAND3_X1  g553(.A1(new_n730), .A2(new_n734), .A3(new_n653), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n730), .A2(new_n734), .A3(KEYINPUT102), .A4(new_n653), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n690), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n726), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n708), .A2(G469), .A3(G902), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n262), .A2(new_n269), .A3(G469), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n286), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n749), .A2(new_n286), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n284), .A2(KEYINPUT103), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n360), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n680), .A2(new_n289), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n360), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n751), .B2(new_n753), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n759), .B1(new_n761), .B2(KEYINPUT104), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n762), .A3(new_n706), .A4(new_n698), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n576), .A2(new_n570), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n562), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n572), .A2(KEYINPUT105), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n705), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n690), .A2(new_n764), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n770), .A2(new_n611), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n754), .A2(KEYINPUT104), .A3(new_n360), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n758), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n765), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  NAND4_X1  g593(.A1(new_n757), .A2(new_n762), .A3(new_n706), .A4(new_n666), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n271), .B2(new_n273), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  OAI21_X1  g597(.A(G469), .B1(new_n270), .B2(new_n783), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n782), .A2(KEYINPUT106), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT106), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n285), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n284), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n790), .B2(KEYINPUT107), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n792), .A3(new_n284), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n360), .A3(new_n671), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n431), .A2(new_n627), .ZN(new_n796));
  XOR2_X1   g610(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  OAI22_X1  g613(.A1(new_n431), .A2(new_n627), .B1(KEYINPUT108), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(KEYINPUT109), .A3(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n801), .B(new_n653), .C1(new_n617), .C2(new_n615), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT109), .B1(new_n798), .B2(new_n800), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n758), .A3(new_n806), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n795), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  NOR4_X1   g623(.A1(new_n578), .A2(new_n759), .A3(new_n690), .A4(new_n611), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT47), .B1(new_n794), .B2(new_n360), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n812), .B(new_n760), .C1(new_n791), .C2(new_n793), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n810), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  INV_X1    g629(.A(new_n811), .ZN(new_n816));
  INV_X1    g630(.A(new_n813), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n284), .A2(new_n709), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT110), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n760), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n661), .B1(new_n798), .B2(new_n800), .ZN(new_n822));
  INV_X1    g636(.A(new_n735), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n758), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT117), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n682), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n711), .A2(new_n713), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n824), .A2(new_n288), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT50), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n830), .A2(new_n759), .ZN(new_n833));
  INV_X1    g647(.A(new_n679), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n611), .A2(new_n833), .A3(new_n491), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n683), .A3(new_n627), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n742), .A2(new_n743), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n833), .A3(new_n822), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT51), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n828), .A2(new_n832), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n833), .A2(new_n770), .A3(new_n822), .A4(new_n611), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n835), .A2(new_n689), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(G952), .A3(new_n252), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n726), .B2(new_n825), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n832), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n821), .B2(new_n827), .ZN(new_n851));
  INV_X1    g665(.A(new_n839), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT51), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n654), .A2(new_n640), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n654), .A2(new_n640), .A3(KEYINPUT112), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n629), .B2(new_n632), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n689), .A2(KEYINPUT111), .A3(new_n358), .A4(new_n495), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n619), .A2(new_n860), .A3(new_n620), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n612), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n728), .A2(new_n717), .A3(new_n720), .A4(new_n738), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n837), .A2(new_n698), .A3(new_n757), .A4(new_n762), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n431), .A2(new_n637), .A3(new_n665), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n688), .A2(new_n758), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n778), .A2(new_n780), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n726), .A2(new_n744), .B1(new_n664), .B2(new_n668), .ZN(new_n874));
  INV_X1    g688(.A(new_n736), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n653), .A2(new_n760), .A3(new_n665), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n679), .A3(new_n876), .A4(new_n754), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n873), .A2(new_n701), .A3(new_n874), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n877), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n696), .B2(new_n700), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n873), .B1(new_n880), .B2(new_n874), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n872), .A2(new_n882), .A3(new_n883), .A4(KEYINPUT53), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n701), .A2(new_n874), .A3(new_n877), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT52), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n873), .A3(new_n874), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n870), .A2(new_n871), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT114), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n878), .B2(new_n881), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n886), .A2(KEYINPUT113), .A3(new_n887), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n895), .B2(new_n872), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT54), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n865), .A2(KEYINPUT116), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n578), .A2(new_n611), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT99), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n830), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n901), .B2(new_n714), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n902), .A2(new_n639), .B1(new_n726), .B2(new_n727), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n714), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n902), .A2(new_n633), .B1(new_n904), .B2(new_n737), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n889), .B1(new_n765), .B2(new_n777), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n898), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n866), .A2(new_n780), .A3(new_n868), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT115), .B1(new_n864), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n866), .A2(new_n780), .A3(new_n868), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n862), .A2(new_n612), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n856), .B2(new_n855), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n912), .A2(new_n913), .A3(new_n858), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n909), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n895), .A2(new_n917), .B1(new_n889), .B2(new_n888), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n897), .A2(new_n920), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n854), .A2(new_n921), .B1(G952), .B2(G953), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n819), .B(KEYINPUT49), .ZN(new_n923));
  NOR4_X1   g737(.A1(new_n829), .A2(new_n618), .A3(new_n289), .A4(new_n760), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n924), .A3(new_n834), .A4(new_n796), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(G75));
  NOR2_X1   g740(.A1(new_n252), .A2(G952), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT120), .Z(new_n928));
  NOR2_X1   g742(.A1(new_n918), .A2(new_n276), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(G210), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n324), .A2(new_n326), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(new_n331), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT56), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n928), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n929), .A2(G210), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT56), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n929), .A2(KEYINPUT119), .A3(G210), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n940), .B2(new_n933), .ZN(G51));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n918), .B2(new_n919), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n898), .A2(new_n907), .A3(new_n908), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n916), .A2(new_n911), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n894), .B2(new_n893), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT53), .B1(new_n872), .B2(new_n882), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT54), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n942), .B(KEYINPUT54), .C1(new_n947), .C2(new_n948), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n285), .B(KEYINPUT57), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n708), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n929), .A2(new_n785), .A3(new_n786), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n927), .B1(new_n955), .B2(new_n956), .ZN(G54));
  AND2_X1   g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n929), .A2(new_n416), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n416), .B1(new_n929), .B2(new_n958), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n927), .ZN(G60));
  XNOR2_X1  g775(.A(new_n625), .B(KEYINPUT59), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n897), .B2(new_n920), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n621), .A2(new_n623), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT122), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n928), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n962), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n951), .A2(new_n950), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(G63));
  XNOR2_X1  g783(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n432), .A2(new_n276), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n918), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n651), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n928), .B1(new_n976), .B2(new_n607), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n976), .A2(new_n607), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(new_n977), .A3(new_n928), .A4(new_n970), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n980), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n493), .B2(new_n329), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n864), .A2(new_n865), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n931), .B1(G898), .B2(new_n252), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  NAND2_X1  g802(.A1(new_n814), .A2(new_n808), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n758), .B1(new_n689), .B2(new_n657), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n899), .A2(new_n672), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n701), .A2(new_n874), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n686), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(KEYINPUT62), .A3(new_n686), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n992), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n990), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n252), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n406), .A2(new_n407), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n550), .B(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1000), .A2(KEYINPUT125), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n770), .A2(new_n611), .A3(new_n875), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n871), .B(new_n993), .C1(new_n795), .C2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(KEYINPUT126), .B1(new_n989), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1005), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1007), .A2(new_n1008), .A3(new_n808), .A4(new_n814), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1006), .A2(new_n252), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1002), .B1(G900), .B2(G953), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1013));
  AOI21_X1  g827(.A(G953), .B1(new_n990), .B2(new_n998), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1002), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1003), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n252), .B1(G227), .B2(G900), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1018), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1003), .A2(new_n1012), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(G72));
  XNOR2_X1  g836(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n985), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n999), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n927), .B1(new_n1027), .B2(new_n677), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n554), .A2(new_n563), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1025), .B(new_n1029), .C1(new_n891), .C2(new_n896), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1006), .A2(new_n985), .A3(new_n1009), .ZN(new_n1032));
  AOI211_X1 g846(.A(new_n558), .B(new_n553), .C1(new_n1032), .C2(new_n1025), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1031), .A2(new_n1033), .ZN(G57));
endmodule


