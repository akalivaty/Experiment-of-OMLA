//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1315,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1381, new_n1382;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT64), .ZN(new_n243));
  XOR2_X1   g0043(.A(G58), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  OR2_X1    g0049(.A1(KEYINPUT65), .A2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT65), .A2(G45), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n206), .A2(G274), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n256), .C2(new_n251), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n227), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT66), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n256), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(G1698), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n272), .B1(new_n228), .B2(new_n270), .C1(new_n273), .C2(new_n221), .ZN(new_n274));
  INV_X1    g0074(.A(new_n257), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n260), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G179), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n216), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT15), .B(G87), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n207), .A2(G33), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n281), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n280), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(G77), .B1(new_n207), .B2(G1), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n293), .A2(new_n294), .B1(G77), .B2(new_n290), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(new_n276), .B2(G169), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n278), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n277), .A2(G200), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n296), .B1(new_n276), .B2(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT67), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n207), .A2(G1), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n202), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n292), .A2(new_n306), .B1(new_n202), .B2(new_n291), .ZN(new_n307));
  INV_X1    g0107(.A(G150), .ZN(new_n308));
  INV_X1    g0108(.A(new_n284), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n282), .A2(new_n287), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(G20), .B2(new_n203), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(new_n281), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G226), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n255), .B1(new_n315), .B2(new_n259), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n317));
  INV_X1    g0117(.A(G223), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n317), .B1(new_n226), .B2(new_n270), .C1(new_n273), .C2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(new_n275), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n314), .B1(G200), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n321), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT68), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT10), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n322), .C1(new_n323), .C2(new_n321), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n321), .A2(G179), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n312), .B1(new_n320), .B2(G169), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n263), .A2(new_n268), .A3(G226), .A4(new_n271), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n263), .A2(new_n268), .A3(G232), .A4(G1698), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G97), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n275), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n255), .A2(KEYINPUT69), .B1(new_n259), .B2(new_n221), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n341), .B2(new_n344), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT14), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT14), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n351), .B(G169), .C1(new_n346), .C2(new_n347), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT71), .B1(new_n348), .B2(G179), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT71), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NOR4_X1   g0155(.A1(new_n346), .A2(new_n347), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n350), .B(new_n352), .C1(new_n353), .C2(new_n356), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n293), .A2(new_n220), .A3(new_n305), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT70), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n284), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n226), .B2(new_n287), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n361), .A2(new_n280), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(KEYINPUT11), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n291), .A2(new_n220), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT12), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(KEYINPUT11), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n341), .A2(new_n344), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT13), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n368), .B1(new_n374), .B2(new_n323), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n348), .A2(new_n325), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n255), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(G223), .A2(G1698), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n315), .B2(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n265), .A2(new_n267), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n383), .A2(new_n384), .B1(G33), .B2(G87), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n275), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n386), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n381), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G190), .ZN(new_n391));
  INV_X1    g0191(.A(G58), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n220), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n393), .B2(new_n201), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n284), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n261), .A2(new_n262), .A3(G20), .ZN(new_n398));
  XOR2_X1   g0198(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n397), .B(KEYINPUT16), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(KEYINPUT7), .ZN(new_n405));
  AOI21_X1  g0205(.A(G20), .B1(new_n263), .B2(new_n268), .ZN(new_n406));
  INV_X1    g0206(.A(new_n399), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n396), .B1(new_n408), .B2(G68), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n280), .B(new_n404), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n282), .A2(new_n305), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(new_n292), .B1(new_n291), .B2(new_n282), .ZN(new_n413));
  INV_X1    g0213(.A(new_n381), .ZN(new_n414));
  INV_X1    g0214(.A(new_n389), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n387), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G200), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n391), .A2(new_n411), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(G68), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n410), .B1(new_n420), .B2(new_n397), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n404), .A2(new_n280), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n413), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  OAI211_X1 g0224(.A(G179), .B(new_n414), .C1(new_n415), .C2(new_n387), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n390), .B2(new_n349), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n423), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n304), .A2(new_n336), .A3(new_n379), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n271), .A2(G244), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n265), .B2(new_n267), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT77), .B1(new_n434), .B2(KEYINPUT4), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT77), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT4), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n261), .A2(new_n262), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(new_n433), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G283), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n263), .A2(new_n268), .A3(G250), .A4(G1698), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n437), .A2(new_n227), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n263), .A2(new_n268), .A3(new_n271), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n275), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT5), .B(G41), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(new_n206), .A3(G45), .A4(G274), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n206), .B(G45), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n257), .ZN(new_n452));
  INV_X1    g0252(.A(G257), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n446), .A2(new_n355), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(G169), .B1(new_n446), .B2(new_n455), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g0258(.A(G97), .B(G107), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT6), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n460), .A2(new_n462), .A3(G107), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n464), .A2(new_n207), .B1(new_n226), .B2(new_n309), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n408), .A2(G107), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(KEYINPUT75), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT75), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n408), .A2(new_n468), .A3(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n281), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n281), .B(new_n290), .C1(G1), .C2(new_n256), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n290), .A2(new_n462), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n472), .A2(KEYINPUT76), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT76), .B1(new_n472), .B2(new_n473), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n458), .B(KEYINPUT78), .C1(new_n470), .C2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n384), .A2(new_n402), .A3(G20), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT66), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n207), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(new_n399), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT75), .B1(new_n483), .B2(new_n228), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n461), .A2(new_n463), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n469), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n476), .B1(new_n487), .B2(new_n280), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n446), .A2(new_n355), .A3(new_n455), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n437), .B1(new_n438), .B2(new_n433), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n491), .A2(new_n439), .A3(new_n442), .A4(new_n444), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n454), .B1(new_n492), .B2(new_n275), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n489), .B1(new_n493), .B2(G169), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n478), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n446), .A2(new_n455), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(G190), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n488), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n477), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n256), .A2(G1), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n291), .A2(new_n280), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n286), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n207), .B(G68), .C1(new_n261), .C2(new_n262), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n287), .B2(new_n462), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n207), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  NOR4_X1   g0311(.A1(new_n511), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G87), .A2(G97), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT79), .B1(new_n513), .B2(new_n228), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n281), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n503), .A2(new_n290), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n516), .A2(KEYINPUT80), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT80), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n222), .A2(new_n462), .A3(new_n228), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n511), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(KEYINPUT79), .A3(new_n228), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(new_n522), .B1(new_n207), .B2(new_n509), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n505), .A2(new_n507), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n280), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n517), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n519), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n504), .B1(new_n518), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n223), .B1(new_n206), .B2(G45), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n257), .A2(new_n529), .B1(new_n254), .B2(G45), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n256), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G238), .A2(G1698), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n227), .B2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n532), .B1(new_n534), .B2(new_n384), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n530), .B1(new_n535), .B2(new_n257), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n349), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G179), .B2(new_n536), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n528), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n471), .A2(new_n222), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n221), .A2(new_n271), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n227), .A2(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n261), .C2(new_n262), .ZN(new_n545));
  INV_X1    g0345(.A(new_n532), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n257), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n257), .A2(new_n529), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n254), .A2(G45), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(G200), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G190), .B(new_n530), .C1(new_n535), .C2(new_n257), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n542), .B(new_n553), .C1(new_n518), .C2(new_n527), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n222), .A2(KEYINPUT22), .A3(G20), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n263), .A2(new_n268), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n207), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT22), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT23), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n207), .B2(G107), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n228), .A2(KEYINPUT23), .A3(G20), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(new_n532), .B2(new_n207), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n560), .B1(new_n559), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n280), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT25), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n290), .A2(new_n568), .A3(G107), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n290), .B2(G107), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n502), .A2(G107), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n451), .A2(G264), .A3(new_n257), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G250), .A2(G1698), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n453), .B2(G1698), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n384), .B1(G33), .B2(G294), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n448), .B(new_n573), .C1(new_n576), .C2(new_n257), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n577), .A2(new_n323), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(G200), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n567), .A2(new_n572), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n540), .A2(new_n554), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n440), .B(new_n207), .C1(G33), .C2(new_n462), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n531), .A2(G20), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n280), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n290), .A2(G116), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n502), .B2(G116), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n269), .A2(G303), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n453), .A2(new_n271), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n229), .A2(G1698), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n261), .C2(new_n262), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(KEYINPUT81), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  INV_X1    g0396(.A(G303), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n263), .B2(new_n268), .ZN(new_n598));
  INV_X1    g0398(.A(new_n594), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n257), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n451), .A2(G270), .A3(new_n257), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G179), .A3(new_n448), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n590), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n448), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n349), .B1(new_n586), .B2(new_n588), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT21), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT21), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n607), .B(new_n610), .C1(new_n601), .C2(new_n605), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n567), .A2(new_n572), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n577), .A2(G179), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n349), .B2(new_n577), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(G200), .B1(new_n601), .B2(new_n605), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT81), .B1(new_n591), .B2(new_n594), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n598), .A2(new_n599), .A3(new_n596), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n275), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n605), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n617), .B(new_n590), .C1(new_n622), .C2(new_n323), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n581), .A2(new_n612), .A3(new_n616), .A4(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n432), .A2(new_n500), .A3(new_n624), .ZN(G372));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n427), .B2(new_n428), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n423), .A2(new_n426), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT18), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(KEYINPUT83), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n351), .B1(new_n374), .B2(G169), .ZN(new_n633));
  INV_X1    g0433(.A(new_n352), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n354), .B1(new_n374), .B2(new_n355), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n348), .A2(KEYINPUT71), .A3(G179), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n368), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n298), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n419), .A2(new_n378), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n632), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n334), .B1(new_n642), .B2(new_n331), .ZN(new_n643));
  INV_X1    g0443(.A(new_n604), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n610), .B1(new_n622), .B2(new_n607), .ZN(new_n645));
  INV_X1    g0445(.A(new_n611), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n616), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n581), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n540), .B1(new_n500), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT82), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n488), .A2(new_n494), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT80), .B1(new_n516), .B2(new_n517), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n525), .A2(new_n519), .A3(new_n526), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n541), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n528), .A2(new_n539), .B1(new_n654), .B2(new_n553), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n650), .B(KEYINPUT26), .C1(new_n651), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n487), .A2(new_n280), .ZN(new_n657));
  INV_X1    g0457(.A(new_n476), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n655), .A2(new_n659), .A3(new_n458), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT82), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT78), .B1(new_n659), .B2(new_n458), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n488), .A2(new_n494), .A3(new_n478), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT26), .B(new_n655), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n649), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n643), .B1(new_n432), .B2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n589), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n612), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n623), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(KEYINPUT84), .B(G330), .Z(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n613), .A2(new_n674), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n580), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n616), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n616), .A2(new_n674), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n612), .A2(new_n674), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(new_n685), .A3(new_n683), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n685), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n210), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n512), .A2(new_n514), .A3(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n214), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n700));
  XNOR2_X1  g0500(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n674), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n655), .B1(new_n664), .B2(new_n665), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT90), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n661), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n652), .A2(new_n653), .B1(new_n503), .B2(new_n502), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n554), .B1(new_n706), .B2(new_n538), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n477), .B2(new_n495), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT90), .B1(new_n708), .B2(KEYINPUT26), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n707), .A2(new_n488), .A3(new_n494), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT26), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n705), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n500), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n647), .A2(new_n581), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n477), .A2(new_n495), .A3(KEYINPUT91), .A4(new_n499), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n540), .B(KEYINPUT89), .Z(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT29), .B(new_n702), .C1(new_n712), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT92), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT88), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n723), .B(new_n724), .C1(new_n667), .C2(new_n674), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n650), .B1(new_n710), .B2(KEYINPUT26), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n660), .A2(KEYINPUT82), .A3(new_n661), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n666), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n540), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n477), .A2(new_n495), .A3(new_n499), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n715), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n674), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT88), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n725), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n705), .A2(new_n709), .A3(new_n711), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n717), .A3(new_n718), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(KEYINPUT92), .A3(KEYINPUT29), .A4(new_n702), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n722), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n573), .B1(new_n576), .B2(new_n257), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n739), .A2(new_n536), .A3(new_n603), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n620), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT87), .A3(KEYINPUT30), .A4(new_n493), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n493), .A2(KEYINPUT30), .A3(new_n620), .A4(new_n740), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT87), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n741), .B2(new_n496), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n577), .A2(new_n355), .A3(new_n536), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n622), .A2(new_n496), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT86), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n747), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(KEYINPUT86), .ZN(new_n756));
  OAI211_X1 g0556(.A(KEYINPUT31), .B(new_n674), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n655), .A2(new_n580), .A3(new_n623), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n647), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n730), .A2(new_n759), .A3(new_n702), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n752), .B1(new_n746), .B2(new_n743), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n702), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n757), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n679), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n738), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n701), .B1(new_n766), .B2(G1), .ZN(G364));
  NOR2_X1   g0567(.A1(new_n678), .A2(new_n679), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT93), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n207), .A2(G13), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n206), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n769), .B(new_n680), .C1(new_n695), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n216), .B1(G20), .B2(new_n349), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n207), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n355), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G77), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n323), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n207), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n462), .ZN(new_n783));
  NAND3_X1  g0583(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(new_n323), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n786), .A2(new_n220), .B1(new_n788), .B2(new_n202), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n783), .B(new_n789), .C1(new_n795), .C2(KEYINPUT32), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n207), .A2(new_n323), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n776), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n325), .A2(G179), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n392), .A2(new_n798), .B1(new_n800), .B2(new_n222), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n790), .A2(new_n799), .A3(new_n791), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n269), .B(new_n801), .C1(new_n803), .C2(G107), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n795), .A2(KEYINPUT32), .ZN(new_n805));
  AND4_X1   g0605(.A1(new_n780), .A2(new_n796), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n794), .A2(G329), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n800), .B(KEYINPUT97), .Z(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n809), .B2(new_n597), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n803), .A2(G283), .ZN(new_n811));
  INV_X1    g0611(.A(new_n777), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G311), .ZN(new_n813));
  INV_X1    g0613(.A(new_n798), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G322), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n811), .A2(new_n269), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G317), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n785), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G326), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n788), .B2(new_n821), .C1(new_n822), .C2(new_n782), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n810), .A2(new_n816), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n774), .B1(new_n806), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n695), .A2(new_n772), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT94), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n270), .A2(G355), .A3(new_n210), .ZN(new_n829));
  INV_X1    g0629(.A(G45), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n245), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n694), .A2(new_n384), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n250), .A2(new_n252), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n215), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n829), .B1(G116), .B2(new_n210), .C1(new_n831), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(G13), .A2(G33), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(G20), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n774), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n828), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n839), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n825), .B(new_n841), .C1(new_n678), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n773), .A2(new_n843), .ZN(G396));
  NOR3_X1   g0644(.A1(new_n278), .A2(new_n297), .A3(new_n674), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n300), .A2(new_n301), .B1(new_n296), .B2(new_n674), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n845), .B1(new_n847), .B2(new_n299), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n732), .B(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(new_n765), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n826), .B1(new_n849), .B2(new_n765), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n786), .A2(new_n308), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(G143), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n788), .A2(new_n854), .B1(new_n798), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n853), .B(new_n856), .C1(new_n779), .C2(G159), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n384), .B1(new_n392), .B2(new_n782), .C1(new_n809), .C2(new_n202), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n220), .A2(new_n802), .B1(new_n793), .B2(new_n861), .ZN(new_n862));
  NOR4_X1   g0662(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n783), .B1(G294), .B2(new_n814), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT98), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n809), .A2(new_n228), .B1(new_n531), .B2(new_n778), .ZN(new_n866));
  INV_X1    g0666(.A(G283), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n269), .B1(new_n786), .B2(new_n867), .C1(new_n597), .C2(new_n788), .ZN(new_n868));
  INV_X1    g0668(.A(G311), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n222), .A2(new_n802), .B1(new_n793), .B2(new_n869), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n865), .A2(new_n866), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n774), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n774), .A2(new_n837), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n828), .B1(new_n226), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n298), .A2(new_n702), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n298), .B2(new_n846), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n837), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n852), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(G384));
  OR2_X1    g0681(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(G116), .A3(new_n217), .A4(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT36), .Z(new_n885));
  OR3_X1    g0685(.A1(new_n214), .A2(new_n226), .A3(new_n393), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n202), .A2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n206), .B(G13), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n732), .A2(new_n848), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n877), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n438), .A2(new_n207), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n220), .B1(new_n892), .B2(KEYINPUT7), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n400), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n410), .B1(new_n894), .B2(new_n397), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n413), .B1(new_n422), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n672), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n419), .B2(new_n429), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n423), .A2(new_n897), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n628), .A2(new_n901), .A3(new_n418), .A4(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT100), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n896), .B1(new_n426), .B2(new_n897), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n902), .B1(new_n909), .B2(new_n418), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n900), .B(KEYINPUT38), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n628), .A2(new_n418), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n913), .A2(KEYINPUT100), .A3(new_n902), .A4(new_n901), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n910), .B1(new_n914), .B2(new_n905), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n912), .B1(new_n915), .B2(new_n899), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n674), .B1(new_n359), .B2(new_n367), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT99), .Z(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n639), .B2(new_n377), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n370), .A2(new_n378), .A3(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n891), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n632), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n672), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(KEYINPUT101), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n632), .A2(new_n419), .ZN(new_n929));
  INV_X1    g0729(.A(new_n901), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n913), .A2(new_n901), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT37), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n906), .B2(new_n907), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n915), .A2(new_n912), .A3(new_n899), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n370), .A2(new_n674), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT39), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n927), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n921), .A2(new_n922), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n890), .B2(new_n877), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n943), .A2(new_n917), .B1(new_n925), .B2(new_n672), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT101), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n722), .A2(new_n734), .A3(new_n431), .A4(new_n737), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n643), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n753), .A2(new_n747), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n760), .A2(new_n763), .A3(new_n951), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n923), .A2(new_n848), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n901), .B1(new_n632), .B2(new_n419), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n914), .A2(new_n905), .B1(new_n932), .B2(KEYINPUT37), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n912), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n911), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT40), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT40), .B1(new_n911), .B2(new_n916), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n953), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n431), .A2(new_n952), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n679), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n949), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n206), .B2(new_n770), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n949), .A2(new_n965), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n889), .B1(new_n967), .B2(new_n968), .ZN(G367));
  NAND2_X1  g0769(.A1(new_n659), .A2(new_n674), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n714), .A2(new_n716), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT102), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n973), .A2(new_n974), .B1(new_n651), .B2(new_n674), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n688), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n495), .B(new_n477), .C1(new_n975), .C2(new_n616), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n702), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n973), .A2(new_n974), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n651), .A2(new_n674), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n690), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT103), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n975), .A2(new_n690), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT42), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR4_X1   g0788(.A1(new_n975), .A2(KEYINPUT103), .A3(KEYINPUT42), .A4(new_n690), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n978), .B(new_n984), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n654), .A2(new_n702), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n729), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n707), .B2(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT104), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT103), .B1(new_n983), .B2(KEYINPUT42), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n986), .A2(new_n985), .A3(new_n987), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n977), .A2(new_n702), .B1(new_n983), .B2(KEYINPUT42), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT104), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n996), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n993), .B(new_n995), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n976), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n976), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1011), .B(new_n1008), .C1(new_n997), .C2(new_n1004), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n695), .B(KEYINPUT41), .Z(new_n1014));
  XOR2_X1   g0814(.A(new_n686), .B(new_n689), .Z(new_n1015));
  XNOR2_X1  g0815(.A(new_n680), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n766), .A2(KEYINPUT107), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT107), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n738), .A2(new_n765), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n1016), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n981), .C2(new_n692), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n1024));
  OR2_X1    g0824(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n975), .A2(new_n691), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(KEYINPUT45), .B1(new_n981), .B2(new_n692), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT45), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n975), .A2(new_n1028), .A3(new_n691), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1023), .B(new_n1026), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT106), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n687), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1029), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1028), .B1(new_n975), .B2(new_n691), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1035), .A2(new_n688), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1030), .A2(new_n687), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT106), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1022), .A2(new_n1032), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1014), .B1(new_n1039), .B2(new_n766), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1013), .B1(new_n1040), .B2(new_n772), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n832), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n840), .B1(new_n210), .B2(new_n286), .C1(new_n1042), .C2(new_n240), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n827), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT108), .Z(new_n1045));
  INV_X1    g0845(.A(new_n774), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n392), .A2(new_n800), .B1(new_n798), .B2(new_n308), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n269), .B(new_n1047), .C1(new_n794), .C2(G137), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n779), .A2(G50), .B1(G77), .B2(new_n803), .ZN(new_n1049));
  INV_X1    g0849(.A(G159), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n786), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n788), .A2(new_n855), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n782), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1051), .B(new_n1052), .C1(G68), .C2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1048), .A2(new_n1049), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n808), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT109), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n802), .A2(new_n462), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n779), .B2(G283), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n438), .B1(new_n798), .B2(new_n597), .C1(new_n822), .C2(new_n786), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G317), .B2(new_n794), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n800), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT46), .B1(new_n1062), .B2(G116), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n782), .A2(new_n228), .B1(new_n788), .B2(new_n869), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1059), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1055), .B1(new_n1057), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT47), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1046), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1045), .A2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT110), .Z(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n842), .B2(new_n993), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1041), .A2(new_n1073), .ZN(G387));
  NAND2_X1  g0874(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n696), .B1(new_n1020), .B2(new_n1016), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n842), .B1(new_n683), .B2(new_n685), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n832), .B1(new_n237), .B2(new_n833), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n270), .A2(new_n210), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n697), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n282), .A2(G50), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT50), .ZN(new_n1083));
  AOI21_X1  g0883(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n697), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1081), .A2(new_n1085), .B1(new_n228), .B2(new_n694), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n840), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n827), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n384), .B1(new_n794), .B2(G326), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n814), .A2(G317), .B1(G311), .B2(new_n785), .ZN(new_n1090));
  INV_X1    g0890(.A(G322), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n788), .C1(new_n778), .C2(new_n597), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1053), .A2(G283), .B1(new_n1062), .B2(G294), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT49), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1089), .B1(new_n531), .B2(new_n802), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n782), .A2(new_n286), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n283), .B2(new_n785), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1050), .B2(new_n788), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n438), .B1(new_n812), .B2(G68), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1062), .A2(G77), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n202), .C2(new_n798), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n1058), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n308), .B2(new_n793), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1099), .A2(new_n1101), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1078), .B(new_n1088), .C1(new_n1110), .C2(new_n774), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1016), .B2(new_n771), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1077), .A2(new_n1114), .ZN(G393));
  NAND2_X1  g0915(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1075), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1038), .A2(new_n1032), .A3(new_n1036), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n695), .B(new_n1117), .C1(new_n1118), .C2(new_n1075), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1116), .A2(new_n771), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n975), .A2(new_n839), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT111), .Z(new_n1122));
  AND2_X1   g0922(.A1(new_n832), .A2(new_n248), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n840), .B1(new_n462), .B2(new_n210), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n788), .A2(new_n308), .B1(new_n798), .B2(new_n1050), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT51), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n384), .B1(new_n800), .B2(new_n220), .C1(new_n202), .C2(new_n786), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n782), .A2(new_n226), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n222), .A2(new_n802), .B1(new_n793), .B2(new_n855), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n283), .B2(new_n779), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n228), .A2(new_n802), .B1(new_n793), .B2(new_n1091), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n269), .B1(new_n867), .B2(new_n800), .C1(new_n822), .C2(new_n777), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n782), .A2(new_n531), .B1(new_n786), .B2(new_n597), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n788), .A2(new_n817), .B1(new_n798), .B2(new_n869), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT52), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1131), .A2(new_n1133), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n827), .B1(new_n1123), .B2(new_n1124), .C1(new_n1140), .C2(new_n1046), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1122), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1120), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n1143), .ZN(G390));
  INV_X1    g0944(.A(KEYINPUT112), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n938), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n957), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n717), .A2(new_n718), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n674), .B1(new_n1149), .B2(new_n735), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n847), .A2(new_n299), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n845), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1145), .B(new_n1148), .C1(new_n1152), .C2(new_n942), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n702), .B(new_n1151), .C1(new_n712), .C2(new_n719), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n942), .B1(new_n1154), .B2(new_n877), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT112), .B1(new_n1155), .B2(new_n1147), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n674), .B(new_n878), .C1(new_n728), .C2(new_n731), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n923), .B1(new_n1158), .B2(new_n845), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1159), .A2(new_n1146), .B1(new_n937), .B2(new_n939), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n764), .A2(new_n923), .A3(new_n679), .A4(new_n848), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1160), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n952), .A2(G330), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n848), .A3(new_n923), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1163), .B(new_n772), .C1(new_n1164), .C2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1130), .B1(G116), .B2(new_n814), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT114), .Z(new_n1169));
  OAI221_X1 g0969(.A(new_n269), .B1(new_n786), .B2(new_n228), .C1(new_n867), .C2(new_n788), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n778), .A2(new_n462), .B1(new_n220), .B2(new_n802), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n809), .A2(new_n222), .B1(new_n822), .B2(new_n793), .ZN(new_n1172));
  OR4_X1    g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n782), .A2(new_n1050), .B1(new_n786), .B2(new_n854), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n269), .B(new_n1174), .C1(G132), .C2(new_n814), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n779), .A2(new_n1177), .B1(G50), .B2(new_n803), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n794), .A2(G125), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n787), .A2(G128), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n800), .A2(new_n308), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT53), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1182), .B2(new_n1181), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1175), .A2(new_n1178), .A3(new_n1179), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1046), .B1(new_n1173), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n828), .B(new_n1186), .C1(new_n282), .C2(new_n874), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n937), .A2(new_n939), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n838), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1167), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n942), .B1(new_n765), .B2(new_n878), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1166), .A2(new_n1192), .B1(new_n877), .B2(new_n890), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n763), .A2(new_n951), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n624), .A2(new_n500), .A3(new_n674), .ZN(new_n1195));
  OAI211_X1 g0995(.A(G330), .B(new_n848), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n942), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1197), .A2(new_n1162), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1152), .A2(new_n1198), .A3(KEYINPUT113), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1154), .A2(new_n877), .A3(new_n1197), .A4(new_n1162), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT113), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1193), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n431), .A2(new_n1165), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n947), .A2(new_n643), .A3(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n696), .B1(new_n1191), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1163), .B(new_n1206), .C1(new_n1164), .C2(new_n1166), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1190), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(G378));
  NAND3_X1  g1011(.A1(new_n1106), .A2(new_n251), .A3(new_n438), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1212), .A2(KEYINPUT115), .B1(new_n803), .B2(G58), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(KEYINPUT115), .B2(new_n1212), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n812), .A2(new_n503), .B1(G97), .B2(new_n785), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT116), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(KEYINPUT116), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT117), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n782), .A2(new_n220), .B1(new_n788), .B2(new_n531), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1217), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1218), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n228), .B2(new_n798), .C1(new_n867), .C2(new_n793), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1214), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n782), .A2(new_n308), .B1(new_n786), .B2(new_n861), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G125), .B2(new_n787), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1177), .A2(new_n1062), .B1(new_n814), .B2(G128), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n854), .C2(new_n777), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT59), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G33), .A2(G41), .ZN(new_n1230));
  INV_X1    g1030(.A(G124), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1230), .B1(new_n802), .B2(new_n1050), .C1(new_n1231), .C2(new_n793), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT118), .Z(new_n1233));
  OAI21_X1  g1033(.A(new_n1224), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1230), .A2(G50), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n384), .B2(G41), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1223), .B2(KEYINPUT58), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n774), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n772), .B(new_n695), .C1(new_n202), .C2(new_n874), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT119), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1242));
  NAND2_X1  g1042(.A1(new_n336), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n312), .A2(new_n897), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT120), .Z(new_n1245));
  INV_X1    g1045(.A(new_n1242), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n331), .A2(new_n335), .A3(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1243), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1241), .B1(new_n1251), .B2(new_n837), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT121), .Z(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n962), .B2(G330), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n958), .A2(KEYINPUT40), .B1(new_n953), .B2(new_n960), .ZN(new_n1255));
  INV_X1    g1055(.A(G330), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1255), .A2(new_n1250), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n927), .A2(new_n940), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n944), .A2(KEYINPUT101), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1254), .A2(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n962), .A2(G330), .A3(new_n1251), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1250), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n941), .A2(new_n945), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1253), .B1(new_n1265), .B2(new_n772), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT57), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1205), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1209), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n695), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT57), .B1(new_n1270), .B2(new_n1265), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1266), .B1(new_n1272), .B2(new_n1273), .ZN(G375));
  AND3_X1   g1074(.A1(new_n1203), .A2(KEYINPUT122), .A3(new_n1205), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT122), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1014), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1207), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n942), .A2(new_n837), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1102), .B1(G283), .B2(new_n814), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT123), .Z(new_n1282));
  OAI221_X1 g1082(.A(new_n269), .B1(new_n786), .B2(new_n531), .C1(new_n822), .C2(new_n788), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n778), .A2(new_n228), .B1(new_n226), .B2(new_n802), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n809), .A2(new_n462), .B1(new_n597), .B2(new_n793), .ZN(new_n1285));
  OR4_X1    g1085(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n808), .A2(G159), .B1(G128), .B2(new_n794), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n782), .A2(new_n202), .B1(new_n788), .B2(new_n861), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n785), .B2(new_n1177), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n384), .B1(new_n777), .B2(new_n308), .C1(new_n854), .C2(new_n798), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(G58), .B2(new_n803), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1046), .B1(new_n1286), .B2(new_n1292), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n828), .B(new_n1293), .C1(new_n220), .C2(new_n874), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1280), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1203), .B2(new_n771), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1279), .A2(new_n1297), .ZN(G381));
  AOI211_X1 g1098(.A(G396), .B(new_n1113), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n880), .ZN(new_n1300));
  OR3_X1    g1100(.A1(G390), .A2(G381), .A3(new_n1300), .ZN(new_n1301));
  OR3_X1    g1101(.A1(G387), .A2(new_n1301), .A3(KEYINPUT124), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1253), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1264), .B2(new_n771), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1166), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1162), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n1160), .B(new_n1306), .C1(new_n1153), .C2(new_n1156), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1205), .B1(new_n1308), .B2(new_n1206), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1267), .B1(new_n1309), .B2(new_n1264), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n696), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1304), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT124), .B1(G387), .B2(new_n1301), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1302), .A2(new_n1210), .A3(new_n1312), .A4(new_n1313), .ZN(G407));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1210), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G407), .B(G213), .C1(G343), .C2(new_n1315), .ZN(G409));
  AOI22_X1  g1116(.A1(new_n1077), .A2(new_n1114), .B1(new_n843), .B2(new_n773), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1317), .A2(new_n1299), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G390), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1119), .B(new_n1143), .C1(new_n1317), .C2(new_n1299), .ZN(new_n1320));
  AND4_X1   g1120(.A1(new_n1041), .A2(new_n1319), .A3(new_n1073), .A4(new_n1320), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1041), .A2(new_n1073), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1260), .A2(new_n1263), .A3(new_n1278), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT125), .B1(new_n1309), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1325), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1270), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1326), .A2(new_n1210), .A3(new_n1266), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n673), .A2(G213), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1330), .B(new_n1331), .C1(new_n1312), .C2(new_n1210), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1193), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1205), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT122), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1203), .A2(KEYINPUT122), .A3(new_n1205), .ZN(new_n1338));
  OAI21_X1  g1138(.A(KEYINPUT60), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1203), .A2(KEYINPUT60), .A3(new_n1205), .ZN(new_n1341));
  AND2_X1   g1141(.A1(new_n1341), .A2(new_n695), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G384), .B1(new_n1343), .B2(new_n1297), .ZN(new_n1344));
  AOI211_X1 g1144(.A(new_n880), .B(new_n1296), .C1(new_n1340), .C2(new_n1342), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(KEYINPUT62), .B1(new_n1332), .B2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1329), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1328), .B1(new_n1270), .B2(new_n1327), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1190), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1352), .A2(new_n1266), .A3(new_n1353), .ZN(new_n1354));
  AOI22_X1  g1154(.A1(new_n1351), .A2(new_n1354), .B1(G213), .B2(new_n673), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G375), .A2(G378), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT62), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1355), .A2(new_n1356), .A3(new_n1357), .A4(new_n1346), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1341), .A2(new_n695), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1359), .B1(new_n1277), .B2(new_n1339), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n880), .B1(new_n1360), .B2(new_n1296), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1343), .A2(G384), .A3(new_n1297), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n673), .A2(G213), .A3(G2897), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1363), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1365), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1366));
  AND2_X1   g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(KEYINPUT61), .B1(new_n1332), .B2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT127), .ZN(new_n1369));
  OAI211_X1 g1169(.A(new_n1348), .B(new_n1358), .C1(new_n1368), .C2(new_n1369), .ZN(new_n1370));
  AOI211_X1 g1170(.A(KEYINPUT127), .B(KEYINPUT61), .C1(new_n1332), .C2(new_n1367), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1324), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1355), .A2(new_n1356), .A3(KEYINPUT63), .A4(new_n1346), .ZN(new_n1373));
  AND2_X1   g1173(.A1(new_n1323), .A2(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1355), .A2(new_n1356), .A3(new_n1346), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT63), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1375), .A2(KEYINPUT126), .A3(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(KEYINPUT126), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1378));
  OAI211_X1 g1178(.A(new_n1374), .B(new_n1368), .C1(new_n1377), .C2(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1372), .A2(new_n1379), .ZN(G405));
  NAND2_X1  g1180(.A1(new_n1356), .A2(new_n1315), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1381), .B(new_n1346), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(new_n1382), .B(new_n1323), .ZN(G402));
endmodule


