//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1316, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT65), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n211), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n212), .B2(new_n218), .ZN(new_n220));
  INV_X1    g0020(.A(G1), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT66), .Z(new_n227));
  INV_X1    g0027(.A(new_n202), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n222), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n224), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n233), .B(new_n236), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n227), .A2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n231), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT68), .B1(new_n258), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(new_n222), .A3(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G150), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT69), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n261), .ZN(new_n266));
  OAI211_X1 g0066(.A(KEYINPUT69), .B(new_n264), .C1(new_n266), .C2(new_n256), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n203), .A2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n255), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n221), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n255), .ZN(new_n273));
  INV_X1    g0073(.A(G50), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n221), .B2(G20), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n273), .A2(new_n275), .B1(new_n274), .B2(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G169), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n221), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G77), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  OAI211_X1 g0094(.A(G222), .B(new_n294), .C1(new_n290), .C2(new_n291), .ZN(new_n295));
  OAI211_X1 g0095(.A(G223), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n284), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n293), .A2(KEYINPUT67), .A3(new_n295), .A4(new_n296), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n289), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n278), .B1(new_n279), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n273), .ZN(new_n307));
  OAI21_X1  g0107(.A(G77), .B1(new_n222), .B2(G1), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n307), .A2(new_n308), .B1(G77), .B2(new_n271), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n257), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n222), .A2(G33), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n309), .B1(new_n313), .B2(new_n255), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n285), .B1(new_n217), .B2(new_n288), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n258), .ZN(new_n318));
  NAND2_X1  g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n294), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(G238), .B1(new_n292), .B2(G107), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n319), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(G232), .A3(new_n294), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n284), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n304), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n315), .B(new_n327), .C1(G169), .C2(new_n326), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(G190), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n314), .C1(new_n330), .C2(new_n326), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT9), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n270), .A2(new_n333), .A3(new_n276), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n333), .B1(new_n270), .B2(new_n276), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n299), .A2(new_n300), .ZN(new_n338));
  INV_X1    g0138(.A(new_n289), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G190), .A3(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n340), .B(KEYINPUT70), .C1(new_n330), .C2(new_n301), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT10), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n301), .A2(new_n330), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n277), .A2(KEYINPUT9), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n334), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n306), .B(new_n332), .C1(new_n342), .C2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n284), .A2(G232), .A3(new_n287), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n285), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n354));
  OR2_X1    g0154(.A1(G223), .A2(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n286), .A2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(new_n356), .C1(new_n290), .C2(new_n291), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n325), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT75), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n285), .A2(new_n352), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n354), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT76), .ZN(new_n364));
  AOI22_X1  g0164(.A1(KEYINPUT75), .A2(new_n353), .B1(new_n359), .B2(new_n325), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT76), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n362), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n363), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n279), .B1(new_n304), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n322), .B2(G20), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n214), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G58), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n214), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n202), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n263), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n371), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n292), .B2(new_n222), .ZN(new_n382));
  NOR4_X1   g0182(.A1(new_n290), .A2(new_n291), .A3(new_n372), .A4(G20), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n380), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n255), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n256), .B1(new_n221), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n273), .B1(new_n272), .B2(new_n256), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n351), .B1(new_n370), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n363), .A2(KEYINPUT76), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n366), .B1(new_n365), .B2(new_n362), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n279), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n369), .A2(new_n304), .ZN(new_n395));
  AND4_X1   g0195(.A1(new_n351), .A2(new_n394), .A3(new_n390), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n389), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n254), .A2(new_n231), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n384), .A2(new_n385), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n371), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(new_n386), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n403));
  AOI21_X1  g0203(.A(G200), .B1(new_n364), .B2(new_n367), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n363), .A2(G190), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n402), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n330), .B1(new_n392), .B2(new_n393), .ZN(new_n407));
  INV_X1    g0207(.A(new_n405), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n390), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n397), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n350), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT12), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n272), .B2(new_n214), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n222), .B2(G1), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n415), .A2(new_n416), .B1(new_n307), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n214), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n266), .B2(new_n216), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n420), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT11), .B1(new_n420), .B2(new_n255), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n285), .B1(new_n215), .B2(new_n288), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  OAI211_X1 g0226(.A(G226), .B(new_n294), .C1(new_n290), .C2(new_n291), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT71), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n322), .A2(new_n430), .A3(G232), .A4(G1698), .ZN(new_n431));
  OAI211_X1 g0231(.A(G232), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT71), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n429), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n425), .B(new_n426), .C1(new_n434), .C2(new_n284), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT73), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n427), .A2(new_n428), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n430), .B1(new_n320), .B2(G232), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n432), .A2(KEYINPUT71), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n325), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT73), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n426), .A4(new_n425), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n426), .B1(new_n441), .B2(new_n425), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n304), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n433), .A2(new_n431), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n284), .B1(new_n447), .B2(new_n437), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT13), .B1(new_n448), .B2(new_n424), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n435), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G169), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n444), .A2(new_n446), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT14), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n453), .A3(G169), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n423), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n448), .A2(KEYINPUT13), .A3(new_n424), .ZN(new_n456));
  OAI21_X1  g0256(.A(G200), .B1(new_n445), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT72), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT72), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(new_n459), .A3(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT74), .ZN(new_n462));
  INV_X1    g0262(.A(new_n423), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n449), .A2(G190), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n444), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n459), .B1(new_n450), .B2(G200), .ZN(new_n468));
  AOI211_X1 g0268(.A(KEYINPUT72), .B(new_n330), .C1(new_n449), .C2(new_n435), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n436), .A2(new_n443), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n423), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT74), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n455), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n413), .A2(new_n474), .A3(KEYINPUT78), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT78), .B1(new_n413), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT88), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n222), .B(G87), .C1(new_n290), .C2(new_n291), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n322), .A2(new_n481), .A3(new_n222), .A4(G87), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G116), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT85), .B1(new_n484), .B2(G20), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT85), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(new_n222), .A3(G33), .A4(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT23), .ZN(new_n489));
  INV_X1    g0289(.A(G107), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(G20), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n222), .A2(G107), .B1(KEYINPUT86), .B2(KEYINPUT23), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n488), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT24), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n491), .B1(new_n493), .B2(new_n492), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n485), .B2(new_n487), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n480), .A2(new_n482), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n399), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT25), .ZN(new_n502));
  AOI211_X1 g0302(.A(G107), .B(new_n271), .C1(KEYINPUT87), .C2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(KEYINPUT87), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n221), .A2(G33), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n399), .A2(new_n271), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n478), .B1(new_n501), .B2(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n499), .B1(new_n497), .B2(new_n498), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n255), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n505), .A2(new_n506), .B1(G107), .B2(new_n510), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(KEYINPUT88), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G257), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n519));
  OAI211_X1 g0319(.A(G250), .B(new_n294), .C1(new_n290), .C2(new_n291), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G294), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n325), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n221), .B(G45), .C1(new_n280), .C2(KEYINPUT5), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT5), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G41), .ZN(new_n526));
  OAI211_X1 g0326(.A(G264), .B(new_n284), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n525), .B2(G41), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n280), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n281), .A2(G1), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(G41), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n284), .A2(G274), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n523), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G179), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n279), .B2(new_n536), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n513), .A2(new_n518), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT89), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n513), .A2(KEYINPUT89), .A3(new_n518), .A4(new_n538), .ZN(new_n542));
  INV_X1    g0342(.A(new_n527), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n325), .B2(new_n522), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n535), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n536), .A2(G190), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n516), .A2(new_n546), .A3(new_n547), .A4(new_n517), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n541), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G264), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n550));
  OAI211_X1 g0350(.A(G257), .B(new_n294), .C1(new_n290), .C2(new_n291), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n318), .A2(G303), .A3(new_n319), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n325), .ZN(new_n554));
  OAI211_X1 g0354(.A(G270), .B(new_n284), .C1(new_n524), .C2(new_n526), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n535), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n273), .A2(G116), .A3(new_n508), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n272), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n254), .A2(new_n231), .B1(G20), .B2(new_n558), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G283), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n222), .C1(G33), .C2(new_n209), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(KEYINPUT20), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT20), .B1(new_n560), .B2(new_n562), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n557), .B(new_n559), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n556), .A2(new_n566), .A3(G169), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n566), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n554), .A2(G190), .A3(new_n535), .A4(new_n555), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n555), .B1(new_n534), .B2(new_n533), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n325), .B2(new_n553), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n570), .B(new_n571), .C1(new_n573), .C2(new_n330), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(G179), .A3(new_n566), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n556), .A2(new_n566), .A3(KEYINPUT21), .A4(G169), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n569), .A2(new_n574), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n222), .B1(new_n428), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n207), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n222), .B(G68), .C1(new_n290), .C2(new_n291), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n578), .B1(new_n311), .B2(new_n209), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT83), .A4(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n255), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n312), .A2(new_n272), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n312), .B(KEYINPUT84), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n510), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n594));
  OAI211_X1 g0394(.A(G238), .B(new_n294), .C1(new_n290), .C2(new_n291), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n484), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n325), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n208), .B1(new_n281), .B2(G1), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n284), .A2(new_n598), .ZN(new_n599));
  OR3_X1    g0399(.A1(new_n281), .A2(G1), .A3(G274), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n279), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n596), .A2(new_n325), .B1(new_n600), .B2(new_n599), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n304), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n593), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n399), .B1(new_n585), .B2(new_n586), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n588), .B1(new_n272), .B2(new_n312), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n602), .A2(G200), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(G190), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n510), .A2(G87), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n608), .A2(new_n609), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n577), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(KEYINPUT79), .B(G107), .C1(new_n382), .C2(new_n383), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n490), .A2(KEYINPUT6), .A3(G97), .ZN(new_n616));
  AND2_X1   g0416(.A1(G97), .A2(G107), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(new_n580), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n618), .B2(KEYINPUT6), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n373), .A2(new_n374), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT79), .B1(new_n622), .B2(G107), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n255), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n284), .B1(new_n524), .B2(new_n526), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n625), .A2(new_n210), .B1(new_n533), .B2(new_n534), .ZN(new_n626));
  OAI211_X1 g0426(.A(G244), .B(new_n294), .C1(new_n290), .C2(new_n291), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT4), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n322), .A2(KEYINPUT4), .A3(G244), .A4(new_n294), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n322), .A2(G250), .A3(G1698), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n561), .A4(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n626), .B1(new_n632), .B2(new_n325), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G190), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n509), .A2(G97), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n271), .A2(new_n209), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT80), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT80), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n639), .A3(new_n636), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n624), .A2(new_n634), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n632), .A2(new_n325), .ZN(new_n643));
  INV_X1    g0443(.A(new_n626), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT82), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(G200), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT82), .B1(new_n633), .B2(new_n330), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI211_X1 g0449(.A(G179), .B(new_n626), .C1(new_n325), .C2(new_n632), .ZN(new_n650));
  AOI21_X1  g0450(.A(G169), .B1(new_n643), .B2(new_n644), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n624), .A2(new_n641), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n642), .A2(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n614), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n477), .A2(new_n549), .A3(new_n655), .ZN(G372));
  NAND2_X1  g0456(.A1(new_n473), .A2(new_n467), .ZN(new_n657));
  INV_X1    g0457(.A(new_n328), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n455), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n411), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n397), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n342), .B2(new_n349), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT10), .B1(new_n337), .B2(new_n341), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n346), .A2(new_n348), .A3(new_n343), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT92), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n661), .A2(new_n667), .B1(new_n305), .B2(new_n303), .ZN(new_n668));
  INV_X1    g0468(.A(new_n606), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(G190), .B2(new_n604), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT90), .A4(new_n611), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n548), .A3(new_n654), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n501), .A2(new_n512), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n279), .B1(new_n544), .B2(new_n535), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(G179), .B2(new_n536), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n676), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n538), .B(KEYINPUT91), .C1(new_n501), .C2(new_n512), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n606), .B1(new_n675), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n652), .A2(new_n653), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT26), .B1(new_n674), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n686), .A2(new_n613), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n668), .B1(new_n477), .B2(new_n692), .ZN(G369));
  NAND3_X1  g0493(.A1(new_n221), .A2(new_n222), .A3(G13), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n682), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n549), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n680), .A2(new_n681), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n700), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n513), .A2(new_n518), .A3(new_n699), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n541), .A2(new_n542), .A3(new_n548), .A4(new_n708), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n539), .A2(new_n700), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n570), .A2(new_n700), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n682), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n577), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n707), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n234), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n581), .A2(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n229), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n700), .B1(new_n685), .B2(new_n691), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n541), .A2(new_n542), .A3(new_n683), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n647), .A2(new_n648), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n624), .A2(new_n634), .A3(new_n641), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n686), .B(new_n548), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n670), .A2(new_n671), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n610), .A3(new_n673), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n606), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n674), .A2(KEYINPUT26), .A3(new_n687), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n689), .B1(new_n686), .B2(new_n613), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n606), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT29), .A3(new_n700), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n728), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n614), .A2(new_n654), .A3(new_n700), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n549), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT93), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n523), .A2(new_n597), .A3(new_n527), .A4(new_n601), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n554), .A2(G179), .A3(new_n535), .A4(new_n555), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT30), .B1(new_n749), .B2(new_n633), .ZN(new_n750));
  AOI21_X1  g0550(.A(G179), .B1(new_n597), .B2(new_n601), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n556), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n752), .A2(new_n536), .A3(new_n633), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n746), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n749), .A2(KEYINPUT30), .A3(new_n633), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n645), .A2(new_n545), .A3(new_n556), .A4(new_n751), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n645), .A2(new_n748), .A3(new_n747), .ZN(new_n758));
  OAI211_X1 g0558(.A(KEYINPUT93), .B(new_n757), .C1(new_n758), .C2(KEYINPUT30), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n754), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n700), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n757), .B1(new_n758), .B2(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n699), .B1(new_n764), .B2(new_n755), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n761), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(G330), .B1(new_n745), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n743), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n725), .B1(new_n770), .B2(G1), .ZN(G364));
  INV_X1    g0571(.A(G13), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n221), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n720), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n716), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n714), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n231), .B1(G20), .B2(new_n279), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n222), .A2(new_n304), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G190), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n788), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n222), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n787), .A2(new_n214), .B1(new_n209), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n222), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G87), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n793), .A2(new_n788), .A3(G200), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n322), .C1(new_n490), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT97), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n784), .A2(G190), .A3(new_n330), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G190), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n784), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n801), .A2(G58), .B1(new_n804), .B2(G77), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n785), .A2(new_n788), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n274), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT32), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n793), .A2(new_n802), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n810), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(KEYINPUT32), .A3(G159), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n808), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n792), .A2(new_n799), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G322), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n800), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n292), .B1(new_n803), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(G329), .C2(new_n813), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n806), .A2(G326), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n786), .A2(new_n823), .B1(new_n795), .B2(G303), .ZN(new_n824));
  INV_X1    g0624(.A(new_n790), .ZN(new_n825));
  INV_X1    g0625(.A(new_n797), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n825), .A2(G294), .B1(new_n826), .B2(G283), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n821), .A2(new_n822), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n783), .B1(new_n816), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n776), .B(KEYINPUT94), .Z(new_n830));
  NAND2_X1  g0630(.A1(new_n234), .A2(new_n322), .ZN(new_n831));
  INV_X1    g0631(.A(G355), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n832), .B1(G116), .B2(new_n234), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n719), .A2(new_n322), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n281), .B2(new_n230), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n252), .A2(G45), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(G13), .A2(G33), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT95), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(G20), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n782), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n830), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n829), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n841), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n714), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n778), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NOR2_X1   g0649(.A1(new_n328), .A2(new_n699), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n331), .B1(new_n314), .B2(new_n700), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n328), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n726), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n700), .B(new_n852), .C1(new_n685), .C2(new_n691), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n768), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT101), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n776), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n858), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n856), .A2(new_n768), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n840), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n782), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n830), .B1(G77), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT99), .Z(new_n868));
  INV_X1    g0668(.A(G303), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n807), .A2(new_n869), .B1(new_n797), .B2(new_n207), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(G107), .B2(new_n795), .ZN(new_n871));
  INV_X1    g0671(.A(G294), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n800), .A2(new_n872), .B1(new_n810), .B2(new_n819), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n322), .B(new_n873), .C1(G116), .C2(new_n804), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G97), .A2(new_n825), .B1(new_n786), .B2(G283), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n801), .A2(G143), .B1(new_n804), .B2(G159), .ZN(new_n877));
  INV_X1    g0677(.A(G150), .ZN(new_n878));
  INV_X1    g0678(.A(G137), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n877), .B1(new_n787), .B2(new_n878), .C1(new_n879), .C2(new_n807), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT34), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n826), .A2(G68), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n292), .B1(new_n813), .B2(G132), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n825), .A2(G58), .B1(new_n795), .B2(G50), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n880), .A2(new_n881), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n876), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT100), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n782), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n868), .B1(new_n852), .B2(new_n840), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n863), .A2(new_n892), .ZN(G384));
  NOR2_X1   g0693(.A1(new_n773), .A2(new_n221), .ZN(new_n894));
  INV_X1    g0694(.A(G330), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n614), .A2(new_n654), .A3(new_n700), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n896), .A2(new_n541), .A3(new_n542), .A4(new_n548), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n765), .B(KEYINPUT31), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n423), .A2(new_n700), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n451), .A2(KEYINPUT14), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n446), .A2(new_n436), .A3(new_n443), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(new_n454), .ZN(new_n903));
  AOI221_X4 g0703(.A(new_n900), .B1(new_n463), .B2(new_n903), .C1(new_n473), .C2(new_n467), .ZN(new_n904));
  INV_X1    g0704(.A(new_n900), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n463), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n657), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n852), .B(new_n899), .C1(new_n904), .C2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  INV_X1    g0711(.A(new_n697), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n390), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n394), .A2(new_n390), .A3(new_n395), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT18), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n370), .A2(new_n351), .A3(new_n390), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT104), .B(new_n914), .C1(new_n660), .C2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT103), .B1(new_n390), .B2(new_n912), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n915), .A3(new_n913), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT104), .B1(new_n412), .B2(new_n914), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n911), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n402), .A2(KEYINPUT102), .A3(new_n697), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT102), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n390), .B2(new_n912), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n660), .B2(new_n918), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n929), .A2(new_n931), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n923), .A2(new_n915), .A3(KEYINPUT37), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(new_n935), .B1(new_n920), .B2(new_n924), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(KEYINPUT38), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n910), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n470), .A2(KEYINPUT74), .A3(new_n472), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n462), .B1(new_n461), .B2(new_n466), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n906), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n900), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n657), .A2(new_n906), .A3(new_n905), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n934), .B1(new_n397), .B2(new_n411), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n924), .A2(new_n920), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n923), .A2(new_n915), .A3(KEYINPUT37), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n946), .B1(new_n932), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n911), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n937), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n944), .A2(new_n950), .A3(new_n852), .A4(new_n899), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n909), .A2(new_n938), .B1(new_n951), .B2(new_n910), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT105), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n477), .B1(new_n897), .B2(new_n898), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n895), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  INV_X1    g0757(.A(new_n850), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n855), .A2(new_n958), .B1(new_n942), .B2(new_n943), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n950), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n918), .A2(new_n697), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n949), .A2(new_n937), .A3(KEYINPUT39), .ZN(new_n962));
  INV_X1    g0762(.A(new_n937), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n412), .A2(new_n914), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT104), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n919), .A3(new_n925), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n963), .B1(new_n967), .B2(new_n911), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n962), .B1(new_n968), .B2(KEYINPUT39), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n455), .A2(new_n700), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n960), .B(new_n961), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n728), .B(new_n742), .C1(new_n475), .C2(new_n476), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n668), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n894), .B1(new_n957), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n957), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n619), .A2(KEYINPUT35), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n619), .A2(KEYINPUT35), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n977), .A2(G116), .A3(new_n232), .A4(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT36), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n229), .A2(new_n216), .A3(new_n377), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G68), .B2(new_n201), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n772), .A2(G1), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n976), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT106), .Z(G367));
  NAND2_X1  g0785(.A1(new_n608), .A2(new_n611), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n699), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n606), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n674), .B2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n841), .ZN(new_n990));
  INV_X1    g0790(.A(new_n830), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n234), .A2(new_n312), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n843), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n834), .A2(new_n245), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(G143), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n996), .A2(new_n807), .B1(new_n787), .B2(new_n811), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n322), .B1(new_n800), .B2(new_n878), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n803), .A2(new_n201), .B1(new_n810), .B2(new_n879), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n797), .A2(new_n216), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G58), .B2(new_n795), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(new_n214), .C2(new_n790), .ZN(new_n1003));
  INV_X1    g0803(.A(G283), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n292), .B1(new_n803), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n800), .A2(new_n869), .B1(new_n810), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n794), .A2(new_n558), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1005), .B(new_n1007), .C1(KEYINPUT46), .C2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n786), .A2(G294), .B1(new_n826), .B2(G97), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G107), .A2(new_n825), .B1(new_n806), .B2(G311), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1008), .A2(KEYINPUT46), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1003), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(KEYINPUT47), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT47), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n782), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n990), .B(new_n995), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT113), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n686), .B1(new_n730), .B2(new_n731), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n700), .B1(new_n624), .B2(new_n641), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT107), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n686), .A2(new_n700), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n1026));
  OR3_X1    g0826(.A1(new_n1025), .A2(new_n706), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n1025), .B2(new_n706), .ZN(new_n1028));
  AOI21_X1  g0828(.A(KEYINPUT44), .B1(new_n1025), .B2(new_n706), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT110), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1027), .A2(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1029), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1025), .A2(KEYINPUT44), .A3(new_n706), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(KEYINPUT110), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n717), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n717), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n709), .A2(new_n710), .A3(new_n701), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT111), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n703), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n715), .A2(KEYINPUT112), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n715), .B(KEYINPUT112), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1043), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(new_n769), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1019), .B1(new_n1038), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1050), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1036), .A2(new_n1037), .A3(new_n1052), .A4(KEYINPUT113), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n770), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n720), .B(KEYINPUT41), .Z(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n775), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT43), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n989), .A2(new_n1058), .ZN(new_n1059));
  OR3_X1    g0859(.A1(new_n1025), .A2(KEYINPUT42), .A3(new_n703), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT42), .B1(new_n1025), .B2(new_n703), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n541), .A2(new_n542), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n687), .B1(new_n1023), .B2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1060), .B(new_n1061), .C1(new_n699), .C2(new_n1063), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n989), .A2(new_n1058), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1059), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1025), .A2(new_n717), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(KEYINPUT108), .A3(new_n1070), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1067), .A2(new_n1070), .A3(new_n1068), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT108), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1018), .B1(new_n1057), .B2(new_n1076), .ZN(G387));
  NAND2_X1  g0877(.A1(new_n1049), .A2(new_n769), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1052), .A2(new_n720), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1049), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n709), .A2(new_n710), .A3(new_n841), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n831), .A2(new_n722), .B1(G107), .B2(new_n234), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n242), .A2(new_n281), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n722), .ZN(new_n1084));
  AOI211_X1 g0884(.A(G45), .B(new_n1084), .C1(G68), .C2(G77), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n256), .A2(G50), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT50), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n835), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1082), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n830), .B1(new_n1089), .B2(new_n843), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n292), .B1(new_n813), .B2(G150), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n216), .B2(new_n794), .C1(new_n209), .C2(new_n797), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n801), .A2(G50), .B1(new_n804), .B2(G68), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n256), .B2(new_n787), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G159), .B2(new_n806), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n591), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1093), .B(new_n1096), .C1(new_n1097), .C2(new_n790), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n825), .A2(G283), .B1(new_n795), .B2(G294), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n801), .A2(G317), .B1(new_n804), .B2(G303), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n787), .B2(new_n819), .C1(new_n817), .C2(new_n807), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT115), .Z(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(KEYINPUT49), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n322), .B1(new_n813), .B2(G326), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n558), .C2(new_n797), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT49), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1098), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1090), .B1(new_n1110), .B2(new_n782), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1080), .A2(new_n775), .B1(new_n1081), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1079), .A2(new_n1112), .ZN(G393));
  NAND3_X1  g0913(.A1(new_n1038), .A2(new_n1019), .A3(new_n1050), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1037), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n1035), .A3(new_n1050), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT113), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n720), .B1(new_n1038), .B2(new_n1050), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1036), .A2(new_n774), .A3(new_n1037), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n843), .B1(G97), .B2(new_n719), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n834), .A2(new_n249), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n991), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n807), .A2(new_n878), .B1(new_n811), .B2(new_n800), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT51), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n787), .A2(new_n201), .B1(new_n207), .B2(new_n797), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n322), .B1(new_n810), .B2(new_n996), .C1(new_n256), .C2(new_n803), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n790), .A2(new_n216), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n794), .A2(new_n214), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n807), .A2(new_n1006), .B1(new_n819), .B2(new_n800), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT52), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n787), .A2(new_n869), .B1(new_n558), .B2(new_n790), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n292), .B1(new_n810), .B2(new_n817), .C1(new_n872), .C2(new_n803), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n490), .A2(new_n797), .B1(new_n794), .B2(new_n1004), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1127), .A2(new_n1132), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1125), .B1(new_n783), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1025), .B2(new_n841), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1122), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1121), .A2(new_n1142), .ZN(G390));
  AOI21_X1  g0943(.A(KEYINPUT39), .B1(new_n928), .B2(new_n937), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n962), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n970), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1144), .A2(new_n1145), .B1(new_n1146), .B2(new_n959), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n851), .A2(new_n328), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n741), .A2(new_n700), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n958), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n944), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1146), .B1(new_n928), .B2(new_n937), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(G330), .B(new_n852), .C1(new_n745), .C2(new_n767), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n943), .B2(new_n942), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1147), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n855), .A2(new_n958), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n904), .A2(new_n907), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n970), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n969), .A2(new_n1161), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n853), .B1(new_n942), .B2(new_n943), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n775), .B(new_n1157), .C1(new_n1162), .C2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n830), .B1(new_n257), .B2(new_n866), .ZN(new_n1167));
  INV_X1    g0967(.A(G125), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n322), .B1(new_n810), .B2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n787), .A2(new_n879), .B1(new_n201), .B2(new_n797), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n807), .A2(new_n1171), .B1(new_n811), .B2(new_n790), .ZN(new_n1172));
  INV_X1    g0972(.A(G132), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n800), .A2(new_n1173), .B1(new_n803), .B2(new_n1174), .ZN(new_n1175));
  OR4_X1    g0975(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n795), .A2(G150), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT53), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1130), .B1(G283), .B2(new_n806), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n490), .B2(new_n787), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n803), .A2(new_n209), .B1(new_n810), .B2(new_n872), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n322), .B(new_n1181), .C1(G116), .C2(new_n801), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n796), .A3(new_n883), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1176), .A2(new_n1178), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1167), .B1(new_n1184), .B2(new_n782), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n840), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1166), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT117), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1155), .A2(new_n1150), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n765), .B(new_n761), .ZN(new_n1192));
  OAI211_X1 g0992(.A(KEYINPUT116), .B(G330), .C1(new_n1192), .C2(new_n745), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n852), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT116), .B1(new_n899), .B2(G330), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1160), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1154), .A2(new_n943), .A3(new_n942), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n852), .B1(new_n904), .B2(new_n907), .ZN(new_n1198));
  OAI21_X1  g0998(.A(G330), .B1(new_n1192), .B2(new_n745), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1191), .A2(new_n1196), .B1(new_n1200), .B2(new_n1158), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1164), .B1(new_n475), .B2(new_n476), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n972), .A2(new_n668), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1190), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n853), .B1(new_n1164), .B2(KEYINPUT116), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT116), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1199), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n944), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n958), .B(new_n1149), .C1(new_n1160), .C2(new_n1154), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1163), .A2(new_n1164), .B1(new_n1160), .B2(new_n1154), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1208), .A2(new_n1209), .B1(new_n1210), .B2(new_n1159), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n972), .A2(new_n668), .A3(new_n1202), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(KEYINPUT117), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1204), .A2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1147), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1165), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n720), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1157), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1204), .B2(new_n1213), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1189), .B1(new_n1218), .B2(new_n1220), .ZN(G378));
  NAND2_X1  g1021(.A1(new_n938), .A2(new_n909), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n951), .A2(new_n910), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(G330), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n663), .A2(new_n306), .A3(new_n666), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT118), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT118), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n663), .A2(new_n1227), .A3(new_n306), .A4(new_n666), .ZN(new_n1228));
  XOR2_X1   g1028(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1226), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1231), .A2(new_n1232), .B1(new_n278), .B2(new_n697), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1229), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n278), .A2(new_n697), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1226), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1224), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n960), .A2(new_n961), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1146), .B2(new_n1186), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1243), .A2(G330), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1240), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1242), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(KEYINPUT57), .C1(new_n1220), .C2(new_n1203), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1203), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1224), .A2(new_n1239), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1243), .B1(new_n952), .B2(G330), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n971), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1240), .A2(new_n1244), .A3(new_n1242), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1249), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1248), .A2(new_n1256), .A3(new_n720), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n860), .B1(new_n865), .B2(new_n201), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1168), .A2(new_n807), .B1(new_n787), .B2(new_n1173), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n801), .A2(G128), .B1(new_n804), .B2(G137), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n794), .B2(new_n1174), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1259), .B(new_n1261), .C1(G150), .C2(new_n825), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n826), .A2(G159), .ZN(new_n1266));
  AOI211_X1 g1066(.A(G33), .B(G41), .C1(new_n813), .C2(G124), .ZN(new_n1267));
  AND4_X1   g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n807), .A2(new_n558), .B1(new_n797), .B2(new_n376), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(G97), .B2(new_n786), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n790), .A2(new_n214), .B1(new_n794), .B2(new_n216), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n322), .A2(G41), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n490), .B2(new_n800), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1271), .B(new_n1273), .C1(G283), .C2(new_n813), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1270), .B(new_n1274), .C1(new_n1097), .C2(new_n803), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT58), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI211_X1 g1077(.A(G50), .B(new_n1272), .C1(new_n258), .C2(new_n280), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(new_n1268), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1258), .B1(new_n783), .B2(new_n1280), .C1(new_n1239), .C2(new_n840), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT119), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1253), .A2(new_n775), .A3(new_n1254), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1257), .A2(new_n1284), .ZN(G375));
  NAND2_X1  g1085(.A1(new_n1160), .A2(new_n864), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n830), .B1(G68), .B2(new_n866), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n787), .A2(new_n558), .B1(new_n794), .B2(new_n209), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1001), .B(new_n1288), .C1(G294), .C2(new_n806), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n800), .A2(new_n1004), .B1(new_n803), .B2(new_n490), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n322), .B(new_n1290), .C1(G303), .C2(new_n813), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1289), .B(new_n1291), .C1(new_n1097), .C2(new_n790), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n794), .A2(new_n811), .B1(new_n810), .B2(new_n1171), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(KEYINPUT121), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n1173), .A2(new_n807), .B1(new_n787), .B2(new_n1174), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n322), .B1(new_n803), .B2(new_n878), .C1(new_n879), .C2(new_n800), .ZN(new_n1296));
  OAI22_X1  g1096(.A1(new_n790), .A2(new_n274), .B1(new_n797), .B2(new_n376), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1292), .A2(KEYINPUT120), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(KEYINPUT120), .B2(new_n1292), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1287), .B1(new_n1300), .B2(new_n782), .ZN(new_n1301));
  XOR2_X1   g1101(.A(new_n1301), .B(KEYINPUT122), .Z(new_n1302));
  AOI22_X1  g1102(.A1(new_n1211), .A2(new_n775), .B1(new_n1286), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1056), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1214), .B2(new_n1305), .ZN(G381));
  NOR2_X1   g1106(.A1(G375), .A2(G378), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1071), .A2(new_n1075), .A3(new_n1072), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1055), .B1(new_n1118), .B2(new_n770), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n775), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(G393), .A2(G396), .ZN(new_n1311));
  INV_X1    g1111(.A(G384), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(G390), .A2(G381), .A3(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1307), .A2(new_n1018), .A3(new_n1310), .A4(new_n1314), .ZN(G407));
  NAND2_X1  g1115(.A1(new_n1307), .A2(new_n698), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(G407), .A2(G213), .A3(new_n1316), .ZN(G409));
  AOI21_X1  g1117(.A(new_n848), .B1(new_n1079), .B2(new_n1112), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1311), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1119), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1142), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1319), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1121), .A2(new_n1323), .A3(new_n1142), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G387), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1310), .A2(new_n1018), .A3(new_n1322), .A4(new_n1324), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT125), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1303), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1201), .A2(KEYINPUT60), .A3(new_n1203), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n720), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1204), .A2(KEYINPUT60), .A3(new_n1213), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1304), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT124), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1332), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1333), .A2(KEYINPUT124), .A3(new_n1304), .ZN(new_n1337));
  AOI211_X1 g1137(.A(new_n1312), .B(new_n1330), .C1(new_n1336), .C2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1332), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n1337), .A3(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G384), .B1(new_n1341), .B2(new_n1303), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1329), .B1(new_n1338), .B2(new_n1342), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1333), .A2(KEYINPUT124), .A3(new_n1304), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT124), .B1(new_n1333), .B2(new_n1304), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1344), .A2(new_n1345), .A3(new_n1332), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1312), .B1(new_n1346), .B2(new_n1330), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1341), .A2(G384), .A3(new_n1303), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1347), .A2(KEYINPUT125), .A3(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(G375), .A2(G378), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT123), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1283), .A2(new_n1351), .A3(new_n1281), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1351), .B1(new_n1283), .B2(new_n1281), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1250), .A2(new_n1255), .A3(new_n1055), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1355), .A2(G378), .ZN(new_n1356));
  AOI22_X1  g1156(.A1(new_n1354), .A2(new_n1356), .B1(G213), .B2(new_n698), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1343), .A2(new_n1349), .A3(new_n1350), .A4(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(KEYINPUT62), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1283), .A2(new_n1281), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(KEYINPUT123), .ZN(new_n1361));
  AND2_X1   g1161(.A1(new_n1204), .A2(new_n1213), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n721), .B1(new_n1362), .B2(new_n1219), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1188), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  OAI211_X1 g1165(.A(new_n1247), .B(new_n1056), .C1(new_n1220), .C2(new_n1203), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1283), .A2(new_n1351), .A3(new_n1281), .ZN(new_n1367));
  NAND4_X1  g1167(.A1(new_n1361), .A2(new_n1365), .A3(new_n1366), .A4(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n698), .A2(G213), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1368), .A2(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1365), .B1(new_n1257), .B2(new_n1284), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT62), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1372), .A2(new_n1373), .A3(new_n1349), .A4(new_n1343), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1359), .A2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT61), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n698), .A2(G213), .A3(G2897), .ZN(new_n1377));
  AND3_X1   g1177(.A1(new_n1343), .A2(new_n1377), .A3(new_n1349), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1338), .A2(new_n1342), .ZN(new_n1379));
  OAI22_X1  g1179(.A1(new_n1379), .A2(new_n1377), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1380));
  OAI21_X1  g1180(.A(new_n1376), .B1(new_n1378), .B2(new_n1380), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1328), .B1(new_n1375), .B2(new_n1381), .ZN(new_n1382));
  NOR2_X1   g1182(.A1(new_n1379), .A2(new_n1377), .ZN(new_n1383));
  NOR2_X1   g1183(.A1(new_n1383), .A2(new_n1372), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1343), .A2(new_n1349), .A3(new_n1377), .ZN(new_n1385));
  AOI21_X1  g1185(.A(KEYINPUT61), .B1(new_n1384), .B2(new_n1385), .ZN(new_n1386));
  XNOR2_X1  g1186(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1387));
  AOI21_X1  g1187(.A(new_n1328), .B1(new_n1358), .B2(new_n1387), .ZN(new_n1388));
  NAND4_X1  g1188(.A1(new_n1372), .A2(KEYINPUT63), .A3(new_n1349), .A4(new_n1343), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1386), .A2(new_n1388), .A3(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1382), .A2(new_n1390), .ZN(G405));
  NOR2_X1   g1191(.A1(new_n1307), .A2(new_n1371), .ZN(new_n1392));
  NAND3_X1  g1192(.A1(new_n1392), .A2(new_n1349), .A3(new_n1343), .ZN(new_n1393));
  OAI22_X1  g1193(.A1(new_n1307), .A2(new_n1371), .B1(new_n1342), .B2(new_n1338), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1393), .A2(new_n1394), .ZN(new_n1395));
  INV_X1    g1195(.A(new_n1328), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1396), .A2(KEYINPUT127), .ZN(new_n1397));
  INV_X1    g1197(.A(KEYINPUT127), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1328), .A2(new_n1398), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1395), .A2(new_n1397), .A3(new_n1399), .ZN(new_n1400));
  NAND4_X1  g1200(.A1(new_n1393), .A2(new_n1396), .A3(KEYINPUT127), .A4(new_n1394), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1400), .A2(new_n1401), .ZN(G402));
endmodule


