//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(KEYINPUT70), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(KEYINPUT70), .B2(new_n188), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT71), .B1(new_n195), .B2(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(G110), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(KEYINPUT73), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(G125), .A3(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT16), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n207), .B2(KEYINPUT16), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n206), .A2(G146), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n201), .A2(G140), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n207), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n207), .B2(new_n213), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n199), .A2(new_n211), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n198), .A2(KEYINPUT72), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT23), .B1(new_n187), .B2(G119), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(new_n197), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT72), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n223), .A3(G110), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n191), .A2(new_n192), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n206), .A2(new_n210), .A3(new_n209), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n212), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n228), .A2(new_n211), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n218), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G953), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT22), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(G137), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n218), .B(new_n234), .C1(new_n226), .C2(new_n229), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n237), .A4(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G217), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G234), .B2(new_n237), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n236), .A2(new_n238), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n251), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n212), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(KEYINPUT1), .A3(G146), .ZN(new_n263));
  XNOR2_X1  g077(.A(G143), .B(G146), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n262), .B(new_n263), .C1(G128), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n261), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n187), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n269), .A2(KEYINPUT66), .A3(new_n263), .A4(new_n262), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT11), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT11), .A3(G134), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(G137), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n274), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n275), .A2(G134), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n273), .A2(G137), .ZN(new_n281));
  OAI21_X1  g095(.A(G131), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n271), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT64), .B1(new_n195), .B2(G116), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G119), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n285), .A2(new_n288), .B1(G116), .B2(new_n195), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT2), .B(G113), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n274), .A2(new_n278), .A3(new_n276), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G131), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n279), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n295));
  AND2_X1   g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n259), .A2(new_n261), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G128), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n264), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n294), .A2(new_n300), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT65), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n284), .A2(new_n291), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n283), .A2(new_n265), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT30), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n284), .A2(new_n301), .A3(new_n303), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(KEYINPUT30), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n257), .B(new_n304), .C1(new_n309), .C2(new_n291), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT31), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n284), .A2(new_n291), .A3(new_n302), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n291), .B1(new_n302), .B2(new_n305), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n294), .A2(new_n295), .A3(new_n300), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n295), .B1(new_n294), .B2(new_n300), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n290), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n289), .B(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n271), .B2(new_n283), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n315), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n314), .B(KEYINPUT68), .C1(new_n322), .C2(new_n313), .ZN(new_n323));
  INV_X1    g137(.A(new_n315), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n304), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT28), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n327), .A3(new_n256), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n306), .B1(new_n318), .B2(new_n284), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n320), .B1(new_n329), .B2(new_n307), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT31), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n257), .A4(new_n304), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n311), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(G472), .A2(G902), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n333), .A2(KEYINPUT32), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT32), .B1(new_n333), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n323), .A2(new_n327), .A3(new_n257), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n330), .A2(new_n256), .A3(new_n304), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n308), .A2(new_n320), .B1(new_n321), .B2(new_n318), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT29), .B(new_n314), .C1(new_n343), .C2(new_n313), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT69), .B1(new_n344), .B2(new_n256), .ZN(new_n345));
  INV_X1    g159(.A(new_n314), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n308), .A2(new_n320), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n304), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n348), .B2(KEYINPUT28), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT69), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT29), .A4(new_n257), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n342), .A2(new_n237), .A3(new_n345), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G472), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n250), .B1(new_n337), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G469), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n357), .B2(G107), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G104), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(G107), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n358), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n360), .A2(G104), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n357), .A2(G107), .ZN(new_n366));
  OAI21_X1  g180(.A(G101), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n293), .A2(new_n279), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n265), .A2(new_n364), .A3(new_n367), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n358), .A2(new_n361), .A3(new_n363), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n378), .A3(G101), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n300), .A3(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n231), .A2(G227), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(G110), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n200), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT12), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n368), .A2(new_n263), .A3(new_n262), .A4(new_n269), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n388), .B(new_n371), .C1(new_n372), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n372), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT12), .B1(new_n391), .B2(new_n294), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n356), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n294), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n388), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(KEYINPUT12), .A3(new_n294), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n398), .A2(KEYINPUT80), .A3(new_n381), .A4(new_n386), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n370), .A2(new_n374), .A3(new_n380), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n294), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n386), .B1(new_n402), .B2(new_n381), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n355), .B(new_n237), .C1(new_n400), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(G469), .A2(G902), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT78), .ZN(new_n406));
  INV_X1    g220(.A(new_n381), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(new_n393), .ZN(new_n408));
  INV_X1    g222(.A(new_n386), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n398), .A2(KEYINPUT78), .A3(new_n381), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n387), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n381), .A2(new_n386), .A3(KEYINPUT79), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n402), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(G469), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n404), .A2(new_n405), .A3(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT9), .B(G234), .Z(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT76), .ZN(new_n419));
  OAI21_X1  g233(.A(G221), .B1(new_n419), .B2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G475), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n357), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT19), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n215), .B2(new_n216), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n202), .A2(KEYINPUT19), .A3(new_n204), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n212), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n211), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT87), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n252), .A2(G214), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G143), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n260), .A2(KEYINPUT85), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n252), .A2(KEYINPUT85), .A3(new_n260), .A4(G214), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n277), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(G131), .A3(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n441), .A3(new_n211), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n430), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(KEYINPUT18), .A2(G131), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT86), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n446));
  INV_X1    g260(.A(new_n444), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n435), .A2(new_n446), .A3(new_n447), .A4(new_n436), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n437), .A2(new_n444), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n217), .B1(new_n212), .B2(new_n205), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n424), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n424), .B(KEYINPUT88), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n435), .A2(KEYINPUT17), .A3(G131), .A4(new_n436), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT89), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT17), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n438), .A2(new_n458), .A3(new_n439), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n228), .A3(new_n211), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n452), .B(new_n454), .C1(new_n457), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n422), .B(new_n237), .C1(new_n453), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n442), .A2(new_n440), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n441), .B1(new_n428), .B2(new_n211), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n452), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n424), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n461), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n471), .A2(KEYINPUT20), .A3(new_n422), .A4(new_n237), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n474));
  INV_X1    g288(.A(G478), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT15), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(G116), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT91), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(KEYINPUT92), .A3(new_n481), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n485), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n287), .A2(G122), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(KEYINPUT14), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n483), .A2(new_n484), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G107), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n260), .A2(G128), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n187), .A2(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G134), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n493), .A3(new_n273), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n479), .A2(new_n488), .A3(new_n360), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT90), .Z(new_n499));
  NAND3_X1  g313(.A1(new_n491), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n479), .A2(new_n488), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G107), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n498), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n493), .B1(new_n492), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT13), .B1(new_n260), .B2(G128), .ZN(new_n506));
  OAI21_X1  g320(.A(G134), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n507), .A3(new_n496), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n419), .A2(new_n244), .A3(G953), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n508), .A3(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n477), .B1(new_n514), .B2(new_n237), .ZN(new_n515));
  AOI211_X1 g329(.A(G902), .B(new_n476), .C1(new_n512), .C2(new_n513), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n474), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n500), .A2(new_n508), .A3(new_n510), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n510), .B1(new_n500), .B2(new_n508), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n237), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n476), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n237), .A3(new_n477), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT93), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(G234), .A2(G237), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(G952), .A3(new_n231), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT21), .B(G898), .Z(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(G902), .A3(G953), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n229), .A2(new_n459), .A3(new_n456), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n424), .B1(new_n530), .B2(new_n452), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n237), .B1(new_n462), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G475), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n473), .A2(new_n524), .A3(new_n529), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n285), .A2(new_n288), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n195), .A2(G116), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(KEYINPUT5), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n536), .A2(KEYINPUT5), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(G113), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n289), .A2(new_n319), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n369), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n377), .A2(new_n379), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n291), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G122), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n541), .B(new_n544), .C1(new_n542), .C2(new_n291), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT6), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT6), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n549), .A3(new_n545), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n299), .A2(G125), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n269), .A2(new_n201), .A3(new_n263), .A4(new_n262), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n231), .A2(G224), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(KEYINPUT81), .Z(new_n555));
  XOR2_X1   g369(.A(new_n553), .B(new_n555), .Z(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n539), .A2(new_n540), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n368), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(KEYINPUT83), .A3(new_n541), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n541), .A2(KEYINPUT83), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n544), .B(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n551), .A2(new_n552), .B1(KEYINPUT84), .B2(new_n555), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n555), .A2(KEYINPUT7), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n565), .B(new_n566), .Z(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n567), .A3(new_n547), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n557), .A2(new_n568), .A3(new_n237), .ZN(new_n569));
  OAI21_X1  g383(.A(G210), .B1(G237), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n557), .A2(new_n568), .A3(new_n237), .A4(new_n570), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G214), .B1(G237), .B2(G902), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n421), .A2(new_n534), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n354), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G101), .ZN(G3));
  NAND2_X1  g393(.A1(new_n333), .A2(new_n237), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n333), .A2(new_n334), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n583), .A2(new_n250), .A3(new_n421), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n465), .A2(new_n533), .A3(new_n472), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT95), .B1(new_n500), .B2(new_n508), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n587), .A2(new_n512), .A3(KEYINPUT33), .A4(new_n513), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  OAI22_X1  g403(.A1(new_n518), .A2(new_n519), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n588), .A2(new_n590), .A3(G478), .A4(new_n237), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n520), .A2(new_n475), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n585), .B(new_n529), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n573), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n569), .A2(new_n599), .A3(new_n571), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n575), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n584), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(KEYINPUT97), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT34), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G104), .ZN(G6));
  INV_X1    g420(.A(new_n529), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n524), .A2(new_n585), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n584), .A2(new_n602), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n333), .B2(new_n237), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n333), .B2(new_n334), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n417), .A2(new_n420), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n517), .A2(new_n523), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n616), .A2(new_n585), .A3(new_n607), .ZN(new_n617));
  INV_X1    g431(.A(new_n576), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n614), .A2(new_n615), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n235), .A2(KEYINPUT36), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n230), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n230), .A2(new_n620), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n243), .A2(new_n245), .B1(new_n248), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT98), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT37), .B(G110), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G12));
  AOI21_X1  g442(.A(new_n624), .B1(new_n337), .B2(new_n353), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n528), .A2(G900), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n526), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n585), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n616), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT99), .B1(new_n634), .B2(new_n601), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n524), .A2(new_n585), .A3(new_n632), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n602), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n629), .A2(new_n635), .A3(new_n615), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  XNOR2_X1  g454(.A(new_n631), .B(KEYINPUT39), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n615), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT40), .Z(new_n643));
  AOI21_X1  g457(.A(new_n256), .B1(new_n330), .B2(new_n304), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n237), .B1(new_n348), .B2(new_n257), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n337), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n624), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n574), .B(KEYINPUT38), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n616), .A2(new_n585), .ZN(new_n652));
  INV_X1    g466(.A(new_n575), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n643), .A2(new_n650), .A3(new_n651), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  OAI211_X1 g470(.A(new_n585), .B(new_n631), .C1(new_n593), .C2(new_n595), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n629), .A2(new_n615), .A3(new_n602), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT100), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  OAI21_X1  g475(.A(new_n237), .B1(new_n400), .B2(new_n403), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G469), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n420), .A3(new_n404), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT101), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n663), .A2(new_n666), .A3(new_n420), .A4(new_n404), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n602), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n354), .A3(new_n597), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  INV_X1    g485(.A(new_n250), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT32), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n582), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n333), .A2(KEYINPUT32), .A3(new_n334), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n351), .A2(new_n345), .ZN(new_n677));
  AOI21_X1  g491(.A(G902), .B1(new_n340), .B2(new_n341), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n612), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n672), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n668), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n597), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT41), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G113), .ZN(G15));
  NAND2_X1  g500(.A1(new_n681), .A2(new_n608), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT103), .B(G116), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G18));
  AOI211_X1 g503(.A(new_n624), .B(new_n534), .C1(new_n337), .C2(new_n353), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n669), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  OAI21_X1  g506(.A(new_n314), .B1(new_n343), .B2(new_n313), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n256), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n311), .A2(new_n694), .A3(new_n332), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n695), .A2(new_n334), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n250), .A2(new_n696), .A3(new_n613), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n652), .A2(new_n607), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n669), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  NOR4_X1   g516(.A1(new_n657), .A2(new_n696), .A3(new_n613), .A4(new_n624), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n602), .A3(new_n667), .A4(new_n665), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  NAND3_X1  g519(.A1(new_n572), .A2(new_n575), .A3(new_n573), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n572), .A2(KEYINPUT107), .A3(new_n575), .A4(new_n573), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n405), .B(KEYINPUT105), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n404), .A2(new_n416), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n420), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n420), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n354), .A3(new_n658), .A4(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n708), .A2(new_n709), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n420), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT106), .B1(new_n713), .B2(new_n420), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n680), .A3(new_n657), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n722), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND3_X1  g544(.A1(new_n718), .A2(new_n354), .A3(new_n636), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  OR2_X1    g546(.A1(new_n593), .A2(new_n595), .ZN(new_n733));
  INV_X1    g547(.A(new_n585), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(KEYINPUT43), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n583), .A3(new_n649), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n723), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n411), .A2(new_n415), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n748), .B2(new_n712), .ZN(new_n749));
  INV_X1    g563(.A(new_n404), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n420), .A3(new_n641), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n742), .A2(new_n755), .A3(new_n723), .A4(new_n743), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n745), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G137), .ZN(G39));
  NAND3_X1  g572(.A1(new_n337), .A2(new_n353), .A3(new_n250), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n657), .A3(new_n710), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT110), .Z(new_n761));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n753), .B2(new_n420), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n420), .ZN(new_n765));
  AOI211_X1 g579(.A(KEYINPUT47), .B(new_n765), .C1(new_n751), .C2(new_n752), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT111), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n200), .ZN(G42));
  NAND2_X1  g584(.A1(new_n663), .A2(new_n404), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT49), .Z(new_n772));
  NOR2_X1   g586(.A1(new_n735), .A2(new_n651), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n250), .A2(new_n653), .A3(new_n765), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n648), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n665), .A2(new_n667), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n723), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n696), .A2(new_n613), .A3(new_n624), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n526), .B1(new_n737), .B2(new_n738), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n648), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n250), .A2(new_n526), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n781), .A2(new_n585), .A3(new_n733), .A4(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n699), .A2(new_n779), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n651), .A2(new_n575), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n776), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n784), .A2(new_n776), .A3(new_n790), .A4(new_n785), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n783), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n764), .A2(new_n767), .A3(KEYINPUT116), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n663), .A2(new_n765), .A3(new_n404), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n763), .B2(new_n766), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n784), .A2(new_n723), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n780), .B(new_n792), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n794), .B1(new_n763), .B2(new_n766), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n723), .A3(new_n784), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n792), .A2(new_n803), .A3(KEYINPUT51), .A4(new_n780), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n699), .A2(new_n779), .A3(new_n669), .ZN(new_n805));
  INV_X1    g619(.A(G952), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT118), .B1(new_n806), .B2(G953), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n781), .A2(new_n782), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n733), .A2(new_n585), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n805), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n777), .A2(new_n354), .A3(new_n779), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT48), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n811), .A2(KEYINPUT48), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n801), .A2(new_n804), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n614), .A2(new_n615), .A3(new_n672), .A4(new_n618), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n734), .B(new_n529), .C1(new_n515), .C2(new_n516), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n624), .A2(new_n619), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n680), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n581), .A2(new_n582), .A3(new_n420), .A4(new_n417), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n823), .A2(new_n250), .A3(new_n576), .A4(new_n596), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n584), .A2(new_n618), .A3(new_n597), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(KEYINPUT112), .A3(new_n578), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n819), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n681), .A2(new_n608), .B1(new_n690), .B2(new_n669), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n684), .A3(new_n701), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n515), .A2(new_n516), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n633), .A2(new_n708), .A3(new_n831), .A4(new_n709), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n624), .B(new_n421), .C1(new_n337), .C2(new_n353), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n834), .A2(new_n835), .B1(new_n703), .B2(new_n718), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n729), .A2(new_n731), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT114), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n682), .B1(new_n681), .B2(new_n597), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n668), .A2(new_n680), .A3(KEYINPUT102), .A4(new_n596), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n829), .B(new_n701), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n729), .A2(new_n731), .A3(new_n836), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n828), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n659), .A2(new_n704), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n714), .A2(new_n652), .A3(new_n601), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n647), .A3(new_n624), .A4(new_n631), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n847), .A3(new_n639), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n639), .A2(new_n659), .A3(new_n704), .A4(new_n849), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n838), .A2(new_n845), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n852), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n830), .A2(new_n837), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n816), .B1(new_n857), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT53), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n830), .A2(new_n853), .A3(new_n856), .A4(new_n837), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n867), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(KEYINPUT118), .A2(G953), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n815), .A2(new_n866), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(G952), .A2(G953), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n775), .B1(new_n871), .B2(new_n872), .ZN(G75));
  NAND2_X1  g687(.A1(new_n548), .A2(new_n550), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(new_n556), .Z(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n859), .A2(new_n860), .A3(new_n858), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT115), .B1(new_n850), .B2(new_n852), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n842), .A2(new_n843), .A3(new_n828), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n856), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n854), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n237), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(G210), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n877), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g701(.A(KEYINPUT56), .B(new_n876), .C1(new_n884), .C2(G210), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n231), .A2(G952), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT119), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(G51));
  XNOR2_X1  g705(.A(new_n711), .B(KEYINPUT57), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n816), .B1(new_n882), .B2(new_n883), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n893), .B2(new_n869), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n403), .B2(new_n400), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n748), .B(KEYINPUT120), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n889), .B1(new_n895), .B2(new_n897), .ZN(G54));
  NAND3_X1  g712(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n461), .A3(new_n470), .ZN(new_n900));
  INV_X1    g714(.A(new_n889), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .A4(new_n471), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n866), .B2(new_n869), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n588), .A2(new_n590), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n905), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n893), .B2(new_n869), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  INV_X1    g726(.A(new_n890), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n910), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT54), .B1(new_n867), .B2(new_n868), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n881), .B1(new_n861), .B2(new_n862), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n816), .B(new_n883), .C1(new_n917), .C2(KEYINPUT53), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT121), .B1(new_n919), .B2(new_n890), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n909), .A2(new_n914), .A3(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT60), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n623), .B(new_n924), .C1(new_n867), .C2(new_n868), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n882), .B2(new_n883), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n913), .B(new_n925), .C1(new_n926), .C2(new_n247), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT61), .B1(new_n925), .B2(KEYINPUT122), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G66));
  AOI21_X1  g743(.A(new_n231), .B1(new_n527), .B2(G224), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n830), .B2(new_n231), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n874), .B1(G898), .B2(new_n231), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(G69));
  NAND2_X1  g747(.A1(new_n729), .A2(new_n731), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT124), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n846), .A2(new_n639), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n354), .A2(new_n585), .A3(new_n616), .A4(new_n602), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n754), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n935), .A2(new_n757), .A3(new_n768), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n231), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n426), .A2(new_n427), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n309), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n941), .B(new_n944), .C1(G227), .C2(new_n231), .ZN(new_n945));
  OAI21_X1  g759(.A(G900), .B1(new_n944), .B2(G227), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(G953), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n655), .A2(new_n639), .A3(new_n846), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  OAI21_X1  g763(.A(new_n809), .B1(new_n585), .B2(new_n831), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  OR4_X1    g765(.A1(new_n680), .A2(new_n951), .A3(new_n642), .A4(new_n710), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n949), .A2(new_n757), .A3(new_n768), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n231), .A3(new_n943), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n945), .A2(new_n947), .A3(new_n954), .ZN(G72));
  XNOR2_X1  g769(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n612), .A2(new_n237), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n953), .B2(new_n830), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n644), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n940), .B2(new_n830), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n339), .B(KEYINPUT126), .Z(new_n962));
  AND2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n644), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n339), .A3(new_n958), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n857), .B2(new_n865), .ZN(new_n967));
  NOR4_X1   g781(.A1(new_n960), .A2(new_n963), .A3(new_n889), .A4(new_n967), .ZN(G57));
endmodule


