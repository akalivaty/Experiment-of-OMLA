//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n453), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI21_X1  g035(.A(KEYINPUT69), .B1(new_n456), .B2(G2106), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(G567), .B2(new_n458), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n456), .A2(KEYINPUT69), .A3(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n470), .A2(new_n472), .A3(G137), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT70), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G137), .A4(new_n473), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n469), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n470), .A2(new_n472), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n486), .A2(new_n473), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n473), .A2(G112), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n489), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n495), .B(new_n496), .ZN(G162));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(G2105), .B1(KEYINPUT74), .B2(G114), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT74), .A2(G114), .ZN(new_n500));
  OAI211_X1 g075(.A(G2104), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n470), .A2(new_n472), .A3(G126), .A4(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n473), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n476), .A2(new_n509), .A3(G138), .A4(new_n473), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n504), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n515), .A2(new_n517), .A3(G50), .A4(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n520), .A2(new_n522), .A3(new_n515), .A4(new_n517), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n520), .A2(new_n522), .A3(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(new_n520), .A2(new_n522), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT77), .Z(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n515), .A2(new_n517), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n534), .B1(new_n523), .B2(new_n535), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n532), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n530), .A2(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n514), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n537), .A2(new_n544), .B1(new_n545), .B2(new_n523), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n530), .A2(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n514), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT78), .B(G81), .Z(new_n552));
  OAI22_X1  g127(.A1(new_n537), .A2(new_n551), .B1(new_n523), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n520), .A2(new_n522), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT79), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n536), .A2(G53), .A3(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  AND4_X1   g144(.A1(new_n520), .A2(new_n522), .A3(new_n515), .A4(new_n517), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G91), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n573));
  XNOR2_X1  g148(.A(G171), .B(new_n573), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  NAND2_X1  g150(.A1(new_n526), .A2(new_n527), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n530), .A2(G88), .A3(new_n536), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n577), .A2(KEYINPUT81), .A3(new_n578), .A4(new_n518), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n525), .B2(new_n528), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G303));
  NAND2_X1  g157(.A1(new_n570), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n537), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n561), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n570), .B2(G86), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n515), .A2(new_n517), .A3(G48), .A4(G543), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n530), .A2(G60), .ZN(new_n595));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n514), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n537), .A2(new_n598), .B1(new_n599), .B2(new_n523), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n561), .B(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n604), .A2(G66), .ZN(new_n605));
  AND2_X1   g180(.A1(G79), .A2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n537), .A2(KEYINPUT83), .ZN(new_n608));
  INV_X1    g183(.A(G54), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n537), .B2(KEYINPUT83), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n570), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n523), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n608), .A2(new_n610), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G301), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G284));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n617), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n617), .B2(G168), .ZN(G297));
  XNOR2_X1  g198(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g199(.A(new_n616), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(new_n554), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n629), .A2(KEYINPUT85), .B1(new_n617), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(KEYINPUT85), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n487), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n473), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(G123), .B2(new_n490), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT86), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n476), .A2(new_n467), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT87), .B(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT15), .B(G2435), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT16), .B(G1341), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n651), .B2(new_n657), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n664), .B1(KEYINPUT89), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(KEYINPUT89), .B2(new_n666), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n671), .C1(new_n662), .C2(new_n663), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT88), .Z(new_n674));
  INV_X1    g249(.A(KEYINPUT18), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n675), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n686), .B1(new_n681), .B2(new_n684), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n689), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1991), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  NAND2_X1  g273(.A1(new_n467), .A2(G105), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n490), .A2(G129), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n487), .A2(G141), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT26), .Z(new_n703));
  AND4_X1   g278(.A1(new_n699), .A2(new_n700), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G29), .B2(G32), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT94), .Z(new_n709));
  INV_X1    g284(.A(G2084), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(KEYINPUT24), .B2(G34), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(KEYINPUT24), .B2(G34), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n484), .B2(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n709), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n710), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n711), .A2(G26), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n490), .A2(G128), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n487), .A2(G140), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n473), .A2(G116), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n717), .B(new_n718), .C1(new_n723), .C2(G29), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n717), .B2(new_n718), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2067), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n715), .A2(new_n716), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(G168), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G21), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT31), .B(G11), .Z(new_n732));
  INV_X1    g307(.A(G28), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n639), .B2(new_n711), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n706), .A2(new_n707), .ZN(new_n738));
  NOR2_X1   g313(.A1(G5), .A2(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G171), .B2(G16), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G1961), .ZN(new_n741));
  NOR4_X1   g316(.A1(new_n731), .A2(new_n737), .A3(new_n738), .A4(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G19), .B(new_n630), .S(G16), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G1341), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(G1341), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n729), .B2(new_n730), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n742), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G33), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n467), .A2(G103), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n487), .A2(G139), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n751), .B(new_n752), .C1(new_n473), .C2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT93), .Z(new_n755));
  AOI21_X1  g330(.A(new_n748), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2072), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n740), .A2(G1961), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT95), .Z(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT101), .ZN(new_n762));
  INV_X1    g337(.A(G20), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1956), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n727), .A2(new_n747), .A3(new_n760), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n711), .A2(G35), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT98), .Z(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n711), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n711), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n711), .ZN(new_n777));
  MUX2_X1   g352(.A(new_n776), .B(new_n777), .S(KEYINPUT96), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2078), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G4), .B(new_n616), .S(G16), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT91), .B(G1348), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n768), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G22), .ZN(new_n790));
  MUX2_X1   g365(.A(new_n790), .B(G166), .S(G16), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1971), .ZN(new_n792));
  MUX2_X1   g367(.A(G23), .B(G288), .S(G16), .Z(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT90), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n789), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n490), .A2(G119), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n487), .A2(G131), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n473), .A2(G107), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G25), .B(new_n803), .S(G29), .Z(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT35), .B(G1991), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G24), .B(G290), .S(G16), .Z(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(G1986), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G1986), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT36), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n773), .A2(new_n774), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT99), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n786), .A2(new_n812), .A3(new_n814), .ZN(G150));
  INV_X1    g390(.A(KEYINPUT102), .ZN(new_n816));
  NAND2_X1  g391(.A1(G150), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n786), .A2(new_n812), .A3(KEYINPUT102), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(G311));
  NAND2_X1  g394(.A1(new_n530), .A2(G67), .ZN(new_n820));
  NAND2_X1  g395(.A1(G80), .A2(G543), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n514), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n537), .A2(new_n823), .B1(new_n824), .B2(new_n523), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G860), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n625), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT103), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n554), .B(new_n826), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n827), .B1(new_n833), .B2(new_n835), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n829), .B1(new_n836), .B2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n803), .B(new_n642), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n484), .B(KEYINPUT104), .Z(new_n840));
  XNOR2_X1  g415(.A(G162), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n487), .A2(G142), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n473), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G130), .B2(new_n490), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n639), .B(new_n846), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n841), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n501), .A2(new_n502), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n511), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n723), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n704), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n754), .ZN(new_n854));
  INV_X1    g429(.A(new_n755), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n853), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n848), .A2(new_n856), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n839), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n841), .B(new_n847), .Z(new_n861));
  INV_X1    g436(.A(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n839), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n848), .A2(new_n856), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n859), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g443(.A(new_n617), .B1(new_n822), .B2(new_n825), .ZN(new_n869));
  INV_X1    g444(.A(G288), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G305), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n601), .B(G166), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT106), .Z(new_n876));
  XOR2_X1   g451(.A(new_n873), .B(KEYINPUT105), .Z(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n878), .B2(new_n874), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n616), .B(G299), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT41), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n628), .B(new_n835), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n879), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n869), .B1(new_n885), .B2(new_n617), .ZN(G295));
  OAI21_X1  g461(.A(new_n869), .B1(new_n885), .B2(new_n617), .ZN(G331));
  NAND2_X1  g462(.A1(G286), .A2(G171), .ZN(new_n888));
  NAND2_X1  g463(.A1(G301), .A2(G168), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n834), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n835), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n880), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n881), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n877), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n860), .B1(new_n895), .B2(new_n877), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n895), .A2(new_n877), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n900), .A2(new_n896), .A3(new_n901), .A4(new_n860), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT44), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n906));
  AOI211_X1 g481(.A(KEYINPUT107), .B(new_n906), .C1(new_n899), .C2(new_n902), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(G397));
  INV_X1    g483(.A(G40), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n482), .B2(G2105), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n479), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT109), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n479), .A2(new_n913), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G1384), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n512), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G2078), .ZN(new_n920));
  AOI21_X1  g495(.A(G1384), .B1(new_n511), .B2(new_n849), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT45), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n915), .A2(new_n919), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT53), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G1961), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n850), .A2(new_n927), .A3(new_n916), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT112), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n921), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI22_X1  g507(.A1(KEYINPUT75), .A2(new_n503), .B1(new_n508), .B2(new_n510), .ZN(new_n933));
  AOI21_X1  g508(.A(G1384), .B1(new_n933), .B2(new_n506), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n479), .A2(new_n913), .A3(new_n910), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n913), .B1(new_n479), .B2(new_n910), .ZN(new_n936));
  OAI22_X1  g511(.A1(new_n934), .A2(new_n927), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n926), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n939));
  INV_X1    g514(.A(new_n921), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n918), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n924), .A2(G2078), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n939), .A2(new_n915), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n925), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT122), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n944), .A2(new_n945), .A3(new_n619), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n944), .B2(new_n619), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n918), .A3(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n911), .A2(new_n924), .A3(G2078), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n922), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n925), .A2(new_n938), .A3(G301), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT54), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n912), .A2(new_n914), .B1(new_n917), .B2(KEYINPUT50), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n503), .B1(new_n508), .B2(new_n510), .ZN(new_n958));
  NOR4_X1   g533(.A1(new_n958), .A2(KEYINPUT112), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n930), .B1(new_n921), .B2(new_n927), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n961), .A3(new_n710), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n935), .A2(new_n936), .B1(KEYINPUT45), .B2(new_n921), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n917), .A2(new_n918), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n963), .B(new_n730), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n939), .A2(new_n915), .A3(new_n941), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n963), .B1(new_n968), .B2(new_n730), .ZN(new_n969));
  OAI21_X1  g544(.A(G8), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(G168), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n972), .B2(KEYINPUT121), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n730), .B1(new_n964), .B2(new_n965), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT115), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(new_n962), .A3(new_n966), .ZN(new_n980));
  OAI211_X1 g555(.A(G8), .B(new_n975), .C1(new_n980), .C2(G286), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n972), .B1(new_n967), .B2(new_n969), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT120), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(new_n984), .A3(new_n972), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n977), .A2(new_n981), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n925), .A2(new_n938), .A3(new_n953), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G171), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n988), .B(KEYINPUT54), .C1(new_n619), .C2(new_n944), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n971), .B1(new_n915), .B2(new_n921), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n870), .A2(G1976), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n590), .B2(new_n593), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n590), .A2(new_n995), .A3(new_n593), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(KEYINPUT49), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  INV_X1    g575(.A(new_n998), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n996), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n990), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n921), .B1(new_n935), .B2(new_n936), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(G8), .A3(new_n991), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n994), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n971), .B1(new_n579), .B2(new_n581), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT55), .B1(new_n1008), .B2(KEYINPUT113), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1008), .A2(KEYINPUT113), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1008), .B2(KEYINPUT113), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND4_X1   g588(.A1(G50), .A2(new_n515), .A3(new_n517), .A4(G543), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n570), .B2(G88), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT81), .B1(new_n1015), .B2(new_n577), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n525), .A2(new_n528), .A3(new_n580), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT113), .B(G8), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT114), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1008), .A2(KEYINPUT113), .A3(new_n1010), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1019), .A2(new_n1022), .A3(KEYINPUT55), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1013), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n957), .A2(new_n961), .A3(new_n774), .ZN(new_n1026));
  INV_X1    g601(.A(G1971), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n922), .B1(new_n935), .B2(new_n936), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n971), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1007), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n912), .A2(new_n914), .B1(KEYINPUT45), .B2(new_n921), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1971), .B1(new_n1033), .B2(new_n919), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT50), .B1(new_n958), .B2(G1384), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n935), .B2(new_n936), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n512), .A2(new_n927), .A3(new_n916), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1036), .A2(G2090), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(G8), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(new_n1024), .A3(new_n1013), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n989), .A2(new_n1032), .A3(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n956), .A2(new_n986), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT61), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT57), .B1(new_n569), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G299), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n569), .A2(new_n571), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n569), .A2(new_n1044), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n567), .B(new_n1047), .C1(new_n1048), .C2(KEYINPUT57), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT56), .B(G2072), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n915), .A2(new_n919), .A3(new_n922), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT118), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1033), .A2(new_n1054), .A3(new_n919), .A4(new_n1051), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n512), .A2(new_n927), .A3(new_n916), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(new_n1035), .C1(new_n936), .C2(new_n935), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND4_X1   g634(.A1(new_n1050), .A2(new_n1053), .A3(new_n1055), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1052), .A2(KEYINPUT118), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1050), .B1(new_n1061), .B2(new_n1055), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1043), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2067), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(new_n921), .C1(new_n935), .C2(new_n936), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n917), .A2(KEYINPUT50), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n915), .A2(new_n1067), .A3(new_n929), .A4(new_n931), .ZN(new_n1068));
  INV_X1    g643(.A(G1348), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1070), .A2(KEYINPUT60), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1072));
  AND4_X1   g647(.A1(KEYINPUT60), .A2(new_n1072), .A3(new_n616), .A4(new_n1065), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n616), .B1(new_n1070), .B2(KEYINPUT60), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1053), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1050), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1061), .A2(new_n1050), .A3(new_n1055), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT61), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1996), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1033), .A2(new_n1081), .A3(new_n919), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT58), .B(G1341), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n1004), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n630), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1063), .A2(new_n1075), .A3(new_n1080), .A4(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1070), .A2(new_n616), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1079), .B1(new_n1062), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(KEYINPUT119), .A3(new_n1090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1042), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1003), .A2(new_n992), .A3(new_n870), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n990), .B1(new_n1096), .B2(new_n1001), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1031), .A2(new_n1025), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n1007), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n994), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1040), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n980), .A2(G8), .A3(G168), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT116), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1102), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1031), .A2(new_n1025), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(new_n1032), .A3(KEYINPUT63), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1099), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n977), .A2(new_n981), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n983), .A2(new_n985), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1032), .B(new_n1040), .C1(new_n946), .C2(new_n947), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(KEYINPUT62), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1111), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n946), .ZN(new_n1121));
  INV_X1    g696(.A(new_n947), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1101), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n986), .B2(new_n1113), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1124), .A2(new_n1115), .A3(KEYINPUT124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1095), .B(new_n1110), .C1(new_n1120), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n915), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n951), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1081), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT110), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n704), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n723), .B(new_n1064), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1081), .B2(new_n704), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1131), .A2(KEYINPUT111), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1131), .A2(KEYINPUT111), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1128), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n803), .B(new_n806), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1134), .B(new_n1135), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n601), .B(G1986), .Z(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1128), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1126), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT46), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1130), .B(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1132), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1128), .B1(new_n852), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT125), .B(KEYINPUT126), .Z(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT47), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1136), .A2(G1986), .A3(G290), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT48), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1149), .A2(new_n1150), .B1(new_n1138), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n803), .A2(new_n805), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1135), .A2(new_n1134), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n723), .A2(G2067), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1136), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1141), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g735(.A1(G227), .A2(new_n464), .A3(G401), .ZN(new_n1162));
  NAND4_X1  g736(.A1(new_n697), .A2(new_n867), .A3(new_n903), .A4(new_n1162), .ZN(G225));
  INV_X1    g737(.A(G225), .ZN(G308));
endmodule


