//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT79), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT80), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(KEYINPUT80), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT2), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n211), .A2(KEYINPUT81), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(KEYINPUT81), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n219), .A2(new_n216), .A3(new_n209), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n218), .A2(new_n221), .ZN(new_n227));
  INV_X1    g026(.A(new_n208), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n223), .B1(new_n228), .B2(KEYINPUT29), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n226), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G78gat), .B(G106gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G228gat), .A2(G233gat), .ZN(new_n233));
  INV_X1    g032(.A(G22gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT31), .B(G50gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n232), .B(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT73), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT34), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT74), .Z(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT27), .B(G183gat), .ZN(new_n242));
  INV_X1    g041(.A(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT28), .B1(new_n244), .B2(KEYINPUT67), .ZN(new_n245));
  INV_X1    g044(.A(G183gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(new_n243), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n249));
  INV_X1    g048(.A(G169gat), .ZN(new_n250));
  INV_X1    g049(.A(G176gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(KEYINPUT26), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n253), .B(KEYINPUT66), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(KEYINPUT26), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n254), .B1(new_n252), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n259), .B2(new_n254), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT24), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(G183gat), .A3(G190gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n247), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT65), .Z(new_n266));
  AOI21_X1  g065(.A(new_n261), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT25), .B(new_n260), .C1(new_n256), .C2(new_n259), .ZN(new_n270));
  INV_X1    g069(.A(new_n265), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n264), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n258), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G120gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n275), .A2(KEYINPUT69), .A3(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G127gat), .ZN(new_n282));
  INV_X1    g081(.A(G134gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n275), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT68), .B(G134gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G127gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n273), .B(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(G227gat), .A2(G233gat), .ZN(new_n290));
  OAI221_X1 g089(.A(new_n241), .B1(new_n239), .B2(KEYINPUT34), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n241), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n281), .A2(new_n287), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n293), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n239), .A2(KEYINPUT34), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  XNOR2_X1  g099(.A(G15gat), .B(G43gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT71), .ZN(new_n302));
  XOR2_X1   g101(.A(G71gat), .B(G99gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n294), .A2(new_n290), .A3(new_n295), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(new_n306), .B2(KEYINPUT32), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT33), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n306), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n306), .B(KEYINPUT32), .C1(new_n309), .C2(new_n305), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n300), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n299), .A2(new_n312), .A3(KEYINPUT72), .A4(new_n313), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n238), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n293), .A2(new_n222), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n322));
  OR3_X1    g121(.A1(new_n288), .A2(new_n227), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n224), .A2(new_n325), .A3(new_n288), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n327), .B(KEYINPUT82), .Z(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n288), .A2(new_n227), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n321), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n322), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n319), .B2(new_n318), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n336), .B2(new_n330), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT6), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n338), .A2(KEYINPUT85), .A3(new_n343), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT84), .B1(new_n338), .B2(new_n343), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n331), .A2(new_n337), .A3(new_n353), .A4(new_n342), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n345), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n347), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n273), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n273), .A2(new_n225), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n208), .B(new_n358), .C1(new_n359), .C2(new_n357), .ZN(new_n360));
  INV_X1    g159(.A(new_n358), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n357), .B1(new_n273), .B2(new_n225), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n228), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  NAND4_X1  g165(.A1(new_n360), .A2(new_n363), .A3(KEYINPUT30), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n360), .A2(new_n363), .ZN(new_n370));
  INV_X1    g169(.A(new_n366), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n368), .A3(new_n367), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n363), .A3(new_n366), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n373), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(KEYINPUT78), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n317), .A2(new_n356), .A3(new_n375), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT35), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n352), .A2(new_n344), .A3(new_n345), .A4(new_n354), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n347), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n379), .B1(new_n369), .B2(new_n373), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n314), .A2(new_n299), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n314), .A2(KEYINPUT76), .A3(new_n299), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n291), .A2(new_n298), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n312), .A2(new_n396), .A3(new_n313), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT75), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n238), .A2(KEYINPUT35), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n383), .B1(new_n390), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n320), .A2(new_n326), .A3(new_n323), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n328), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n403), .A2(KEYINPUT39), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n318), .A2(new_n329), .A3(new_n332), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(KEYINPUT39), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n342), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT40), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n404), .A2(KEYINPUT40), .A3(new_n342), .A4(new_n406), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n409), .A2(new_n344), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n387), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n238), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n370), .A2(KEYINPUT37), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n360), .A2(new_n363), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n371), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT38), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n417), .A2(KEYINPUT38), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(KEYINPUT86), .A3(KEYINPUT38), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n376), .A4(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n413), .B1(new_n423), .B2(new_n385), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n381), .A2(new_n375), .ZN(new_n425));
  INV_X1    g224(.A(new_n355), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n342), .B1(new_n331), .B2(new_n337), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(new_n348), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n346), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n238), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n315), .A2(KEYINPUT36), .A3(new_n316), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT36), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n395), .A2(new_n398), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n424), .A2(new_n430), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n401), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G229gat), .A2(G233gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(KEYINPUT13), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n234), .A2(G15gat), .ZN(new_n439));
  INV_X1    g238(.A(G15gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G22gat), .ZN(new_n441));
  INV_X1    g240(.A(G1gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT92), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G22gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT92), .A3(new_n443), .ZN(new_n448));
  INV_X1    g247(.A(G8gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n444), .A2(KEYINPUT91), .A3(G8gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n447), .A2(G1gat), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G43gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G50gat), .ZN(new_n460));
  INV_X1    g259(.A(G50gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G43gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT15), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT14), .ZN(new_n464));
  INV_X1    g263(.A(G29gat), .ZN(new_n465));
  INV_X1    g264(.A(G36gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g268(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT88), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT89), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n463), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n459), .B2(G50gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n461), .A2(KEYINPUT90), .A3(G43gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n460), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT15), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n472), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n475), .A2(new_n463), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n458), .B1(new_n476), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n476), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n450), .B(new_n454), .C1(new_n456), .C2(new_n455), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n438), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT17), .B1(new_n485), .B2(new_n476), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n472), .B1(new_n470), .B2(KEYINPUT88), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n467), .A2(new_n468), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n475), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n463), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n497), .A2(new_n463), .A3(new_n475), .A4(new_n483), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n458), .B1(new_n491), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n487), .A2(new_n488), .ZN(new_n502));
  INV_X1    g301(.A(new_n436), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n490), .B1(new_n504), .B2(KEYINPUT18), .ZN(new_n505));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G197gat), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT11), .B(G169gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT12), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n505), .B(new_n510), .C1(KEYINPUT18), .C2(new_n504), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n504), .B2(KEYINPUT18), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n491), .A2(new_n500), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n488), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n486), .A3(new_n436), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT93), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(new_n505), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n510), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n519), .A2(KEYINPUT94), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT94), .B1(new_n519), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT95), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n525), .A2(KEYINPUT97), .A3(new_n526), .A4(new_n529), .ZN(new_n533));
  INV_X1    g332(.A(G57gat), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n534), .A2(G64gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(G64gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n524), .ZN(new_n537));
  OAI22_X1  g336(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(KEYINPUT9), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(KEYINPUT98), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT98), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G57gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n542), .A3(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n536), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n543), .A2(KEYINPUT99), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT99), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT100), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n537), .B1(KEYINPUT9), .B2(new_n527), .ZN(new_n548));
  NOR4_X1   g347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n543), .A2(new_n544), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT99), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT98), .B(G57gat), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n536), .B1(new_n553), .B2(G64gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT99), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT100), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n539), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G127gat), .ZN(new_n562));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n488), .B1(new_n557), .B2(new_n558), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT101), .Z(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n214), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n563), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n562), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT102), .Z(new_n577));
  XOR2_X1   g376(.A(G134gat), .B(G162gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT103), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT103), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT8), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n588), .A2(KEYINPUT104), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT104), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n582), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n594), .B(new_n582), .C1(new_n591), .C2(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n514), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n598), .B2(new_n487), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n580), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n599), .B2(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT105), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT105), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n608), .B(new_n603), .C1(new_n599), .C2(new_n601), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT106), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT106), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n605), .A2(new_n607), .A3(new_n612), .A4(new_n609), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n602), .A2(new_n604), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n606), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n580), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT108), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n557), .A2(new_n598), .ZN(new_n620));
  INV_X1    g419(.A(new_n548), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n554), .B2(KEYINPUT99), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n547), .B1(new_n622), .B2(new_n545), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n552), .A2(KEYINPUT100), .A3(new_n555), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n625), .A2(new_n539), .A3(new_n597), .A4(new_n596), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n619), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AOI211_X1 g429(.A(KEYINPUT108), .B(new_n628), .C1(new_n620), .C2(new_n626), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n626), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n598), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n639), .A2(KEYINPUT10), .A3(new_n625), .A4(new_n539), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n628), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n629), .B1(new_n638), .B2(new_n640), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT107), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n636), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n630), .A2(new_n631), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n634), .B1(new_n649), .B2(new_n642), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n575), .A2(new_n618), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n435), .A2(new_n523), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n356), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n442), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n654), .A2(new_n387), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n449), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n654), .A2(new_n387), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(KEYINPUT42), .B2(new_n660), .ZN(G1325gat));
  NAND2_X1  g461(.A1(new_n395), .A2(new_n398), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n440), .B1(new_n654), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT109), .Z(new_n665));
  AOI211_X1 g464(.A(new_n440), .B(new_n654), .C1(new_n431), .C2(new_n433), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(G1326gat));
  INV_X1    g466(.A(new_n238), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n654), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n618), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n401), .B2(new_n434), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n570), .A2(new_n574), .ZN(new_n674));
  INV_X1    g473(.A(new_n523), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n674), .A2(new_n675), .A3(new_n652), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n465), .A3(new_n429), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT45), .ZN(new_n680));
  AND4_X1   g479(.A1(new_n424), .A2(new_n431), .A3(new_n430), .A4(new_n433), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n385), .A2(new_n387), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT87), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n685), .A2(new_n686), .B1(KEYINPUT35), .B2(new_n382), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n618), .B1(new_n681), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n673), .A2(KEYINPUT44), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n676), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n356), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n680), .A2(new_n694), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n692), .A2(new_n412), .A3(new_n676), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n692), .A2(KEYINPUT110), .A3(new_n412), .A4(new_n676), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(G36gat), .A3(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n677), .A2(G36gat), .A3(new_n387), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1329gat));
  OAI21_X1  g502(.A(new_n459), .B1(new_n677), .B2(new_n663), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n433), .A2(new_n431), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G43gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n693), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT47), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n709), .B(new_n704), .C1(new_n693), .C2(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1330gat));
  NAND4_X1  g510(.A1(new_n690), .A2(new_n238), .A3(new_n691), .A4(new_n676), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n677), .A2(G50gat), .A3(new_n668), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT48), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n714), .B1(new_n712), .B2(G50gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n719), .A2(KEYINPUT111), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n721), .ZN(G1331gat));
  NAND4_X1  g521(.A1(new_n674), .A2(new_n675), .A3(new_n672), .A4(new_n652), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n401), .B2(new_n434), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n429), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(new_n553), .Z(G1332gat));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n412), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT49), .B(G64gat), .Z(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(G1333gat));
  NAND2_X1  g529(.A1(new_n724), .A2(new_n705), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n663), .A2(G71gat), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n731), .A2(G71gat), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n724), .A2(new_n238), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n674), .A2(new_n523), .A3(new_n651), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n692), .A2(new_n429), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n584), .A2(new_n586), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n692), .A2(KEYINPUT112), .A3(new_n429), .A4(new_n737), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n674), .A2(new_n523), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n673), .A2(KEYINPUT51), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT51), .B1(new_n673), .B2(new_n744), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT113), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(KEYINPUT113), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n356), .A2(new_n741), .A3(new_n651), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n743), .A2(new_n750), .ZN(G1336gat));
  NOR3_X1   g550(.A1(new_n387), .A2(new_n651), .A3(G92gat), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n747), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n690), .A2(new_n412), .A3(new_n691), .A4(new_n737), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n435), .A2(new_n618), .A3(new_n744), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n673), .A2(KEYINPUT51), .A3(new_n744), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI22_X1  g561(.A1(G92gat), .A2(new_n754), .B1(new_n762), .B2(new_n752), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n753), .A2(new_n757), .B1(new_n763), .B2(new_n756), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n692), .A2(new_n705), .A3(new_n737), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G99gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n747), .A2(new_n748), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n663), .A2(G99gat), .A3(new_n651), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT114), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n767), .B2(new_n769), .ZN(G1338gat));
  NOR3_X1   g569(.A1(new_n668), .A2(G106gat), .A3(new_n651), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n745), .B2(new_n746), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT115), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n762), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n690), .A2(new_n238), .A3(new_n691), .A4(new_n737), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT53), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n747), .A2(new_n748), .A3(new_n771), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT53), .B1(new_n776), .B2(G106gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT107), .B1(new_n641), .B2(new_n628), .ZN(new_n785));
  AOI211_X1 g584(.A(new_n643), .B(new_n629), .C1(new_n638), .C2(new_n640), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n638), .A2(new_n640), .A3(new_n629), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT54), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n634), .B1(new_n645), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT55), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n647), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n787), .A2(KEYINPUT54), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n644), .A2(new_n794), .A3(new_n646), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT55), .B1(new_n795), .B2(new_n791), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n436), .B1(new_n515), .B2(new_n486), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n489), .A2(new_n486), .A3(new_n438), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n509), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n511), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(new_n618), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n650), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n801), .B1(new_n804), .B2(new_n647), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n797), .B2(new_n523), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT116), .B(new_n803), .C1(new_n806), .C2(new_n618), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  INV_X1    g608(.A(new_n791), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n789), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g610(.A(new_n809), .B(new_n634), .C1(new_n645), .C2(new_n790), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n785), .A2(new_n786), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n795), .A2(new_n812), .B1(new_n813), .B2(new_n636), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n523), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n805), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n618), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND4_X1   g616(.A1(new_n618), .A2(new_n811), .A3(new_n814), .A4(new_n802), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n808), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n807), .A2(new_n819), .A3(new_n575), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n674), .A2(new_n675), .A3(new_n672), .A4(new_n651), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n238), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n356), .A2(new_n412), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n663), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n822), .A2(KEYINPUT117), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n822), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n523), .A2(G113gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n356), .B1(new_n820), .B2(new_n821), .ZN(new_n832));
  INV_X1    g631(.A(new_n317), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n412), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n675), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(G113gat), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n784), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  OAI221_X1 g637(.A(KEYINPUT118), .B1(G113gat), .B2(new_n836), .C1(new_n829), .C2(new_n830), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1340gat));
  INV_X1    g639(.A(new_n835), .ZN(new_n841));
  AOI21_X1  g640(.A(G120gat), .B1(new_n841), .B2(new_n652), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n652), .A2(G120gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n828), .B2(new_n843), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n829), .B2(new_n575), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n282), .A3(new_n674), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  OAI21_X1  g646(.A(G134gat), .B1(new_n829), .B2(new_n672), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n835), .A2(new_n285), .A3(new_n672), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT56), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(G141gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n705), .A2(new_n824), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n238), .A2(KEYINPUT57), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n575), .B1(new_n817), .B2(new_n818), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n821), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n820), .A2(new_n821), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n858), .B2(new_n238), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n859), .B2(KEYINPUT119), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n668), .B1(new_n820), .B2(new_n821), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(KEYINPUT57), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n854), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n852), .B1(new_n864), .B2(new_n523), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n705), .A2(new_n668), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n832), .A2(new_n387), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n523), .A2(new_n852), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT58), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n859), .A2(KEYINPUT119), .ZN(new_n873));
  INV_X1    g672(.A(new_n857), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n863), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n523), .A3(new_n853), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G141gat), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n870), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n872), .A2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n881), .A3(new_n652), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT59), .B(new_n881), .C1(new_n864), .C2(new_n652), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n855), .B1(new_n820), .B2(new_n821), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n821), .A2(new_n856), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n238), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n652), .B(new_n853), .C1(new_n885), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n884), .B1(new_n888), .B2(G148gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n882), .B1(new_n883), .B2(new_n889), .ZN(G1345gat));
  AOI21_X1  g689(.A(G155gat), .B1(new_n867), .B2(new_n674), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n575), .A2(new_n214), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT121), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n864), .B2(new_n893), .ZN(G1346gat));
  NAND3_X1  g693(.A1(new_n867), .A2(new_n215), .A3(new_n618), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n864), .A2(new_n618), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n215), .ZN(G1347gat));
  AOI21_X1  g696(.A(new_n429), .B1(new_n820), .B2(new_n821), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n898), .A2(new_n317), .A3(new_n412), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n250), .A3(new_n523), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n356), .A2(new_n412), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n663), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n822), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n675), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(KEYINPUT122), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(KEYINPUT122), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n899), .A2(new_n251), .A3(new_n652), .ZN(new_n908));
  OAI21_X1  g707(.A(G176gat), .B1(new_n903), .B2(new_n651), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1349gat));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n899), .A2(new_n242), .A3(new_n674), .ZN(new_n913));
  OAI21_X1  g712(.A(G183gat), .B1(new_n903), .B2(new_n575), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n915), .B(new_n916), .Z(G1350gat));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n243), .A3(new_n618), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n822), .A2(new_n618), .A3(new_n902), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  AND4_X1   g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(G190gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n243), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n920), .A2(new_n923), .B1(new_n919), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n918), .B1(new_n922), .B2(new_n924), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n866), .A2(new_n412), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT125), .Z(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n898), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n523), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n885), .A2(new_n887), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n705), .A3(new_n901), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(G197gat), .A3(new_n523), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n930), .A2(new_n934), .ZN(G1352gat));
  INV_X1    g734(.A(G204gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n652), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  OR3_X1    g738(.A1(new_n928), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n932), .A2(new_n652), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n928), .B2(new_n937), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n203), .A3(new_n674), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n705), .A2(new_n901), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n674), .B(new_n946), .C1(new_n885), .C2(new_n887), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(G211gat), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  NAND3_X1  g754(.A1(new_n929), .A2(new_n204), .A3(new_n618), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n932), .A2(new_n618), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n958), .B2(new_n204), .ZN(G1355gat));
endmodule


