

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731;

  AND2_X1 U368 ( .A1(n650), .A2(n612), .ZN(n420) );
  NOR2_X1 U369 ( .A1(n642), .A2(n639), .ZN(n658) );
  INV_X1 U370 ( .A(n540), .ZN(n639) );
  BUF_X1 U371 ( .A(G128), .Z(n355) );
  INV_X2 U372 ( .A(G953), .ZN(n722) );
  NOR2_X2 U373 ( .A1(n577), .A2(n574), .ZN(n595) );
  XNOR2_X2 U374 ( .A(n560), .B(KEYINPUT6), .ZN(n594) );
  NOR2_X2 U375 ( .A1(n667), .A2(n668), .ZN(n599) );
  XNOR2_X2 U376 ( .A(n532), .B(n459), .ZN(n668) );
  OR2_X1 U377 ( .A1(n622), .A2(G902), .ZN(n361) );
  INV_X1 U378 ( .A(KEYINPUT95), .ZN(n442) );
  AND2_X1 U379 ( .A1(n357), .A2(n356), .ZN(n615) );
  NOR2_X1 U380 ( .A1(n675), .A2(n575), .ZN(n576) );
  XNOR2_X1 U381 ( .A(n408), .B(KEYINPUT32), .ZN(n729) );
  XNOR2_X1 U382 ( .A(n544), .B(KEYINPUT80), .ZN(n634) );
  INV_X1 U383 ( .A(n534), .ZN(n387) );
  NAND2_X1 U384 ( .A1(n523), .A2(n660), .ZN(n542) );
  XNOR2_X1 U385 ( .A(n498), .B(n432), .ZN(n375) );
  OR2_X2 U386 ( .A1(n704), .A2(G902), .ZN(n475) );
  AND2_X1 U387 ( .A1(n394), .A2(n392), .ZN(n551) );
  AND2_X1 U388 ( .A1(n395), .A2(n637), .ZN(n394) );
  NOR2_X1 U389 ( .A1(n634), .A2(n550), .ZN(n393) );
  XNOR2_X1 U390 ( .A(G146), .B(G125), .ZN(n469) );
  XNOR2_X1 U391 ( .A(n375), .B(n448), .ZN(n717) );
  XNOR2_X1 U392 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U393 ( .A(G134), .ZN(n446) );
  XNOR2_X1 U394 ( .A(G137), .B(G131), .ZN(n447) );
  INV_X1 U395 ( .A(n539), .ZN(n546) );
  XNOR2_X1 U396 ( .A(KEYINPUT69), .B(G469), .ZN(n389) );
  OR2_X1 U397 ( .A1(n695), .A2(G902), .ZN(n390) );
  XNOR2_X1 U398 ( .A(n422), .B(G110), .ZN(n450) );
  XNOR2_X1 U399 ( .A(n427), .B(n426), .ZN(n487) );
  XOR2_X1 U400 ( .A(G113), .B(G116), .Z(n426) );
  XNOR2_X1 U401 ( .A(n717), .B(n449), .ZN(n486) );
  INV_X1 U402 ( .A(G146), .ZN(n449) );
  NOR2_X1 U403 ( .A1(n534), .A2(n365), .ZN(n364) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(KEYINPUT104), .Z(n504) );
  XNOR2_X1 U405 ( .A(G113), .B(G131), .ZN(n503) );
  XNOR2_X1 U406 ( .A(n368), .B(G122), .ZN(n502) );
  INV_X1 U407 ( .A(KEYINPUT11), .ZN(n368) );
  NAND2_X1 U408 ( .A1(G234), .A2(G237), .ZN(n476) );
  XOR2_X1 U409 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n477) );
  XNOR2_X1 U410 ( .A(n554), .B(n353), .ZN(n377) );
  XNOR2_X1 U411 ( .A(n542), .B(n541), .ZN(n567) );
  XNOR2_X1 U412 ( .A(n486), .B(n415), .ZN(n622) );
  XNOR2_X1 U413 ( .A(n487), .B(n349), .ZN(n415) );
  XOR2_X1 U414 ( .A(KEYINPUT5), .B(KEYINPUT101), .Z(n485) );
  XNOR2_X1 U415 ( .A(n406), .B(n707), .ZN(n441) );
  XNOR2_X1 U416 ( .A(n369), .B(n438), .ZN(n406) );
  XNOR2_X1 U417 ( .A(n375), .B(n437), .ZN(n369) );
  XNOR2_X1 U418 ( .A(n401), .B(n530), .ZN(n400) );
  OR2_X1 U419 ( .A1(n410), .A2(KEYINPUT39), .ZN(n384) );
  NAND2_X1 U420 ( .A1(n386), .A2(n388), .ZN(n385) );
  XNOR2_X1 U421 ( .A(n573), .B(KEYINPUT22), .ZN(n577) );
  XNOR2_X1 U422 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U423 ( .A(n414), .B(n413), .ZN(n412) );
  INV_X1 U424 ( .A(KEYINPUT30), .ZN(n413) );
  AND2_X1 U425 ( .A1(n604), .A2(n411), .ZN(n410) );
  INV_X1 U426 ( .A(n533), .ZN(n411) );
  XNOR2_X1 U427 ( .A(n403), .B(n402), .ZN(n704) );
  XNOR2_X1 U428 ( .A(n468), .B(n350), .ZN(n402) );
  XNOR2_X1 U429 ( .A(n467), .B(n716), .ZN(n403) );
  XNOR2_X1 U430 ( .A(n486), .B(n456), .ZN(n695) );
  XNOR2_X1 U431 ( .A(n453), .B(n452), .ZN(n455) );
  NOR2_X1 U432 ( .A1(G952), .A2(n722), .ZN(n706) );
  INV_X1 U433 ( .A(n658), .ZN(n397) );
  NOR2_X1 U434 ( .A1(G953), .A2(G237), .ZN(n507) );
  OR2_X1 U435 ( .A1(n671), .A2(n533), .ZN(n483) );
  OR2_X1 U436 ( .A1(G237), .A2(G902), .ZN(n518) );
  XNOR2_X1 U437 ( .A(n405), .B(G119), .ZN(n425) );
  INV_X1 U438 ( .A(KEYINPUT70), .ZN(n405) );
  XOR2_X1 U439 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n509) );
  XNOR2_X1 U440 ( .A(G143), .B(G104), .ZN(n501) );
  XNOR2_X1 U441 ( .A(G902), .B(KEYINPUT15), .ZN(n460) );
  XNOR2_X1 U442 ( .A(n431), .B(KEYINPUT64), .ZN(n432) );
  INV_X1 U443 ( .A(KEYINPUT4), .ZN(n431) );
  XNOR2_X1 U444 ( .A(KEYINPUT17), .B(KEYINPUT78), .ZN(n436) );
  XOR2_X1 U445 ( .A(KEYINPUT93), .B(KEYINPUT18), .Z(n434) );
  INV_X1 U446 ( .A(n410), .ZN(n365) );
  XNOR2_X1 U447 ( .A(n407), .B(KEYINPUT0), .ZN(n572) );
  NOR2_X1 U448 ( .A1(n567), .A2(n568), .ZN(n407) );
  NOR2_X1 U449 ( .A1(n648), .A2(n359), .ZN(n358) );
  INV_X1 U450 ( .A(n727), .ZN(n359) );
  XNOR2_X1 U451 ( .A(G140), .B(KEYINPUT10), .ZN(n470) );
  XNOR2_X1 U452 ( .A(G119), .B(G137), .ZN(n464) );
  XOR2_X1 U453 ( .A(G110), .B(n355), .Z(n465) );
  XNOR2_X1 U454 ( .A(KEYINPUT106), .B(KEYINPUT9), .ZN(n490) );
  XOR2_X1 U455 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n491) );
  XNOR2_X1 U456 ( .A(G116), .B(G134), .ZN(n488) );
  XOR2_X1 U457 ( .A(G122), .B(G107), .Z(n489) );
  XNOR2_X1 U458 ( .A(G101), .B(n450), .ZN(n453) );
  INV_X1 U459 ( .A(KEYINPUT77), .ZN(n451) );
  XNOR2_X1 U460 ( .A(n378), .B(KEYINPUT87), .ZN(n611) );
  AND2_X1 U461 ( .A1(n559), .A2(n379), .ZN(n376) );
  XNOR2_X1 U462 ( .A(n528), .B(KEYINPUT41), .ZN(n687) );
  XNOR2_X1 U463 ( .A(n588), .B(KEYINPUT35), .ZN(n590) );
  NOR2_X1 U464 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U465 ( .A(KEYINPUT34), .ZN(n584) );
  XNOR2_X1 U466 ( .A(n515), .B(n514), .ZN(n539) );
  OR2_X1 U467 ( .A1(n543), .A2(n567), .ZN(n544) );
  XNOR2_X1 U468 ( .A(n600), .B(KEYINPUT98), .ZN(n602) );
  XNOR2_X1 U469 ( .A(n423), .B(n450), .ZN(n428) );
  XNOR2_X1 U470 ( .A(n421), .B(KEYINPUT16), .ZN(n423) );
  NAND2_X1 U471 ( .A1(n382), .A2(n639), .ZN(n381) );
  NOR2_X1 U472 ( .A1(n668), .A2(n526), .ZN(n646) );
  AND2_X1 U473 ( .A1(n374), .A2(n373), .ZN(n525) );
  INV_X1 U474 ( .A(n542), .ZN(n373) );
  OR2_X1 U475 ( .A1(n577), .A2(n409), .ZN(n408) );
  NAND2_X1 U476 ( .A1(n348), .A2(n347), .ZN(n409) );
  NAND2_X1 U477 ( .A1(n410), .A2(n412), .ZN(n547) );
  INV_X1 U478 ( .A(KEYINPUT63), .ZN(n391) );
  XNOR2_X1 U479 ( .A(n702), .B(n360), .ZN(n705) );
  XNOR2_X1 U480 ( .A(n704), .B(n703), .ZN(n360) );
  XNOR2_X1 U481 ( .A(n695), .B(n354), .ZN(n417) );
  INV_X1 U482 ( .A(n706), .ZN(n356) );
  INV_X1 U483 ( .A(KEYINPUT53), .ZN(n366) );
  AND2_X1 U484 ( .A1(n412), .A2(KEYINPUT39), .ZN(n346) );
  NOR2_X1 U485 ( .A1(n668), .A2(n671), .ZN(n347) );
  XOR2_X1 U486 ( .A(KEYINPUT79), .B(n594), .Z(n348) );
  XOR2_X1 U487 ( .A(n485), .B(n484), .Z(n349) );
  INV_X1 U488 ( .A(n648), .ZN(n379) );
  XNOR2_X1 U489 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n350) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n351) );
  INV_X1 U491 ( .A(KEYINPUT39), .ZN(n388) );
  XNOR2_X1 U492 ( .A(KEYINPUT45), .B(KEYINPUT86), .ZN(n352) );
  XOR2_X1 U493 ( .A(KEYINPUT48), .B(KEYINPUT88), .Z(n353) );
  XNOR2_X1 U494 ( .A(n428), .B(n487), .ZN(n707) );
  XOR2_X1 U495 ( .A(n697), .B(n696), .Z(n354) );
  XNOR2_X1 U496 ( .A(n372), .B(n351), .ZN(n357) );
  NOR2_X1 U497 ( .A1(n731), .A2(n730), .ZN(n536) );
  XNOR2_X1 U498 ( .A(n531), .B(KEYINPUT42), .ZN(n731) );
  NAND2_X1 U499 ( .A1(n377), .A2(n358), .ZN(n720) );
  NAND2_X1 U500 ( .A1(n419), .A2(G210), .ZN(n372) );
  NOR2_X1 U501 ( .A1(n381), .A2(n383), .ZN(n535) );
  XNOR2_X2 U502 ( .A(n361), .B(G472), .ZN(n560) );
  XNOR2_X1 U503 ( .A(n362), .B(n391), .ZN(G57) );
  NOR2_X2 U504 ( .A1(n625), .A2(n706), .ZN(n362) );
  XNOR2_X1 U505 ( .A(n363), .B(n621), .ZN(G60) );
  NOR2_X2 U506 ( .A1(n620), .A2(n706), .ZN(n363) );
  NAND2_X1 U507 ( .A1(n346), .A2(n364), .ZN(n382) );
  NOR2_X2 U508 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U509 ( .A(n367), .B(n366), .ZN(G75) );
  NAND2_X1 U510 ( .A1(n694), .A2(n693), .ZN(n367) );
  INV_X1 U511 ( .A(n572), .ZN(n600) );
  XNOR2_X1 U512 ( .A(n585), .B(n584), .ZN(n587) );
  NAND2_X1 U513 ( .A1(n633), .A2(n729), .ZN(n580) );
  NAND2_X1 U514 ( .A1(n576), .A2(n598), .ZN(n633) );
  NAND2_X1 U515 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U516 ( .A1(n371), .A2(n370), .ZN(n614) );
  INV_X1 U517 ( .A(KEYINPUT2), .ZN(n370) );
  NAND2_X1 U518 ( .A1(n404), .A2(n613), .ZN(n371) );
  INV_X1 U519 ( .A(n614), .ZN(n649) );
  XNOR2_X1 U520 ( .A(n524), .B(KEYINPUT112), .ZN(n374) );
  NAND2_X1 U521 ( .A1(n377), .A2(n376), .ZN(n378) );
  NAND2_X1 U522 ( .A1(n387), .A2(n412), .ZN(n386) );
  NAND2_X1 U523 ( .A1(n380), .A2(n382), .ZN(n555) );
  INV_X1 U524 ( .A(n383), .ZN(n380) );
  NAND2_X1 U525 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X2 U526 ( .A(n390), .B(n389), .ZN(n532) );
  XNOR2_X1 U527 ( .A(n393), .B(KEYINPUT73), .ZN(n392) );
  NAND2_X1 U528 ( .A1(n396), .A2(KEYINPUT47), .ZN(n395) );
  NAND2_X1 U529 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U530 ( .A(n634), .ZN(n398) );
  NAND2_X1 U531 ( .A1(n400), .A2(n399), .ZN(n543) );
  INV_X1 U532 ( .A(n532), .ZN(n399) );
  NAND2_X1 U533 ( .A1(n529), .A2(n560), .ZN(n401) );
  NOR2_X2 U534 ( .A1(n483), .A2(n569), .ZN(n529) );
  NAND2_X1 U535 ( .A1(n404), .A2(n720), .ZN(n652) );
  NAND2_X1 U536 ( .A1(n404), .A2(n722), .ZN(n713) );
  NAND2_X1 U537 ( .A1(n611), .A2(n404), .ZN(n650) );
  XNOR2_X2 U538 ( .A(n610), .B(n352), .ZN(n404) );
  NAND2_X1 U539 ( .A1(n560), .A2(n660), .ZN(n414) );
  NOR2_X1 U540 ( .A1(n416), .A2(n706), .ZN(G54) );
  XNOR2_X1 U541 ( .A(n418), .B(n417), .ZN(n416) );
  NAND2_X1 U542 ( .A1(n419), .A2(G469), .ZN(n418) );
  AND2_X2 U543 ( .A1(n420), .A2(n614), .ZN(n419) );
  XNOR2_X1 U544 ( .A(n578), .B(KEYINPUT91), .ZN(n579) );
  NOR2_X1 U545 ( .A1(n594), .A2(n581), .ZN(n583) );
  XNOR2_X1 U546 ( .A(n451), .B(G140), .ZN(n452) );
  INV_X1 U547 ( .A(KEYINPUT65), .ZN(n429) );
  INV_X1 U548 ( .A(KEYINPUT1), .ZN(n457) );
  XNOR2_X1 U549 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U550 ( .A(n617), .B(KEYINPUT59), .ZN(n618) );
  XNOR2_X1 U551 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n621) );
  XOR2_X1 U552 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n440) );
  XOR2_X1 U553 ( .A(KEYINPUT71), .B(G122), .Z(n421) );
  XNOR2_X1 U554 ( .A(G104), .B(G107), .ZN(n422) );
  XNOR2_X1 U555 ( .A(KEYINPUT3), .B(G101), .ZN(n424) );
  XNOR2_X1 U556 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X2 U557 ( .A(G143), .B(G128), .ZN(n430) );
  XNOR2_X2 U558 ( .A(n430), .B(n429), .ZN(n498) );
  NAND2_X1 U559 ( .A1(G224), .A2(n722), .ZN(n433) );
  XNOR2_X1 U560 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U561 ( .A(n435), .B(KEYINPUT94), .Z(n438) );
  XNOR2_X1 U562 ( .A(n436), .B(n469), .ZN(n437) );
  XNOR2_X1 U563 ( .A(n441), .B(KEYINPUT83), .ZN(n439) );
  INV_X1 U564 ( .A(n460), .ZN(n612) );
  NOR2_X2 U565 ( .A1(n612), .A2(n441), .ZN(n445) );
  NAND2_X1 U566 ( .A1(G210), .A2(n518), .ZN(n443) );
  XNOR2_X2 U567 ( .A(n445), .B(n444), .ZN(n523) );
  NAND2_X1 U568 ( .A1(G227), .A2(n722), .ZN(n454) );
  XNOR2_X1 U569 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U570 ( .A(KEYINPUT66), .ZN(n458) );
  INV_X1 U571 ( .A(n668), .ZN(n574) );
  XOR2_X1 U572 ( .A(KEYINPUT21), .B(KEYINPUT100), .Z(n463) );
  NAND2_X1 U573 ( .A1(G234), .A2(n460), .ZN(n461) );
  XNOR2_X1 U574 ( .A(KEYINPUT20), .B(n461), .ZN(n471) );
  NAND2_X1 U575 ( .A1(n471), .A2(G221), .ZN(n462) );
  XOR2_X1 U576 ( .A(n463), .B(n462), .Z(n569) );
  XNOR2_X1 U577 ( .A(n465), .B(n464), .ZN(n468) );
  NAND2_X1 U578 ( .A1(G234), .A2(n722), .ZN(n466) );
  XOR2_X1 U579 ( .A(KEYINPUT8), .B(n466), .Z(n494) );
  NAND2_X1 U580 ( .A1(n494), .A2(G221), .ZN(n467) );
  XOR2_X1 U581 ( .A(n470), .B(n469), .Z(n716) );
  NAND2_X1 U582 ( .A1(n471), .A2(G217), .ZN(n472) );
  XNOR2_X1 U583 ( .A(n472), .B(KEYINPUT25), .ZN(n473) );
  XNOR2_X1 U584 ( .A(KEYINPUT99), .B(n473), .ZN(n474) );
  XNOR2_X2 U585 ( .A(n475), .B(n474), .ZN(n671) );
  XNOR2_X1 U586 ( .A(n477), .B(n476), .ZN(n479) );
  NAND2_X1 U587 ( .A1(G902), .A2(n479), .ZN(n564) );
  NOR2_X1 U588 ( .A1(G900), .A2(n564), .ZN(n478) );
  NAND2_X1 U589 ( .A1(G953), .A2(n478), .ZN(n481) );
  NAND2_X1 U590 ( .A1(G952), .A2(n479), .ZN(n686) );
  NOR2_X1 U591 ( .A1(G953), .A2(n686), .ZN(n480) );
  XOR2_X1 U592 ( .A(KEYINPUT96), .B(n480), .Z(n561) );
  NAND2_X1 U593 ( .A1(n481), .A2(n561), .ZN(n482) );
  XNOR2_X1 U594 ( .A(KEYINPUT81), .B(n482), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n507), .A2(G210), .ZN(n484) );
  XNOR2_X1 U596 ( .A(KEYINPUT107), .B(G478), .ZN(n500) );
  XNOR2_X1 U597 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U599 ( .A(n493), .B(n492), .Z(n496) );
  NAND2_X1 U600 ( .A1(G217), .A2(n494), .ZN(n495) );
  XNOR2_X1 U601 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n498), .B(n497), .ZN(n698) );
  NOR2_X1 U603 ( .A1(G902), .A2(n698), .ZN(n499) );
  XOR2_X1 U604 ( .A(n500), .B(n499), .Z(n545) );
  INV_X1 U605 ( .A(n716), .ZN(n513) );
  XNOR2_X1 U606 ( .A(n502), .B(n501), .ZN(n506) );
  XNOR2_X1 U607 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U608 ( .A(n506), .B(n505), .ZN(n511) );
  NAND2_X1 U609 ( .A1(G214), .A2(n507), .ZN(n508) );
  XNOR2_X1 U610 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U611 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U612 ( .A(n512), .B(n513), .Z(n616) );
  NOR2_X1 U613 ( .A1(G902), .A2(n616), .ZN(n515) );
  XNOR2_X1 U614 ( .A(KEYINPUT13), .B(G475), .ZN(n514) );
  NAND2_X1 U615 ( .A1(n545), .A2(n539), .ZN(n540) );
  NOR2_X1 U616 ( .A1(n594), .A2(n540), .ZN(n516) );
  NAND2_X1 U617 ( .A1(n529), .A2(n516), .ZN(n517) );
  XNOR2_X1 U618 ( .A(KEYINPUT109), .B(n517), .ZN(n524) );
  NAND2_X1 U619 ( .A1(G214), .A2(n518), .ZN(n660) );
  NAND2_X1 U620 ( .A1(n524), .A2(n660), .ZN(n519) );
  NOR2_X1 U621 ( .A1(n574), .A2(n519), .ZN(n521) );
  XNOR2_X1 U622 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n521), .B(n520), .ZN(n522) );
  NOR2_X1 U624 ( .A1(n523), .A2(n522), .ZN(n648) );
  XOR2_X1 U625 ( .A(KEYINPUT36), .B(n525), .Z(n526) );
  INV_X1 U626 ( .A(KEYINPUT46), .ZN(n537) );
  XOR2_X1 U627 ( .A(KEYINPUT38), .B(KEYINPUT76), .Z(n527) );
  XOR2_X1 U628 ( .A(n523), .B(n527), .Z(n534) );
  NAND2_X1 U629 ( .A1(n387), .A2(n660), .ZN(n657) );
  NAND2_X1 U630 ( .A1(n546), .A2(n545), .ZN(n662) );
  NOR2_X1 U631 ( .A1(n657), .A2(n662), .ZN(n528) );
  XNOR2_X1 U632 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n530) );
  NOR2_X1 U633 ( .A1(n687), .A2(n543), .ZN(n531) );
  INV_X1 U634 ( .A(n569), .ZN(n672) );
  NAND2_X1 U635 ( .A1(n672), .A2(n671), .ZN(n667) );
  NOR2_X1 U636 ( .A1(n532), .A2(n667), .ZN(n604) );
  XNOR2_X1 U637 ( .A(n535), .B(KEYINPUT40), .ZN(n730) );
  XNOR2_X1 U638 ( .A(n537), .B(n536), .ZN(n538) );
  NOR2_X1 U639 ( .A1(n646), .A2(n538), .ZN(n553) );
  NOR2_X1 U640 ( .A1(n539), .A2(n545), .ZN(n642) );
  XNOR2_X1 U641 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n541) );
  OR2_X1 U642 ( .A1(n546), .A2(n545), .ZN(n586) );
  NOR2_X1 U643 ( .A1(n547), .A2(n586), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n523), .A2(n548), .ZN(n637) );
  NOR2_X1 U645 ( .A1(KEYINPUT47), .A2(n658), .ZN(n549) );
  XOR2_X1 U646 ( .A(KEYINPUT74), .B(n549), .Z(n550) );
  XNOR2_X1 U647 ( .A(n551), .B(KEYINPUT72), .ZN(n552) );
  NAND2_X1 U648 ( .A1(n553), .A2(n552), .ZN(n554) );
  INV_X1 U649 ( .A(n642), .ZN(n556) );
  NOR2_X1 U650 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U651 ( .A(n557), .B(KEYINPUT113), .ZN(n727) );
  NAND2_X1 U652 ( .A1(KEYINPUT2), .A2(n727), .ZN(n558) );
  XOR2_X1 U653 ( .A(KEYINPUT82), .B(n558), .Z(n559) );
  INV_X1 U654 ( .A(n671), .ZN(n598) );
  BUF_X1 U655 ( .A(n560), .Z(n675) );
  INV_X1 U656 ( .A(n561), .ZN(n566) );
  NOR2_X1 U657 ( .A1(G898), .A2(n722), .ZN(n562) );
  XOR2_X1 U658 ( .A(KEYINPUT97), .B(n562), .Z(n708) );
  INV_X1 U659 ( .A(n708), .ZN(n563) );
  NOR2_X1 U660 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U661 ( .A1(n566), .A2(n565), .ZN(n568) );
  OR2_X1 U662 ( .A1(n569), .A2(n662), .ZN(n570) );
  XOR2_X1 U663 ( .A(KEYINPUT108), .B(n570), .Z(n571) );
  NAND2_X1 U664 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U665 ( .A(n595), .ZN(n575) );
  INV_X1 U666 ( .A(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n591), .A2(KEYINPUT90), .ZN(n578) );
  XNOR2_X1 U668 ( .A(n580), .B(n579), .ZN(n589) );
  INV_X1 U669 ( .A(n599), .ZN(n581) );
  XNOR2_X1 U670 ( .A(KEYINPUT92), .B(KEYINPUT33), .ZN(n582) );
  XNOR2_X1 U671 ( .A(n583), .B(n582), .ZN(n688) );
  NOR2_X1 U672 ( .A1(n688), .A2(n602), .ZN(n585) );
  NAND2_X1 U673 ( .A1(n589), .A2(n590), .ZN(n593) );
  INV_X1 U674 ( .A(n590), .ZN(n728) );
  NAND2_X1 U675 ( .A1(n728), .A2(n591), .ZN(n592) );
  NAND2_X1 U676 ( .A1(n593), .A2(n592), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U678 ( .A(KEYINPUT89), .B(n596), .Z(n597) );
  NOR2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n626) );
  NAND2_X1 U680 ( .A1(n675), .A2(n599), .ZN(n678) );
  NOR2_X1 U681 ( .A1(n600), .A2(n678), .ZN(n601) );
  XOR2_X1 U682 ( .A(KEYINPUT31), .B(n601), .Z(n643) );
  INV_X1 U683 ( .A(n602), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U685 ( .A1(n675), .A2(n605), .ZN(n628) );
  NOR2_X1 U686 ( .A1(n643), .A2(n628), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n658), .A2(n606), .ZN(n607) );
  NOR2_X1 U688 ( .A1(n626), .A2(n607), .ZN(n608) );
  INV_X1 U689 ( .A(n720), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U691 ( .A1(n419), .A2(G475), .ZN(n619) );
  INV_X1 U692 ( .A(n616), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n419), .A2(G472), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT62), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(n625) );
  XOR2_X1 U697 ( .A(G101), .B(n626), .Z(G3) );
  NAND2_X1 U698 ( .A1(n628), .A2(n639), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n627), .B(G104), .ZN(G6) );
  XNOR2_X1 U700 ( .A(G107), .B(KEYINPUT27), .ZN(n632) );
  XOR2_X1 U701 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n630) );
  NAND2_X1 U702 ( .A1(n628), .A2(n642), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n632), .B(n631), .ZN(G9) );
  XNOR2_X1 U705 ( .A(n633), .B(G110), .ZN(G12) );
  XOR2_X1 U706 ( .A(n355), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U707 ( .A1(n642), .A2(n398), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G30) );
  XNOR2_X1 U709 ( .A(G143), .B(n637), .ZN(G45) );
  NAND2_X1 U710 ( .A1(n398), .A2(n639), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n638), .B(G146), .ZN(G48) );
  XOR2_X1 U712 ( .A(G113), .B(KEYINPUT115), .Z(n641) );
  NAND2_X1 U713 ( .A1(n643), .A2(n639), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G15) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(KEYINPUT116), .ZN(n645) );
  XNOR2_X1 U717 ( .A(G116), .B(n645), .ZN(G18) );
  XNOR2_X1 U718 ( .A(G125), .B(n646), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U720 ( .A(G140), .B(n648), .Z(G42) );
  NAND2_X1 U721 ( .A1(n649), .A2(KEYINPUT84), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n655) );
  NOR2_X1 U723 ( .A1(KEYINPUT2), .A2(n652), .ZN(n653) );
  NOR2_X1 U724 ( .A1(KEYINPUT84), .A2(n653), .ZN(n654) );
  XNOR2_X1 U725 ( .A(KEYINPUT85), .B(n656), .ZN(n694) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT119), .B(n659), .Z(n665) );
  NOR2_X1 U728 ( .A1(n387), .A2(n660), .ZN(n661) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U730 ( .A(KEYINPUT118), .B(n663), .ZN(n664) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n688), .A2(n666), .ZN(n683) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT50), .B(n669), .Z(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT117), .ZN(n677) );
  NOR2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U737 ( .A(KEYINPUT49), .B(n673), .Z(n674) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U741 ( .A(KEYINPUT51), .B(n680), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n681), .A2(n687), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U744 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n691) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U747 ( .A(KEYINPUT120), .B(n689), .ZN(n690) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n692) );
  AND2_X1 U749 ( .A1(n692), .A2(n722), .ZN(n693) );
  XOR2_X1 U750 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n697) );
  XNOR2_X1 U751 ( .A(KEYINPUT122), .B(KEYINPUT121), .ZN(n696) );
  XOR2_X1 U752 ( .A(n698), .B(KEYINPUT123), .Z(n700) );
  NAND2_X1 U753 ( .A1(n419), .A2(G478), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n706), .A2(n701), .ZN(G63) );
  XOR2_X1 U756 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n703) );
  NAND2_X1 U757 ( .A1(n419), .A2(G217), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(G66) );
  NOR2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n715) );
  NAND2_X1 U760 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n709), .B(KEYINPUT61), .ZN(n710) );
  XNOR2_X1 U762 ( .A(KEYINPUT126), .B(n710), .ZN(n711) );
  NAND2_X1 U763 ( .A1(G898), .A2(n711), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U765 ( .A(n715), .B(n714), .ZN(G69) );
  XOR2_X1 U766 ( .A(n717), .B(n716), .Z(n721) );
  XNOR2_X1 U767 ( .A(n721), .B(G227), .ZN(n718) );
  NOR2_X1 U768 ( .A1(n722), .A2(n718), .ZN(n719) );
  NAND2_X1 U769 ( .A1(n719), .A2(G900), .ZN(n725) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U773 ( .A(n726), .B(KEYINPUT127), .ZN(G72) );
  XNOR2_X1 U774 ( .A(G134), .B(n727), .ZN(G36) );
  XOR2_X1 U775 ( .A(n728), .B(G122), .Z(G24) );
  XNOR2_X1 U776 ( .A(G119), .B(n729), .ZN(G21) );
  XOR2_X1 U777 ( .A(n730), .B(G131), .Z(G33) );
  XOR2_X1 U778 ( .A(G137), .B(n731), .Z(G39) );
endmodule

