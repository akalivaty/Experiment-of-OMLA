

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U326 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n362) );
  XNOR2_X1 U327 ( .A(n363), .B(n362), .ZN(n381) );
  XNOR2_X1 U328 ( .A(n331), .B(KEYINPUT72), .ZN(n332) );
  XNOR2_X1 U329 ( .A(n413), .B(n332), .ZN(n336) );
  XNOR2_X1 U330 ( .A(n340), .B(n432), .ZN(n341) );
  XNOR2_X1 U331 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n391) );
  XNOR2_X1 U332 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U333 ( .A(n392), .B(n391), .ZN(n546) );
  XNOR2_X1 U334 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n295) );
  XNOR2_X1 U337 ( .A(G134GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U339 ( .A(n296), .B(G99GAT), .Z(n298) );
  XOR2_X1 U340 ( .A(G113GAT), .B(KEYINPUT0), .Z(n417) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(n417), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n304) );
  XOR2_X1 U343 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n300) );
  XNOR2_X1 U344 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n401) );
  XOR2_X1 U346 ( .A(n401), .B(G183GAT), .Z(n302) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n312) );
  XOR2_X1 U350 ( .A(G71GAT), .B(KEYINPUT20), .Z(n306) );
  XNOR2_X1 U351 ( .A(KEYINPUT85), .B(KEYINPUT66), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U353 ( .A(G176GAT), .B(G120GAT), .Z(n308) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n558) );
  INV_X1 U358 ( .A(n558), .ZN(n561) );
  XOR2_X1 U359 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n314) );
  XNOR2_X1 U360 ( .A(G106GAT), .B(G92GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n329) );
  XNOR2_X1 U362 ( .A(G99GAT), .B(G85GAT), .ZN(n343) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n315), .B(KEYINPUT78), .ZN(n397) );
  XNOR2_X1 U365 ( .A(n343), .B(n397), .ZN(n317) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U368 ( .A(G162GAT), .B(n318), .ZN(n323) );
  XOR2_X1 U369 ( .A(G29GAT), .B(G134GAT), .Z(n412) );
  XOR2_X1 U370 ( .A(KEYINPUT77), .B(n412), .Z(n320) );
  XOR2_X1 U371 ( .A(G50GAT), .B(KEYINPUT74), .Z(n433) );
  XNOR2_X1 U372 ( .A(G218GAT), .B(n433), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U374 ( .A(n321), .B(KEYINPUT10), .Z(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U376 ( .A(n324), .B(KEYINPUT76), .Z(n327) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n325), .B(KEYINPUT7), .ZN(n357) );
  XNOR2_X1 U379 ( .A(n357), .B(KEYINPUT9), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n384) );
  NAND2_X1 U382 ( .A1(n561), .A2(n384), .ZN(n447) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(G148GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n330), .B(G57GAT), .ZN(n413) );
  AND2_X1 U385 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XOR2_X1 U386 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n334) );
  XNOR2_X1 U387 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U389 ( .A(n336), .B(n335), .Z(n342) );
  XNOR2_X1 U390 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n337), .B(KEYINPUT13), .ZN(n367) );
  XOR2_X1 U392 ( .A(G64GAT), .B(G92GAT), .Z(n339) );
  XNOR2_X1 U393 ( .A(G176GAT), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n393) );
  XNOR2_X1 U395 ( .A(n367), .B(n393), .ZN(n340) );
  XOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .Z(n432) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n578) );
  XNOR2_X1 U398 ( .A(KEYINPUT41), .B(n578), .ZN(n505) );
  XOR2_X1 U399 ( .A(G1GAT), .B(G141GAT), .Z(n346) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(G197GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U402 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n348) );
  XNOR2_X1 U403 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n361) );
  XOR2_X1 U406 ( .A(G15GAT), .B(G22GAT), .Z(n377) );
  XOR2_X1 U407 ( .A(G113GAT), .B(G36GAT), .Z(n352) );
  XNOR2_X1 U408 ( .A(G29GAT), .B(G50GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(n377), .B(n353), .Z(n355) );
  NAND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(n356), .B(KEYINPUT30), .Z(n359) );
  XNOR2_X1 U414 ( .A(n357), .B(KEYINPUT70), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n573) );
  NAND2_X1 U417 ( .A1(n505), .A2(n573), .ZN(n363) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n369) );
  XOR2_X1 U419 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n365) );
  XNOR2_X1 U420 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U424 ( .A(G8GAT), .B(G183GAT), .Z(n394) );
  XOR2_X1 U425 ( .A(G1GAT), .B(G127GAT), .Z(n410) );
  XOR2_X1 U426 ( .A(n394), .B(n410), .Z(n371) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U429 ( .A(n373), .B(n372), .Z(n379) );
  XOR2_X1 U430 ( .A(G57GAT), .B(G78GAT), .Z(n375) );
  XNOR2_X1 U431 ( .A(G155GAT), .B(G211GAT), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n488) );
  INV_X1 U435 ( .A(n488), .ZN(n583) );
  OR2_X1 U436 ( .A1(n384), .A2(n583), .ZN(n380) );
  NOR2_X1 U437 ( .A1(n381), .A2(n380), .ZN(n383) );
  INV_X1 U438 ( .A(KEYINPUT47), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n390) );
  XNOR2_X1 U440 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n586) );
  NOR2_X1 U442 ( .A1(n488), .A2(n586), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n386), .B(KEYINPUT45), .ZN(n387) );
  NAND2_X1 U444 ( .A1(n387), .A2(n578), .ZN(n388) );
  NOR2_X1 U445 ( .A1(n388), .A2(n573), .ZN(n389) );
  NOR2_X1 U446 ( .A1(n390), .A2(n389), .ZN(n392) );
  XOR2_X1 U447 ( .A(n394), .B(n393), .Z(n396) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U450 ( .A(n398), .B(n397), .Z(n403) );
  XOR2_X1 U451 ( .A(G211GAT), .B(KEYINPUT21), .Z(n400) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n441) );
  XNOR2_X1 U454 ( .A(n401), .B(n441), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n523) );
  XNOR2_X1 U456 ( .A(n523), .B(KEYINPUT121), .ZN(n404) );
  NOR2_X1 U457 ( .A1(n546), .A2(n404), .ZN(n405) );
  XNOR2_X1 U458 ( .A(n405), .B(KEYINPUT54), .ZN(n427) );
  XOR2_X1 U459 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n407) );
  XNOR2_X1 U460 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n421) );
  XOR2_X1 U462 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n409) );
  XNOR2_X1 U463 ( .A(G85GAT), .B(KEYINPUT1), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U465 ( .A(n411), .B(n410), .Z(n419) );
  XOR2_X1 U466 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U471 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U472 ( .A(KEYINPUT86), .B(KEYINPUT3), .Z(n423) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(G155GAT), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U475 ( .A(G162GAT), .B(KEYINPUT2), .Z(n424) );
  XNOR2_X1 U476 ( .A(n425), .B(n424), .ZN(n429) );
  XNOR2_X1 U477 ( .A(n426), .B(n429), .ZN(n465) );
  XNOR2_X1 U478 ( .A(KEYINPUT92), .B(n465), .ZN(n475) );
  NAND2_X1 U479 ( .A1(n427), .A2(n475), .ZN(n428) );
  XNOR2_X1 U480 ( .A(n428), .B(KEYINPUT65), .ZN(n571) );
  INV_X1 U481 ( .A(n429), .ZN(n445) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n431) );
  XNOR2_X1 U483 ( .A(G22GAT), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n437) );
  XOR2_X1 U485 ( .A(G204GAT), .B(KEYINPUT88), .Z(n435) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U488 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U491 ( .A(n440), .B(KEYINPUT87), .Z(n443) );
  XNOR2_X1 U492 ( .A(n441), .B(KEYINPUT24), .ZN(n442) );
  XNOR2_X1 U493 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U494 ( .A(n445), .B(n444), .ZN(n458) );
  AND2_X1 U495 ( .A1(n571), .A2(n458), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n446), .B(KEYINPUT55), .ZN(n562) );
  OR2_X1 U497 ( .A1(n447), .A2(n562), .ZN(n451) );
  XOR2_X1 U498 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n449) );
  INV_X1 U499 ( .A(G190GAT), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n453) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n453), .B(n452), .ZN(n477) );
  NAND2_X1 U503 ( .A1(n573), .A2(n578), .ZN(n492) );
  INV_X1 U504 ( .A(n475), .ZN(n521) );
  XNOR2_X1 U505 ( .A(n523), .B(KEYINPUT27), .ZN(n457) );
  NAND2_X1 U506 ( .A1(n521), .A2(n457), .ZN(n549) );
  XNOR2_X1 U507 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(n458), .ZN(n527) );
  NOR2_X1 U509 ( .A1(n549), .A2(n527), .ZN(n532) );
  NAND2_X1 U510 ( .A1(n558), .A2(n532), .ZN(n468) );
  NOR2_X1 U511 ( .A1(n561), .A2(n458), .ZN(n456) );
  XNOR2_X1 U512 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n455) );
  XOR2_X1 U513 ( .A(n456), .B(n455), .Z(n572) );
  NAND2_X1 U514 ( .A1(n457), .A2(n572), .ZN(n464) );
  XNOR2_X1 U515 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n462) );
  NAND2_X1 U516 ( .A1(n561), .A2(n523), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT95), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n487) );
  NOR2_X1 U523 ( .A1(n488), .A2(n384), .ZN(n471) );
  XOR2_X1 U524 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT82), .B(n469), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n487), .A2(n472), .ZN(n473) );
  XNOR2_X1 U528 ( .A(KEYINPUT96), .B(n473), .ZN(n508) );
  NOR2_X1 U529 ( .A1(n492), .A2(n508), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n474), .B(KEYINPUT97), .ZN(n482) );
  NOR2_X1 U531 ( .A1(n475), .A2(n482), .ZN(n476) );
  XOR2_X1 U532 ( .A(n477), .B(n476), .Z(G1324GAT) );
  INV_X1 U533 ( .A(n523), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n478), .A2(n482), .ZN(n479) );
  XOR2_X1 U535 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U536 ( .A1(n558), .A2(n482), .ZN(n481) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  INV_X1 U539 ( .A(n527), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n483), .A2(n482), .ZN(n485) );
  XNOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U545 ( .A1(n488), .A2(n487), .ZN(n489) );
  NOR2_X1 U546 ( .A1(n586), .A2(n489), .ZN(n491) );
  XNOR2_X1 U547 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n520) );
  NOR2_X1 U549 ( .A1(n492), .A2(n520), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n493), .B(KEYINPUT38), .ZN(n502) );
  NAND2_X1 U551 ( .A1(n502), .A2(n521), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n496), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(G36GAT), .B(KEYINPUT105), .Z(n498) );
  NAND2_X1 U555 ( .A1(n523), .A2(n502), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n500) );
  NAND2_X1 U558 ( .A1(n502), .A2(n561), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U560 ( .A(G43GAT), .B(n501), .Z(G1330GAT) );
  XOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U562 ( .A1(n502), .A2(n527), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n510) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT108), .ZN(n560) );
  INV_X1 U566 ( .A(n573), .ZN(n506) );
  NAND2_X1 U567 ( .A1(n560), .A2(n506), .ZN(n507) );
  XOR2_X1 U568 ( .A(KEYINPUT109), .B(n507), .Z(n519) );
  NOR2_X1 U569 ( .A1(n508), .A2(n519), .ZN(n516) );
  NAND2_X1 U570 ( .A1(n516), .A2(n521), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n511), .Z(G1332GAT) );
  XOR2_X1 U573 ( .A(G64GAT), .B(KEYINPUT111), .Z(n513) );
  NAND2_X1 U574 ( .A1(n516), .A2(n523), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n561), .A2(n516), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT112), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U580 ( .A1(n516), .A2(n527), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n520), .A2(n519), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n528), .A2(n521), .ZN(n522) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n528), .A2(n523), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT113), .Z(n526) );
  NAND2_X1 U588 ( .A1(n528), .A2(n561), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n530) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U593 ( .A(G106GAT), .B(n531), .Z(G1339GAT) );
  NAND2_X1 U594 ( .A1(n532), .A2(n561), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n546), .A2(n533), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n542), .A2(n573), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(KEYINPUT116), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n537) );
  NAND2_X1 U600 ( .A1(n542), .A2(n560), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U604 ( .A1(n542), .A2(n583), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U608 ( .A1(n542), .A2(n384), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U610 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  INV_X1 U611 ( .A(n546), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n547), .A2(n572), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n573), .A2(n555), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U617 ( .A1(n555), .A2(n505), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n583), .A2(n555), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n384), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n562), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n568), .A2(n573), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  OR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n565) );
  XOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT123), .Z(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n583), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .Z(n575) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n585) );
  INV_X1 U639 ( .A(n585), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n580) );
  OR2_X1 U645 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

