

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  INV_X1 U325 ( .A(n461), .ZN(n529) );
  NOR2_X1 U326 ( .A1(n486), .A2(n580), .ZN(n386) );
  XNOR2_X2 U327 ( .A(n454), .B(KEYINPUT119), .ZN(n565) );
  XOR2_X1 U328 ( .A(n340), .B(n339), .Z(n293) );
  XNOR2_X1 U329 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n398) );
  XNOR2_X1 U330 ( .A(n399), .B(n398), .ZN(n526) );
  XOR2_X1 U331 ( .A(n346), .B(n345), .Z(n576) );
  XOR2_X1 U332 ( .A(n465), .B(KEYINPUT28), .Z(n532) );
  XNOR2_X1 U333 ( .A(n455), .B(G190GAT), .ZN(n456) );
  XNOR2_X1 U334 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n295) );
  XNOR2_X1 U336 ( .A(G197GAT), .B(G204GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(G211GAT), .B(n296), .Z(n401) );
  XOR2_X1 U339 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n298) );
  XNOR2_X1 U340 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n401), .B(n299), .ZN(n313) );
  XOR2_X1 U343 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n301) );
  XNOR2_X1 U344 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U346 ( .A(KEYINPUT3), .B(n302), .Z(n430) );
  XOR2_X1 U347 ( .A(G78GAT), .B(G148GAT), .Z(n333) );
  XOR2_X1 U348 ( .A(G22GAT), .B(G155GAT), .Z(n369) );
  XOR2_X1 U349 ( .A(n333), .B(n369), .Z(n304) );
  XNOR2_X1 U350 ( .A(G218GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U352 ( .A(n430), .B(n305), .Z(n307) );
  NAND2_X1 U353 ( .A1(G228GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(n308), .B(KEYINPUT23), .Z(n311) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n309), .B(G162GAT), .ZN(n354) );
  XNOR2_X1 U358 ( .A(n354), .B(KEYINPUT88), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n465) );
  XOR2_X1 U361 ( .A(KEYINPUT66), .B(KEYINPUT7), .Z(n315) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G29GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U364 ( .A(KEYINPUT8), .B(n316), .Z(n358) );
  XOR2_X1 U365 ( .A(G197GAT), .B(KEYINPUT68), .Z(n318) );
  XNOR2_X1 U366 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n358), .B(n319), .ZN(n330) );
  XOR2_X1 U369 ( .A(G169GAT), .B(G8GAT), .Z(n408) );
  XOR2_X1 U370 ( .A(KEYINPUT29), .B(G22GAT), .Z(n321) );
  XNOR2_X1 U371 ( .A(G36GAT), .B(G50GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U373 ( .A(n408), .B(n322), .Z(n324) );
  NAND2_X1 U374 ( .A1(G229GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U376 ( .A(n325), .B(G113GAT), .Z(n328) );
  XNOR2_X1 U377 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n326), .B(G15GAT), .ZN(n372) );
  XNOR2_X1 U379 ( .A(n372), .B(G141GAT), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U381 ( .A(n330), .B(n329), .Z(n570) );
  INV_X1 U382 ( .A(n570), .ZN(n556) );
  XOR2_X1 U383 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n332) );
  XNOR2_X1 U384 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n346) );
  XOR2_X1 U386 ( .A(G176GAT), .B(G64GAT), .Z(n400) );
  XOR2_X1 U387 ( .A(KEYINPUT73), .B(n400), .Z(n335) );
  XNOR2_X1 U388 ( .A(G92GAT), .B(n333), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U390 ( .A(KEYINPUT13), .B(G57GAT), .Z(n373) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n336), .B(G106GAT), .ZN(n355) );
  XNOR2_X1 U393 ( .A(n373), .B(n355), .ZN(n338) );
  AND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U396 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XOR2_X1 U397 ( .A(KEYINPUT71), .B(G204GAT), .Z(n342) );
  XNOR2_X1 U398 ( .A(KEYINPUT69), .B(KEYINPUT31), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n437), .B(n343), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n293), .B(n344), .ZN(n345) );
  INV_X1 U402 ( .A(KEYINPUT78), .ZN(n364) );
  INV_X1 U403 ( .A(KEYINPUT11), .ZN(n350) );
  XOR2_X1 U404 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n348) );
  XNOR2_X1 U405 ( .A(KEYINPUT9), .B(KEYINPUT64), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n352) );
  NAND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(G134GAT), .B(KEYINPUT76), .Z(n425) );
  XNOR2_X1 U411 ( .A(n353), .B(n425), .ZN(n357) );
  XOR2_X1 U412 ( .A(n355), .B(n354), .Z(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U415 ( .A(G218GAT), .B(G92GAT), .Z(n361) );
  XNOR2_X1 U416 ( .A(G190GAT), .B(KEYINPUT77), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U418 ( .A(G36GAT), .B(n362), .Z(n404) );
  XOR2_X1 U419 ( .A(n363), .B(n404), .Z(n392) );
  XNOR2_X1 U420 ( .A(n364), .B(n392), .ZN(n540) );
  XOR2_X1 U421 ( .A(KEYINPUT36), .B(KEYINPUT100), .Z(n365) );
  XNOR2_X1 U422 ( .A(n540), .B(n365), .ZN(n486) );
  XOR2_X1 U423 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n367) );
  XNOR2_X1 U424 ( .A(G71GAT), .B(G78GAT), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U426 ( .A(n368), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U427 ( .A(G8GAT), .B(n369), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n377) );
  XOR2_X1 U429 ( .A(n373), .B(n372), .Z(n375) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U432 ( .A(n377), .B(n376), .Z(n385) );
  XOR2_X1 U433 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n379) );
  XNOR2_X1 U434 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U436 ( .A(G211GAT), .B(KEYINPUT12), .Z(n381) );
  XNOR2_X1 U437 ( .A(G183GAT), .B(G127GAT), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U440 ( .A(n385), .B(n384), .Z(n580) );
  XNOR2_X1 U441 ( .A(KEYINPUT45), .B(n386), .ZN(n387) );
  NAND2_X1 U442 ( .A1(n576), .A2(n387), .ZN(n388) );
  NOR2_X1 U443 ( .A1(n556), .A2(n388), .ZN(n397) );
  XOR2_X1 U444 ( .A(KEYINPUT109), .B(KEYINPUT47), .Z(n395) );
  INV_X1 U445 ( .A(n580), .ZN(n564) );
  XOR2_X1 U446 ( .A(KEYINPUT41), .B(n576), .Z(n500) );
  OR2_X1 U447 ( .A1(n500), .A2(n570), .ZN(n390) );
  INV_X1 U448 ( .A(KEYINPUT46), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n391) );
  NOR2_X1 U450 ( .A1(n564), .A2(n391), .ZN(n393) );
  BUF_X1 U451 ( .A(n392), .Z(n554) );
  NAND2_X1 U452 ( .A1(n393), .A2(n554), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  NOR2_X1 U454 ( .A1(n397), .A2(n396), .ZN(n399) );
  XOR2_X1 U455 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U458 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U459 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n407) );
  XNOR2_X1 U460 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n442) );
  XNOR2_X1 U462 ( .A(n408), .B(n442), .ZN(n409) );
  XOR2_X1 U463 ( .A(n410), .B(n409), .Z(n517) );
  XOR2_X1 U464 ( .A(n517), .B(KEYINPUT118), .Z(n411) );
  NOR2_X1 U465 ( .A1(n526), .A2(n411), .ZN(n412) );
  XOR2_X1 U466 ( .A(KEYINPUT54), .B(n412), .Z(n435) );
  XOR2_X1 U467 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n414) );
  XNOR2_X1 U468 ( .A(G113GAT), .B(G127GAT), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n438) );
  XOR2_X1 U470 ( .A(n438), .B(KEYINPUT94), .Z(n416) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n434) );
  XOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n418) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(G155GAT), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U476 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n420) );
  XNOR2_X1 U477 ( .A(KEYINPUT95), .B(KEYINPUT4), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n432) );
  XOR2_X1 U480 ( .A(G148GAT), .B(G57GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(G120GAT), .B(G162GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U483 ( .A(n426), .B(n425), .Z(n428) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G85GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n470) );
  INV_X1 U489 ( .A(n470), .ZN(n515) );
  NOR2_X2 U490 ( .A1(n435), .A2(n515), .ZN(n569) );
  NAND2_X1 U491 ( .A1(n465), .A2(n569), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n436), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U493 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n441), .B(KEYINPUT85), .Z(n444) );
  XNOR2_X1 U497 ( .A(n442), .B(KEYINPUT20), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n452) );
  XOR2_X1 U499 ( .A(G134GAT), .B(G99GAT), .Z(n446) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G190GAT), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT86), .B(G176GAT), .Z(n448) );
  XNOR2_X1 U503 ( .A(G169GAT), .B(G15GAT), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U505 ( .A(n450), .B(n449), .Z(n451) );
  XOR2_X1 U506 ( .A(n452), .B(n451), .Z(n461) );
  NAND2_X1 U507 ( .A1(n453), .A2(n529), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n565), .A2(n540), .ZN(n457) );
  XOR2_X1 U509 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n455) );
  NAND2_X1 U510 ( .A1(n556), .A2(n576), .ZN(n491) );
  OR2_X1 U511 ( .A1(n540), .A2(n580), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n458), .B(KEYINPUT16), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT83), .ZN(n474) );
  XNOR2_X1 U514 ( .A(n517), .B(KEYINPUT27), .ZN(n467) );
  NAND2_X1 U515 ( .A1(n515), .A2(n467), .ZN(n525) );
  NOR2_X1 U516 ( .A1(n532), .A2(n525), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n473) );
  NAND2_X1 U518 ( .A1(n529), .A2(n517), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n462), .A2(n465), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT96), .B(n463), .Z(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT25), .ZN(n469) );
  NOR2_X1 U522 ( .A1(n529), .A2(n465), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U524 ( .A1(n467), .A2(n568), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n487) );
  NAND2_X1 U528 ( .A1(n474), .A2(n487), .ZN(n501) );
  NOR2_X1 U529 ( .A1(n491), .A2(n501), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT97), .B(n475), .Z(n482) );
  NAND2_X1 U531 ( .A1(n482), .A2(n515), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(KEYINPUT34), .ZN(n477) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n517), .A2(n482), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U537 ( .A1(n482), .A2(n529), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U540 ( .A1(n482), .A2(n532), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n485) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n494) );
  NAND2_X1 U545 ( .A1(n580), .A2(n487), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT101), .B(n488), .Z(n489) );
  NOR2_X1 U547 ( .A1(n486), .A2(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n490), .ZN(n512) );
  NOR2_X1 U549 ( .A1(n512), .A2(n491), .ZN(n492) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n492), .ZN(n498) );
  NAND2_X1 U551 ( .A1(n498), .A2(n515), .ZN(n493) );
  XOR2_X1 U552 ( .A(n494), .B(n493), .Z(G1328GAT) );
  NAND2_X1 U553 ( .A1(n498), .A2(n517), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n529), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U558 ( .A1(n498), .A2(n532), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U560 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  INV_X1 U561 ( .A(n500), .ZN(n561) );
  NAND2_X1 U562 ( .A1(n570), .A2(n561), .ZN(n513) );
  NOR2_X1 U563 ( .A1(n513), .A2(n501), .ZN(n508) );
  NAND2_X1 U564 ( .A1(n515), .A2(n508), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  XOR2_X1 U566 ( .A(G64GAT), .B(KEYINPUT103), .Z(n505) );
  NAND2_X1 U567 ( .A1(n508), .A2(n517), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n529), .A2(n508), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT104), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n510) );
  NAND2_X1 U573 ( .A1(n508), .A2(n532), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U575 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT106), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n515), .A2(n522), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  XOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U581 ( .A1(n522), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n522), .A2(n529), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT108), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n522), .A2(n532), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U589 ( .A(G113GAT), .B(KEYINPUT113), .Z(n534) );
  INV_X1 U590 ( .A(KEYINPUT111), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n544) );
  NAND2_X1 U593 ( .A1(n544), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(KEYINPUT112), .B(n530), .ZN(n531) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n556), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U599 ( .A1(n541), .A2(n561), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n538) );
  NAND2_X1 U602 ( .A1(n541), .A2(n564), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n544), .A2(n568), .ZN(n553) );
  NOR2_X1 U609 ( .A1(n570), .A2(n553), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n550) );
  NOR2_X1 U615 ( .A1(n500), .A2(n553), .ZN(n549) );
  XOR2_X1 U616 ( .A(n550), .B(n549), .Z(G1345GAT) );
  NOR2_X1 U617 ( .A1(n580), .A2(n553), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NAND2_X1 U622 ( .A1(n565), .A2(n556), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n559) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(n560), .Z(n563) );
  NAND2_X1 U628 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G183GAT), .B(n567), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n582) );
  NOR2_X1 U634 ( .A1(n570), .A2(n582), .ZN(n575) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT124), .B(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n582), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n486), .A2(n582), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

