//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n471), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n477), .A2(G124), .B1(G136), .B2(new_n467), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT68), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n478), .A2(new_n481), .ZN(G162));
  NAND2_X1  g057(.A1(G126), .A2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n465), .B2(new_n466), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n467), .B2(G138), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n462), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n488), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n502), .A2(new_n503), .A3(new_n509), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n508), .A2(new_n515), .ZN(G166));
  OR2_X1    g091(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(G76), .A2(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G651), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(new_n517), .A3(new_n518), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n510), .A2(G51), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n502), .A2(G89), .A3(new_n503), .A4(new_n509), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n502), .A2(G63), .A3(G651), .A4(new_n503), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n524), .A2(KEYINPUT71), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(new_n523), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n509), .A2(G51), .A3(G543), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n528), .A2(new_n525), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n527), .A2(new_n532), .ZN(G168));
  NAND4_X1  g108(.A1(new_n502), .A2(G90), .A3(new_n503), .A4(new_n509), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n509), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n502), .A2(G64), .A3(new_n503), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n507), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n537), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(new_n510), .A2(G43), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n502), .A2(G81), .A3(new_n503), .A4(new_n509), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n504), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n545), .B1(G651), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g126(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n552));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n536), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n536), .B2(new_n556), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(new_n558), .B1(G91), .B2(new_n512), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n504), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  OAI21_X1  g141(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n512), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n510), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  AOI22_X1  g145(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n507), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n512), .A2(G86), .B1(G48), .B2(new_n510), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(G72), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G60), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n504), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n577), .A2(KEYINPUT73), .A3(G651), .ZN(new_n581));
  XOR2_X1   g156(.A(KEYINPUT74), .B(G85), .Z(new_n582));
  AOI22_X1  g157(.A1(new_n512), .A2(new_n582), .B1(G47), .B2(new_n510), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n504), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n502), .A2(G92), .A3(new_n503), .A4(new_n509), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n585), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n585), .B1(new_n594), .B2(G868), .ZN(G321));
  NOR2_X1   g171(.A1(G299), .A2(G868), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g173(.A(new_n597), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n467), .A2(G135), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT76), .Z(new_n607));
  OAI21_X1  g182(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n608));
  INV_X1    g183(.A(G111), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G2105), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n477), .B2(G123), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(G2096), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n471), .A2(new_n463), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n613), .A2(G2096), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n614), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT78), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT79), .ZN(G401));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT80), .Z(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n644), .B(new_n646), .C1(new_n642), .C2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n643), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(new_n641), .A3(new_n645), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n642), .A2(new_n648), .A3(new_n645), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1991), .B(G1996), .Z(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT83), .ZN(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT85), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n664), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n659), .A2(new_n660), .ZN(new_n670));
  MUX2_X1   g245(.A(new_n669), .B(new_n664), .S(new_n670), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n672), .B1(new_n668), .B2(new_n671), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n657), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n675), .ZN(new_n677));
  INV_X1    g252(.A(new_n657), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n678), .A3(new_n673), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n680), .B1(new_n676), .B2(new_n679), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G29), .A2(G33), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT25), .Z(new_n687));
  INV_X1    g262(.A(G139), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n468), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n471), .A2(G127), .ZN(new_n690));
  NAND2_X1  g265(.A1(G115), .A2(G2104), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n462), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n685), .B1(new_n693), .B2(G29), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G34), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT86), .B(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(G34), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G160), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G2084), .ZN(new_n703));
  AOI22_X1  g278(.A1(G2072), .A2(new_n694), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G2072), .B2(new_n694), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT31), .B(G11), .Z(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT91), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n613), .A2(new_n697), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT92), .B(KEYINPUT30), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G28), .ZN(new_n710));
  AOI21_X1  g285(.A(G29), .B1(new_n709), .B2(G28), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n707), .B(new_n708), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n703), .B2(new_n702), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT89), .B(KEYINPUT26), .ZN(new_n715));
  AND3_X1   g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n463), .A2(G105), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n467), .A2(G141), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n471), .A2(G129), .A3(G2105), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(new_n701), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(KEYINPUT90), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G29), .B2(G32), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n723), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  AOI211_X1 g301(.A(new_n705), .B(new_n713), .C1(new_n714), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(G301), .A2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G5), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n549), .B2(G16), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n732), .A2(G1961), .B1(G1341), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2090), .ZN(new_n736));
  INV_X1    g311(.A(new_n697), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G35), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n735), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n732), .A2(G1961), .B1(G1341), .B2(new_n734), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n727), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n594), .A2(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G4), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n726), .A2(new_n714), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n697), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  OAI211_X1 g326(.A(G140), .B(new_n462), .C1(new_n491), .C2(new_n492), .ZN(new_n752));
  OAI211_X1 g327(.A(G128), .B(G2105), .C1(new_n491), .C2(new_n492), .ZN(new_n753));
  INV_X1    g328(.A(G116), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G104), .C2(G2105), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n751), .B1(new_n701), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2067), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(G164), .A2(new_n697), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G27), .B2(new_n697), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n761), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n748), .A2(new_n749), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n741), .A2(new_n736), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT94), .Z(new_n768));
  NOR2_X1   g343(.A1(G16), .A2(G21), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G168), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1966), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n729), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1956), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n747), .B2(new_n746), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n744), .A2(new_n766), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n729), .A2(G22), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G166), .B2(new_n729), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G1971), .Z(new_n782));
  NOR2_X1   g357(.A1(G6), .A2(G16), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n571), .A2(new_n507), .ZN(new_n784));
  INV_X1    g359(.A(new_n573), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n783), .B1(new_n786), .B2(G16), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n729), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(G288), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n729), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n782), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n467), .A2(G131), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n462), .A2(G107), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G119), .ZN(new_n803));
  OAI221_X1 g378(.A(new_n800), .B1(new_n801), .B2(new_n802), .C1(new_n803), .C2(new_n476), .ZN(new_n804));
  MUX2_X1   g379(.A(G25), .B(new_n804), .S(new_n737), .Z(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n729), .A2(G24), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G290), .B2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n798), .A2(new_n799), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT36), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n779), .A2(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NAND2_X1  g391(.A1(new_n594), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(G80), .A2(G543), .ZN(new_n819));
  INV_X1    g394(.A(G67), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n504), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G651), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n510), .A2(G55), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n502), .A2(G93), .A3(new_n503), .A4(new_n509), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT95), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n823), .A2(KEYINPUT95), .A3(new_n824), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n549), .B(new_n822), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n822), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n548), .A2(G651), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n829), .A2(new_n543), .A3(new_n544), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n818), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n835), .A2(new_n836), .A3(G860), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n828), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n757), .B(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n715), .A2(new_n716), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n715), .A2(new_n716), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n718), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n719), .A2(new_n720), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT96), .B1(new_n484), .B2(new_n487), .ZN(new_n849));
  OAI211_X1 g424(.A(G126), .B(G2105), .C1(new_n491), .C2(new_n492), .ZN(new_n850));
  INV_X1    g425(.A(G114), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n849), .B(new_n855), .C1(new_n490), .C2(new_n494), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n757), .A2(new_n841), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n721), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n848), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n857), .B1(new_n848), .B2(new_n860), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT98), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n860), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n721), .B1(new_n859), .B2(new_n858), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n848), .A2(new_n857), .A3(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n693), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n693), .B1(new_n861), .B2(new_n862), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT99), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI211_X1 g448(.A(KEYINPUT99), .B(new_n693), .C1(new_n863), .C2(new_n869), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n617), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n693), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT98), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n871), .A2(KEYINPUT99), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n617), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n870), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n804), .B(KEYINPUT100), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n467), .A2(G142), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n462), .A2(G118), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(G130), .ZN(new_n890));
  OAI221_X1 g465(.A(new_n887), .B1(new_n888), .B2(new_n889), .C1(new_n890), .C2(new_n476), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n886), .B(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n875), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n875), .B2(new_n885), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(G162), .B(new_n700), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n612), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n892), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n873), .A2(new_n874), .A3(new_n617), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n882), .B1(new_n881), .B2(new_n884), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n875), .A2(new_n885), .A3(new_n892), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n897), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g482(.A(G868), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n828), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G305), .B(G290), .ZN(new_n910));
  XNOR2_X1  g485(.A(G166), .B(G288), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT42), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n832), .B(new_n602), .Z(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n593), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n559), .A2(new_n589), .A3(new_n592), .A4(new_n563), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT41), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n917), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(KEYINPUT101), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n922), .B1(new_n914), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n913), .B(new_n928), .Z(new_n929));
  OAI21_X1  g504(.A(new_n909), .B1(new_n929), .B2(new_n908), .ZN(G295));
  XOR2_X1   g505(.A(G295), .B(KEYINPUT102), .Z(G331));
  OR3_X1    g506(.A1(new_n537), .A2(new_n540), .A3(KEYINPUT103), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT103), .B1(new_n537), .B2(new_n540), .ZN(new_n933));
  NAND3_X1  g508(.A1(G168), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(G301), .A2(new_n527), .A3(new_n532), .A4(KEYINPUT103), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n832), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n934), .A2(new_n827), .A3(new_n831), .A4(new_n935), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n833), .A2(KEYINPUT104), .A3(new_n935), .A4(new_n934), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n923), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n910), .B(new_n911), .Z(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n921), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT105), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n946), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n912), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n943), .A2(new_n944), .A3(new_n952), .A4(new_n946), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n948), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n953), .A2(new_n951), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n920), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n915), .A2(KEYINPUT106), .A3(new_n919), .A4(new_n916), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n960), .A2(new_n918), .A3(new_n961), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n942), .A2(new_n962), .B1(new_n927), .B2(new_n945), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n912), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n958), .A2(new_n948), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n957), .A2(KEYINPUT108), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT108), .B1(new_n957), .B2(new_n966), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT43), .B1(new_n963), .B2(new_n912), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n948), .A2(new_n969), .A3(new_n951), .A4(new_n953), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT107), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n958), .A2(new_n973), .A3(new_n948), .A4(new_n969), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OAI22_X1  g550(.A1(new_n967), .A2(new_n968), .B1(KEYINPUT44), .B2(new_n975), .ZN(G397));
  XNOR2_X1  g551(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n856), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n470), .A2(new_n474), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n721), .B(G1996), .ZN(new_n987));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n757), .B(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n804), .B(new_n806), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(G290), .A2(G1986), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n856), .A2(KEYINPUT112), .A3(new_n979), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT112), .B1(new_n856), .B2(new_n979), .ZN(new_n997));
  NAND2_X1  g572(.A1(G160), .A2(G40), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G305), .A2(G1981), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n784), .A2(new_n785), .A3(G1981), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1004), .A3(KEYINPUT49), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n1006));
  INV_X1    g581(.A(G1981), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n572), .B2(new_n573), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(new_n1008), .B2(new_n1003), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1001), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1012), .A2(G1976), .A3(G288), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1001), .B1(new_n1013), .B2(new_n1003), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1001), .B1(new_n1015), .B2(G288), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI22_X1  g593(.A1(new_n1016), .A2(new_n1018), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1016), .A2(KEYINPUT52), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n856), .A2(new_n979), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n856), .A2(KEYINPUT112), .A3(new_n979), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1028), .A2(KEYINPUT113), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n996), .A2(new_n997), .A3(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n495), .A2(new_n979), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(new_n1029), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1031), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT114), .B(G2090), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(new_n982), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n977), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n856), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n982), .A3(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT110), .B(G1971), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1025), .B(G8), .C1(new_n1039), .C2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1014), .B1(new_n1022), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT50), .B1(new_n996), .B2(new_n997), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n998), .B1(new_n1035), .B2(new_n1029), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1052), .A2(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1024), .B1(new_n1053), .B2(new_n1000), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1021), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n982), .A2(new_n703), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n996), .B2(new_n997), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1034), .B2(new_n977), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n495), .A2(KEYINPUT115), .A3(new_n979), .A4(new_n978), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1064), .A3(new_n982), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n771), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(G8), .B(G168), .C1(new_n1058), .C2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1048), .B1(new_n1055), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1048), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1024), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(new_n1046), .A3(new_n1072), .A4(new_n1021), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1047), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1042), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1956), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1051), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(G299), .B(KEYINPUT57), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1956), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1083), .B2(new_n1077), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(KEYINPUT61), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1028), .A2(new_n982), .A3(new_n1030), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT116), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1028), .A2(new_n1089), .A3(new_n982), .A4(new_n1030), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT58), .B(G1341), .Z(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1042), .A2(G1996), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1086), .B1(new_n1094), .B2(new_n549), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT59), .B(new_n830), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1085), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT120), .B(new_n1080), .C1(new_n1083), .C2(new_n1077), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT120), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1084), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1037), .A2(new_n982), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT117), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1037), .A2(new_n1106), .A3(new_n982), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n747), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n988), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n593), .A4(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1110), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n594), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT60), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1103), .B(new_n1111), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n593), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1084), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1116), .B(new_n1082), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1082), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT118), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1115), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  INV_X1    g698(.A(G1961), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1105), .A2(new_n1124), .A3(new_n1107), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1042), .B2(G2078), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1041), .A2(new_n982), .ZN(new_n1128));
  NOR4_X1   g703(.A1(new_n1128), .A2(new_n980), .A3(new_n1126), .A4(G2078), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT123), .Z(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1123), .B1(new_n1131), .B2(G171), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1065), .A2(new_n1126), .A3(G2078), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1133), .A2(new_n1127), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1125), .A3(G301), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1055), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(G168), .A3(new_n1066), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n1139));
  AND2_X1   g714(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(G8), .B(G286), .C1(new_n1058), .C2(new_n1067), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT51), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n1148), .A3(new_n1142), .A4(new_n1141), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1131), .A2(G171), .ZN(new_n1151));
  AOI21_X1  g726(.A(G301), .B1(new_n1134), .B2(new_n1125), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1123), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1136), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1074), .B1(new_n1122), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1150), .B2(KEYINPUT62), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n1158));
  AOI211_X1 g733(.A(KEYINPUT124), .B(new_n1158), .C1(new_n1145), .C2(new_n1149), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1145), .A2(new_n1158), .A3(new_n1149), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1054), .A2(new_n1152), .A3(new_n1046), .A4(new_n1021), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n995), .B1(new_n1155), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n806), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n804), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n991), .B2(new_n983), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(G2067), .B2(new_n757), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1169), .A2(new_n1170), .A3(new_n983), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1172), .A2(KEYINPUT126), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(KEYINPUT126), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n983), .A2(G1996), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT46), .Z(new_n1176));
  OAI21_X1  g751(.A(new_n984), .B1(new_n721), .B2(new_n990), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT47), .Z(new_n1179));
  NOR2_X1   g754(.A1(new_n986), .A2(new_n983), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1180), .A2(KEYINPUT48), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1180), .A2(KEYINPUT48), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n983), .B1(new_n991), .B2(new_n992), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NOR4_X1   g759(.A1(new_n1173), .A2(new_n1174), .A3(new_n1179), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1164), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g761(.A(new_n639), .ZN(new_n1188));
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  NOR3_X1   g763(.A1(new_n1188), .A2(new_n1189), .A3(G227), .ZN(new_n1190));
  INV_X1    g764(.A(new_n1190), .ZN(new_n1191));
  INV_X1    g765(.A(new_n683), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1192), .B2(new_n681), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n902), .A2(new_n897), .A3(new_n903), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1194), .A2(new_n951), .ZN(new_n1195));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1195), .B2(new_n904), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n1197));
  NOR3_X1   g771(.A1(new_n975), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  OAI21_X1  g772(.A(new_n1190), .B1(new_n682), .B2(new_n683), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n1199), .B1(new_n898), .B2(new_n905), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n1201));
  AOI21_X1  g775(.A(KEYINPUT127), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n1198), .A2(new_n1202), .ZN(G308));
  OAI21_X1  g777(.A(new_n1197), .B1(new_n975), .B2(new_n1196), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n1200), .A2(KEYINPUT127), .A3(new_n1201), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1205), .ZN(G225));
endmodule


