

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733;

  XNOR2_X1 U380 ( .A(G113), .B(G104), .ZN(n432) );
  XNOR2_X1 U381 ( .A(n432), .B(G122), .ZN(n510) );
  INV_X1 U382 ( .A(G953), .ZN(n688) );
  OR2_X1 U383 ( .A1(n532), .A2(n531), .ZN(n386) );
  AND2_X4 U384 ( .A1(n412), .A2(n411), .ZN(n701) );
  AND2_X2 U385 ( .A1(n681), .A2(n619), .ZN(n411) );
  XNOR2_X2 U386 ( .A(n382), .B(KEYINPUT3), .ZN(n381) );
  INV_X2 U387 ( .A(KEYINPUT70), .ZN(n382) );
  XNOR2_X2 U388 ( .A(n386), .B(n385), .ZN(n730) );
  NAND2_X1 U389 ( .A1(n397), .A2(n396), .ZN(n681) );
  AND2_X1 U390 ( .A1(n552), .A2(n551), .ZN(n553) );
  INV_X2 U391 ( .A(n581), .ZN(n613) );
  XNOR2_X1 U392 ( .A(n459), .B(n426), .ZN(n489) );
  XNOR2_X1 U393 ( .A(G146), .B(n719), .ZN(n485) );
  XOR2_X1 U394 ( .A(G131), .B(G134), .Z(n719) );
  XOR2_X1 U395 ( .A(KEYINPUT73), .B(KEYINPUT16), .Z(n433) );
  XNOR2_X1 U396 ( .A(n613), .B(KEYINPUT38), .ZN(n662) );
  XOR2_X2 U397 ( .A(G143), .B(G128), .Z(n497) );
  XNOR2_X1 U398 ( .A(KEYINPUT71), .B(G110), .ZN(n426) );
  NAND2_X1 U399 ( .A1(n701), .A2(G472), .ZN(n408) );
  NOR2_X1 U400 ( .A1(n731), .A2(n732), .ZN(n373) );
  NOR2_X1 U401 ( .A1(n631), .A2(n641), .ZN(n594) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n512) );
  AND2_X1 U403 ( .A1(n404), .A2(n403), .ZN(n617) );
  INV_X1 U404 ( .A(n644), .ZN(n403) );
  XNOR2_X1 U405 ( .A(KEYINPUT93), .B(KEYINPUT45), .ZN(n555) );
  XNOR2_X1 U406 ( .A(n496), .B(n360), .ZN(n374) );
  XOR2_X1 U407 ( .A(G116), .B(G107), .Z(n500) );
  XNOR2_X1 U408 ( .A(n706), .B(n410), .ZN(n409) );
  XNOR2_X1 U409 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U410 ( .A(n491), .B(KEYINPUT33), .ZN(n687) );
  XNOR2_X1 U411 ( .A(n576), .B(KEYINPUT41), .ZN(n659) );
  XNOR2_X1 U412 ( .A(n391), .B(KEYINPUT39), .ZN(n614) );
  INV_X1 U413 ( .A(n662), .ZN(n413) );
  OR2_X1 U414 ( .A1(n589), .A2(n663), .ZN(n609) );
  NOR2_X1 U415 ( .A1(n526), .A2(n525), .ZN(n528) );
  INV_X1 U416 ( .A(KEYINPUT28), .ZN(n378) );
  XNOR2_X1 U417 ( .A(n375), .B(KEYINPUT111), .ZN(n503) );
  OR2_X1 U418 ( .A1(n699), .A2(G902), .ZN(n375) );
  XNOR2_X1 U419 ( .A(n478), .B(n477), .ZN(n479) );
  OR2_X1 U420 ( .A1(n532), .A2(n646), .ZN(n384) );
  AND2_X1 U421 ( .A1(n729), .A2(KEYINPUT65), .ZN(n537) );
  XNOR2_X1 U422 ( .A(G146), .B(G125), .ZN(n464) );
  XNOR2_X1 U423 ( .A(n373), .B(KEYINPUT46), .ZN(n608) );
  INV_X1 U424 ( .A(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U425 ( .A(G143), .B(G131), .ZN(n504) );
  AND2_X1 U426 ( .A1(G224), .A2(n688), .ZN(n428) );
  NAND2_X1 U427 ( .A1(G234), .A2(G237), .ZN(n442) );
  XOR2_X1 U428 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n443) );
  XNOR2_X1 U429 ( .A(n372), .B(KEYINPUT116), .ZN(n668) );
  NOR2_X1 U430 ( .A1(n662), .A2(n663), .ZN(n372) );
  OR2_X1 U431 ( .A1(n694), .A2(G902), .ZN(n419) );
  AND2_X1 U432 ( .A1(n570), .A2(n363), .ZN(n647) );
  XNOR2_X1 U433 ( .A(G113), .B(G116), .ZN(n453) );
  XOR2_X1 U434 ( .A(KEYINPUT105), .B(G137), .Z(n454) );
  XOR2_X1 U435 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n452) );
  XNOR2_X1 U436 ( .A(G128), .B(G119), .ZN(n466) );
  XNOR2_X1 U437 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  XNOR2_X1 U438 ( .A(G104), .B(G107), .ZN(n483) );
  XOR2_X1 U439 ( .A(G137), .B(G140), .Z(n487) );
  AND2_X1 U440 ( .A1(G227), .A2(n688), .ZN(n421) );
  AND2_X1 U441 ( .A1(n617), .A2(n361), .ZN(n396) );
  XNOR2_X1 U442 ( .A(KEYINPUT84), .B(n492), .ZN(n493) );
  AND2_X1 U443 ( .A1(n392), .A2(n365), .ZN(n582) );
  XNOR2_X1 U444 ( .A(n563), .B(KEYINPUT30), .ZN(n564) );
  XNOR2_X1 U445 ( .A(n499), .B(n374), .ZN(n502) );
  XNOR2_X1 U446 ( .A(n579), .B(n578), .ZN(n731) );
  NOR2_X1 U447 ( .A1(n609), .A2(n590), .ZN(n591) );
  INV_X1 U448 ( .A(KEYINPUT32), .ZN(n385) );
  NAND2_X1 U449 ( .A1(n649), .A2(n651), .ZN(n383) );
  INV_X1 U450 ( .A(n384), .ZN(n548) );
  NAND2_X1 U451 ( .A1(n407), .A2(n692), .ZN(n406) );
  XNOR2_X1 U452 ( .A(n408), .B(n368), .ZN(n407) );
  INV_X1 U453 ( .A(KEYINPUT60), .ZN(n399) );
  NAND2_X1 U454 ( .A1(n401), .A2(n692), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n402), .B(n367), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n695) );
  XNOR2_X1 U457 ( .A(n694), .B(n693), .ZN(n394) );
  NAND2_X1 U458 ( .A1(n701), .A2(G469), .ZN(n395) );
  NAND2_X1 U459 ( .A1(n388), .A2(n692), .ZN(n387) );
  XNOR2_X1 U460 ( .A(n389), .B(n370), .ZN(n388) );
  INV_X1 U461 ( .A(KEYINPUT53), .ZN(n414) );
  NOR2_X1 U462 ( .A1(n686), .A2(n366), .ZN(n416) );
  XOR2_X1 U463 ( .A(KEYINPUT68), .B(G469), .Z(n359) );
  XNOR2_X1 U464 ( .A(KEYINPUT9), .B(KEYINPUT110), .ZN(n360) );
  XOR2_X1 U465 ( .A(KEYINPUT86), .B(n616), .Z(n361) );
  XOR2_X1 U466 ( .A(KEYINPUT101), .B(KEYINPUT23), .Z(n362) );
  XOR2_X1 U467 ( .A(KEYINPUT104), .B(n652), .Z(n363) );
  AND2_X1 U468 ( .A1(n649), .A2(n542), .ZN(n364) );
  XOR2_X1 U469 ( .A(n565), .B(n564), .Z(n365) );
  XNOR2_X1 U470 ( .A(n480), .B(n479), .ZN(n570) );
  NAND2_X1 U471 ( .A1(n689), .A2(n688), .ZN(n366) );
  XOR2_X1 U472 ( .A(n697), .B(n696), .Z(n367) );
  XOR2_X1 U473 ( .A(n620), .B(KEYINPUT62), .Z(n368) );
  XNOR2_X1 U474 ( .A(n409), .B(n489), .ZN(n690) );
  XOR2_X1 U475 ( .A(KEYINPUT48), .B(KEYINPUT96), .Z(n369) );
  XOR2_X1 U476 ( .A(n690), .B(n691), .Z(n370) );
  NOR2_X1 U477 ( .A1(G952), .A2(n688), .ZN(n705) );
  XNOR2_X1 U478 ( .A(KEYINPUT95), .B(KEYINPUT56), .ZN(n371) );
  NAND2_X1 U479 ( .A1(n701), .A2(G210), .ZN(n389) );
  XNOR2_X1 U480 ( .A(n400), .B(n399), .ZN(G60) );
  XNOR2_X2 U481 ( .A(n522), .B(n521), .ZN(n729) );
  NOR2_X1 U482 ( .A1(n607), .A2(n606), .ZN(n376) );
  XNOR2_X1 U483 ( .A(n405), .B(n369), .ZN(n404) );
  XNOR2_X2 U484 ( .A(n462), .B(n463), .ZN(n649) );
  NAND2_X1 U485 ( .A1(n376), .A2(n608), .ZN(n405) );
  NOR2_X1 U486 ( .A1(n390), .A2(n714), .ZN(n615) );
  NOR2_X1 U487 ( .A1(n703), .A2(G902), .ZN(n480) );
  XNOR2_X1 U488 ( .A(n468), .B(n377), .ZN(n472) );
  XNOR2_X1 U489 ( .A(n465), .B(n362), .ZN(n377) );
  XNOR2_X1 U490 ( .A(n379), .B(n378), .ZN(n573) );
  NOR2_X1 U491 ( .A1(n572), .A2(n649), .ZN(n379) );
  XNOR2_X2 U492 ( .A(n450), .B(n433), .ZN(n434) );
  XNOR2_X2 U493 ( .A(n381), .B(n380), .ZN(n450) );
  XNOR2_X2 U494 ( .A(G119), .B(KEYINPUT69), .ZN(n380) );
  NOR2_X2 U495 ( .A1(n730), .A2(n628), .ZN(n536) );
  NOR2_X2 U496 ( .A1(n384), .A2(n383), .ZN(n628) );
  XNOR2_X1 U497 ( .A(n387), .B(n371), .ZN(G51) );
  XNOR2_X1 U498 ( .A(n390), .B(n724), .ZN(n723) );
  NAND2_X1 U499 ( .A1(n679), .A2(n390), .ZN(n680) );
  NAND2_X2 U500 ( .A1(n617), .A2(n643), .ZN(n390) );
  NAND2_X1 U501 ( .A1(n582), .A2(n413), .ZN(n391) );
  XNOR2_X1 U502 ( .A(n562), .B(n393), .ZN(n392) );
  INV_X1 U503 ( .A(KEYINPUT77), .ZN(n393) );
  INV_X1 U504 ( .A(n570), .ZN(n651) );
  NAND2_X1 U505 ( .A1(n541), .A2(n647), .ZN(n561) );
  INV_X1 U506 ( .A(n714), .ZN(n397) );
  NAND2_X1 U507 ( .A1(n398), .A2(n687), .ZN(n494) );
  AND2_X1 U508 ( .A1(n398), .A2(n364), .ZN(n624) );
  XNOR2_X1 U509 ( .A(n539), .B(KEYINPUT100), .ZN(n398) );
  NAND2_X1 U510 ( .A1(n701), .A2(G475), .ZN(n402) );
  NAND2_X1 U511 ( .A1(n668), .A2(n665), .ZN(n576) );
  XNOR2_X1 U512 ( .A(n406), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U513 ( .A1(n690), .A2(n618), .ZN(n438) );
  XNOR2_X1 U514 ( .A(n429), .B(n436), .ZN(n410) );
  XNOR2_X2 U515 ( .A(n434), .B(n435), .ZN(n706) );
  NOR2_X1 U516 ( .A1(n412), .A2(KEYINPUT91), .ZN(n683) );
  OR2_X2 U517 ( .A1(n615), .A2(KEYINPUT2), .ZN(n412) );
  XNOR2_X1 U518 ( .A(n415), .B(n414), .ZN(G75) );
  NAND2_X1 U519 ( .A1(n417), .A2(n416), .ZN(n415) );
  XNOR2_X1 U520 ( .A(n685), .B(n418), .ZN(n417) );
  INV_X1 U521 ( .A(KEYINPUT92), .ZN(n418) );
  XNOR2_X2 U522 ( .A(n419), .B(n359), .ZN(n574) );
  XNOR2_X1 U523 ( .A(n489), .B(n420), .ZN(n694) );
  XNOR2_X1 U524 ( .A(n490), .B(n488), .ZN(n420) );
  XNOR2_X1 U525 ( .A(n535), .B(n534), .ZN(n554) );
  INV_X1 U526 ( .A(n464), .ZN(n427) );
  INV_X1 U527 ( .A(KEYINPUT114), .ZN(n563) );
  NAND2_X1 U528 ( .A1(n665), .A2(n363), .ZN(n525) );
  NOR2_X1 U529 ( .A1(n581), .A2(n663), .ZN(n441) );
  XNOR2_X1 U530 ( .A(KEYINPUT117), .B(KEYINPUT42), .ZN(n578) );
  XNOR2_X2 U531 ( .A(n497), .B(KEYINPUT4), .ZN(n722) );
  INV_X1 U532 ( .A(n722), .ZN(n423) );
  INV_X1 U533 ( .A(G101), .ZN(n422) );
  NAND2_X1 U534 ( .A1(n423), .A2(n422), .ZN(n425) );
  NAND2_X1 U535 ( .A1(G101), .A2(n722), .ZN(n424) );
  NAND2_X1 U536 ( .A1(n425), .A2(n424), .ZN(n459) );
  XOR2_X1 U537 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n431) );
  XNOR2_X1 U538 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n430) );
  XNOR2_X1 U539 ( .A(n431), .B(n430), .ZN(n436) );
  XNOR2_X1 U540 ( .A(n510), .B(n500), .ZN(n435) );
  OR2_X1 U541 ( .A1(G237), .A2(G902), .ZN(n439) );
  NAND2_X1 U542 ( .A1(G210), .A2(n439), .ZN(n437) );
  XNOR2_X2 U543 ( .A(n438), .B(n437), .ZN(n581) );
  NAND2_X1 U544 ( .A1(n439), .A2(G214), .ZN(n440) );
  XNOR2_X1 U545 ( .A(n440), .B(KEYINPUT97), .ZN(n663) );
  XNOR2_X1 U546 ( .A(n441), .B(KEYINPUT19), .ZN(n597) );
  XNOR2_X1 U547 ( .A(n443), .B(n442), .ZN(n445) );
  NAND2_X1 U548 ( .A1(n445), .A2(G952), .ZN(n444) );
  XNOR2_X1 U549 ( .A(n444), .B(KEYINPUT98), .ZN(n678) );
  NOR2_X1 U550 ( .A1(G953), .A2(n678), .ZN(n560) );
  NAND2_X1 U551 ( .A1(G902), .A2(n445), .ZN(n557) );
  XNOR2_X1 U552 ( .A(G898), .B(KEYINPUT99), .ZN(n712) );
  NAND2_X1 U553 ( .A1(G953), .A2(n712), .ZN(n708) );
  NOR2_X1 U554 ( .A1(n557), .A2(n708), .ZN(n446) );
  NOR2_X1 U555 ( .A1(n560), .A2(n446), .ZN(n447) );
  NOR2_X2 U556 ( .A1(n597), .A2(n447), .ZN(n448) );
  XNOR2_X2 U557 ( .A(n448), .B(KEYINPUT0), .ZN(n539) );
  XNOR2_X1 U558 ( .A(G472), .B(KEYINPUT106), .ZN(n463) );
  INV_X1 U559 ( .A(n485), .ZN(n449) );
  XNOR2_X1 U560 ( .A(n450), .B(n449), .ZN(n458) );
  NAND2_X1 U561 ( .A1(n512), .A2(G210), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n452), .B(n451), .ZN(n456) );
  XNOR2_X1 U563 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U564 ( .A(n456), .B(n455), .Z(n457) );
  XNOR2_X1 U565 ( .A(n458), .B(n457), .ZN(n461) );
  INV_X1 U566 ( .A(n459), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n620) );
  NOR2_X1 U568 ( .A1(n620), .A2(G902), .ZN(n462) );
  XOR2_X1 U569 ( .A(n649), .B(KEYINPUT6), .Z(n586) );
  XNOR2_X1 U570 ( .A(KEYINPUT10), .B(n464), .ZN(n511) );
  XOR2_X1 U571 ( .A(n487), .B(n511), .Z(n720) );
  XOR2_X1 U572 ( .A(KEYINPUT24), .B(KEYINPUT79), .Z(n465) );
  XOR2_X1 U573 ( .A(KEYINPUT89), .B(G110), .Z(n467) );
  XNOR2_X1 U574 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U575 ( .A(KEYINPUT90), .B(KEYINPUT8), .Z(n470) );
  NAND2_X1 U576 ( .A1(G234), .A2(n688), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n470), .B(n469), .ZN(n495) );
  NAND2_X1 U578 ( .A1(n495), .A2(G221), .ZN(n471) );
  XNOR2_X1 U579 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U580 ( .A(n720), .B(n473), .ZN(n703) );
  NAND2_X1 U581 ( .A1(G234), .A2(n618), .ZN(n474) );
  XNOR2_X1 U582 ( .A(KEYINPUT20), .B(n474), .ZN(n481) );
  NAND2_X1 U583 ( .A1(G217), .A2(n481), .ZN(n478) );
  XOR2_X1 U584 ( .A(KEYINPUT102), .B(KEYINPUT25), .Z(n476) );
  XNOR2_X1 U585 ( .A(KEYINPUT103), .B(KEYINPUT78), .ZN(n475) );
  XNOR2_X1 U586 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U587 ( .A1(n481), .A2(G221), .ZN(n482) );
  XNOR2_X1 U588 ( .A(n482), .B(KEYINPUT21), .ZN(n652) );
  XOR2_X1 U589 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n484) );
  XNOR2_X1 U590 ( .A(n484), .B(n483), .ZN(n486) );
  XNOR2_X1 U591 ( .A(n486), .B(n485), .ZN(n490) );
  XNOR2_X1 U592 ( .A(n487), .B(n421), .ZN(n488) );
  XOR2_X1 U593 ( .A(n574), .B(KEYINPUT1), .Z(n523) );
  NAND2_X1 U594 ( .A1(n647), .A2(n523), .ZN(n538) );
  OR2_X1 U595 ( .A1(n586), .A2(n538), .ZN(n491) );
  XOR2_X1 U596 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n492) );
  XNOR2_X1 U597 ( .A(n494), .B(n493), .ZN(n520) );
  NAND2_X1 U598 ( .A1(G217), .A2(n495), .ZN(n496) );
  XNOR2_X1 U599 ( .A(n497), .B(G134), .ZN(n498) );
  XNOR2_X1 U600 ( .A(n498), .B(G122), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n500), .B(KEYINPUT7), .ZN(n501) );
  XNOR2_X1 U602 ( .A(n502), .B(n501), .ZN(n699) );
  XNOR2_X1 U603 ( .A(G478), .B(n503), .ZN(n543) );
  INV_X1 U604 ( .A(n543), .ZN(n524) );
  XNOR2_X1 U605 ( .A(KEYINPUT13), .B(G475), .ZN(n518) );
  XOR2_X1 U606 ( .A(KEYINPUT109), .B(G140), .Z(n505) );
  XNOR2_X1 U607 ( .A(n505), .B(n504), .ZN(n509) );
  XOR2_X1 U608 ( .A(KEYINPUT108), .B(KEYINPUT11), .Z(n507) );
  XNOR2_X1 U609 ( .A(KEYINPUT12), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U610 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U611 ( .A(n509), .B(n508), .ZN(n516) );
  XOR2_X1 U612 ( .A(n511), .B(n510), .Z(n514) );
  NAND2_X1 U613 ( .A1(G214), .A2(n512), .ZN(n513) );
  XNOR2_X1 U614 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n516), .B(n515), .ZN(n697) );
  NOR2_X1 U616 ( .A1(G902), .A2(n697), .ZN(n517) );
  XNOR2_X1 U617 ( .A(n518), .B(n517), .ZN(n544) );
  NAND2_X1 U618 ( .A1(n524), .A2(n544), .ZN(n584) );
  INV_X1 U619 ( .A(n584), .ZN(n519) );
  NAND2_X1 U620 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U621 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n521) );
  NOR2_X1 U622 ( .A1(n729), .A2(KEYINPUT65), .ZN(n533) );
  BUF_X1 U623 ( .A(n523), .Z(n646) );
  INV_X1 U624 ( .A(n539), .ZN(n526) );
  NOR2_X1 U625 ( .A1(n524), .A2(n544), .ZN(n665) );
  INV_X1 U626 ( .A(KEYINPUT22), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n528), .B(n527), .ZN(n532) );
  NAND2_X1 U628 ( .A1(n646), .A2(n586), .ZN(n529) );
  NOR2_X1 U629 ( .A1(n570), .A2(n529), .ZN(n530) );
  XNOR2_X1 U630 ( .A(n530), .B(KEYINPUT85), .ZN(n531) );
  NAND2_X1 U631 ( .A1(n533), .A2(n536), .ZN(n535) );
  NAND2_X1 U632 ( .A1(n537), .A2(n536), .ZN(n552) );
  NOR2_X1 U633 ( .A1(n649), .A2(n538), .ZN(n657) );
  NAND2_X1 U634 ( .A1(n539), .A2(n657), .ZN(n540) );
  XNOR2_X1 U635 ( .A(n540), .B(KEYINPUT31), .ZN(n639) );
  INV_X1 U636 ( .A(n574), .ZN(n541) );
  INV_X1 U637 ( .A(n561), .ZN(n542) );
  NOR2_X1 U638 ( .A1(n639), .A2(n624), .ZN(n545) );
  NOR2_X1 U639 ( .A1(n544), .A2(n543), .ZN(n638) );
  NAND2_X1 U640 ( .A1(n544), .A2(n543), .ZN(n585) );
  INV_X1 U641 ( .A(n585), .ZN(n635) );
  NOR2_X1 U642 ( .A1(n638), .A2(n635), .ZN(n596) );
  XNOR2_X1 U643 ( .A(KEYINPUT88), .B(n596), .ZN(n601) );
  NOR2_X1 U644 ( .A1(n545), .A2(n601), .ZN(n546) );
  XNOR2_X1 U645 ( .A(KEYINPUT112), .B(n546), .ZN(n550) );
  AND2_X1 U646 ( .A1(n570), .A2(n586), .ZN(n547) );
  NAND2_X1 U647 ( .A1(n548), .A2(n547), .ZN(n621) );
  INV_X1 U648 ( .A(n621), .ZN(n549) );
  NOR2_X1 U649 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U650 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X2 U651 ( .A(n556), .B(n555), .ZN(n714) );
  OR2_X1 U652 ( .A1(n688), .A2(n557), .ZN(n558) );
  NOR2_X1 U653 ( .A1(G900), .A2(n558), .ZN(n559) );
  NOR2_X1 U654 ( .A1(n560), .A2(n559), .ZN(n567) );
  NOR2_X1 U655 ( .A1(n561), .A2(n567), .ZN(n562) );
  NOR2_X1 U656 ( .A1(n649), .A2(n663), .ZN(n565) );
  AND2_X1 U657 ( .A1(n614), .A2(n635), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n566), .B(KEYINPUT40), .ZN(n732) );
  NOR2_X1 U659 ( .A1(n567), .A2(n652), .ZN(n568) );
  XNOR2_X1 U660 ( .A(n568), .B(KEYINPUT67), .ZN(n569) );
  NOR2_X1 U661 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U662 ( .A(KEYINPUT66), .B(n571), .ZN(n587) );
  INV_X1 U663 ( .A(n587), .ZN(n572) );
  NOR2_X1 U664 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U665 ( .A(n575), .B(KEYINPUT115), .ZN(n598) );
  INV_X1 U666 ( .A(n598), .ZN(n577) );
  NAND2_X1 U667 ( .A1(n577), .A2(n659), .ZN(n579) );
  NAND2_X1 U668 ( .A1(KEYINPUT47), .A2(n596), .ZN(n580) );
  NAND2_X1 U669 ( .A1(n580), .A2(KEYINPUT87), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n613), .A2(n582), .ZN(n583) );
  NOR2_X1 U671 ( .A1(n584), .A2(n583), .ZN(n631) );
  INV_X1 U672 ( .A(n646), .ZN(n593) );
  INV_X1 U673 ( .A(n613), .ZN(n590) );
  NOR2_X1 U674 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U675 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U676 ( .A(KEYINPUT36), .B(n591), .Z(n592) );
  NOR2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n641) );
  NAND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n607) );
  INV_X1 U679 ( .A(n596), .ZN(n667) );
  OR2_X1 U680 ( .A1(KEYINPUT87), .A2(n667), .ZN(n599) );
  NOR2_X1 U681 ( .A1(n598), .A2(n597), .ZN(n633) );
  NAND2_X1 U682 ( .A1(n599), .A2(n633), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n600), .A2(KEYINPUT47), .ZN(n605) );
  NOR2_X1 U684 ( .A1(KEYINPUT47), .A2(n601), .ZN(n602) );
  XNOR2_X1 U685 ( .A(KEYINPUT74), .B(n602), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n603), .A2(n633), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U688 ( .A(n609), .B(KEYINPUT113), .Z(n610) );
  NOR2_X1 U689 ( .A1(n646), .A2(n610), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT43), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n644) );
  NAND2_X1 U692 ( .A1(n614), .A2(n638), .ZN(n643) );
  NAND2_X1 U693 ( .A1(KEYINPUT2), .A2(n643), .ZN(n616) );
  INV_X1 U694 ( .A(n618), .ZN(n619) );
  XNOR2_X1 U695 ( .A(G101), .B(n621), .ZN(G3) );
  NAND2_X1 U696 ( .A1(n624), .A2(n635), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT118), .ZN(n623) );
  XNOR2_X1 U698 ( .A(G104), .B(n623), .ZN(G6) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n626) );
  NAND2_X1 U700 ( .A1(n624), .A2(n638), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U702 ( .A(G107), .B(n627), .ZN(G9) );
  XOR2_X1 U703 ( .A(G110), .B(n628), .Z(G12) );
  XOR2_X1 U704 ( .A(G128), .B(KEYINPUT29), .Z(n630) );
  NAND2_X1 U705 ( .A1(n633), .A2(n638), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(n631), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(KEYINPUT119), .ZN(G45) );
  NAND2_X1 U709 ( .A1(n633), .A2(n635), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n634), .B(G146), .ZN(G48) );
  NAND2_X1 U711 ( .A1(n639), .A2(n635), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(KEYINPUT120), .ZN(n637) );
  XNOR2_X1 U713 ( .A(G113), .B(n637), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(G116), .ZN(G18) );
  XNOR2_X1 U716 ( .A(G125), .B(n641), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n642), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U718 ( .A(G134), .B(n643), .ZN(G36) );
  XNOR2_X1 U719 ( .A(G140), .B(n644), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(KEYINPUT121), .ZN(G42) );
  OR2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U722 ( .A(KEYINPUT50), .B(n648), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT49), .B(n653), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(KEYINPUT51), .B(n658), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U730 ( .A(KEYINPUT122), .B(n661), .Z(n674) );
  NAND2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U733 ( .A(KEYINPUT123), .B(n666), .Z(n670) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n687), .A2(n671), .ZN(n672) );
  XOR2_X1 U737 ( .A(n672), .B(KEYINPUT124), .Z(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U739 ( .A(KEYINPUT125), .B(n675), .Z(n676) );
  XNOR2_X1 U740 ( .A(n676), .B(KEYINPUT52), .ZN(n677) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n686) );
  NOR2_X1 U742 ( .A1(KEYINPUT2), .A2(n714), .ZN(n679) );
  NAND2_X1 U743 ( .A1(n680), .A2(KEYINPUT91), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U746 ( .A1(n659), .A2(n687), .ZN(n689) );
  INV_X1 U747 ( .A(n705), .ZN(n692) );
  XNOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n691) );
  XOR2_X1 U749 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n693) );
  NOR2_X1 U750 ( .A1(n705), .A2(n695), .ZN(G54) );
  XOR2_X1 U751 ( .A(KEYINPUT59), .B(KEYINPUT64), .Z(n696) );
  NAND2_X1 U752 ( .A1(G478), .A2(n701), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n705), .A2(n700), .ZN(G63) );
  NAND2_X1 U755 ( .A1(G217), .A2(n701), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n705), .A2(n704), .ZN(G66) );
  XNOR2_X1 U758 ( .A(G101), .B(G110), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n718) );
  XOR2_X1 U761 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n711) );
  NAND2_X1 U762 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n711), .B(n710), .ZN(n713) );
  NOR2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U765 ( .A1(G953), .A2(n714), .ZN(n715) );
  NOR2_X1 U766 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U768 ( .A(n719), .B(n720), .Z(n721) );
  XNOR2_X1 U769 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U770 ( .A1(n723), .A2(n688), .ZN(n728) );
  XNOR2_X1 U771 ( .A(G227), .B(n724), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G953), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n728), .A2(n727), .ZN(G72) );
  XOR2_X1 U775 ( .A(n729), .B(G122), .Z(G24) );
  XOR2_X1 U776 ( .A(G119), .B(n730), .Z(G21) );
  XOR2_X1 U777 ( .A(n731), .B(G137), .Z(G39) );
  XNOR2_X1 U778 ( .A(G131), .B(KEYINPUT127), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(n732), .ZN(G33) );
endmodule

