//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n194), .A3(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G128), .B1(new_n200), .B2(KEYINPUT68), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n202), .B1(new_n205), .B2(new_n194), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n197), .B1(new_n201), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n194), .A2(new_n196), .A3(G128), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n208), .A2(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(G107), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n211), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT10), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT0), .A4(G128), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n226));
  XNOR2_X1  g040(.A(G143), .B(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT0), .A4(G128), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT0), .B(G128), .Z(new_n230));
  AOI22_X1  g044(.A1(new_n226), .A2(new_n229), .B1(new_n197), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n212), .B1(new_n213), .B2(G104), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n213), .A2(G104), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n211), .B1(new_n237), .B2(new_n214), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n239));
  AOI21_X1  g053(.A(KEYINPUT82), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND4_X1   g054(.A1(KEYINPUT82), .A2(new_n232), .A3(G101), .A4(new_n239), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n231), .B(new_n234), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  INV_X1    g057(.A(new_n196), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n197), .A2(new_n243), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n209), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n221), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n222), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n224), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT11), .B1(new_n251), .B2(G137), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(G137), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT65), .B(G131), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n252), .A2(new_n255), .B1(new_n251), .B2(G137), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n250), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT84), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n250), .A2(new_n265), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT83), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n259), .B(KEYINPUT83), .C1(new_n260), .C2(new_n261), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n224), .A2(new_n242), .A3(new_n249), .A4(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n192), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n221), .B1(new_n209), .B2(new_n245), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n208), .A2(new_n205), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n200), .A2(KEYINPUT68), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n205), .A2(new_n202), .A3(new_n194), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G128), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n278), .B2(new_n197), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n274), .B1(new_n279), .B2(new_n221), .ZN(new_n280));
  INV_X1    g094(.A(new_n262), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT12), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n248), .B1(new_n210), .B2(new_n247), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n262), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n285), .A3(new_n272), .ZN(new_n286));
  INV_X1    g100(.A(new_n192), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n187), .B(new_n188), .C1(new_n273), .C2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n187), .A2(new_n188), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n267), .A2(new_n192), .A3(new_n272), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n192), .B(KEYINPUT80), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(G469), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n289), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G214), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G110), .B(G122), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT8), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G116), .ZN(new_n305));
  INV_X1    g119(.A(G116), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT2), .B(G113), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G113), .B1(new_n305), .B2(KEYINPUT5), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT5), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(new_n308), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n247), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT69), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT69), .B1(new_n305), .B2(new_n307), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n319), .A2(new_n320), .A3(new_n314), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n321), .B2(new_n312), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n308), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G116), .B(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT69), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT5), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT85), .A3(new_n313), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n311), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n221), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n317), .B1(new_n330), .B2(KEYINPUT88), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n313), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n310), .B1(new_n332), .B2(new_n318), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n247), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n303), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n210), .A2(G125), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n231), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT7), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT87), .B(G224), .Z(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n190), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n338), .A2(new_n340), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n322), .A2(new_n311), .A3(new_n247), .A4(new_n328), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n309), .B1(new_n319), .B2(new_n320), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n311), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(new_n234), .C1(new_n240), .C2(new_n241), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n349), .A3(new_n301), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n279), .A2(new_n339), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n231), .A2(new_n339), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT7), .A4(new_n343), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n188), .B1(new_n337), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n344), .B1(new_n338), .B2(new_n340), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n352), .A3(new_n343), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n346), .A2(new_n349), .A3(new_n301), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n346), .A2(new_n349), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n301), .B(KEYINPUT86), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n362), .B1(new_n346), .B2(new_n349), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT6), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n359), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n300), .B1(new_n355), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n316), .B1(new_n334), .B2(new_n335), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n330), .A2(KEYINPUT88), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n302), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n354), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n368), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n350), .B1(new_n367), .B2(KEYINPUT6), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n358), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n299), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n298), .B1(new_n370), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT9), .B(G234), .ZN(new_n381));
  OAI21_X1  g195(.A(G221), .B1(new_n381), .B2(G902), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n296), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT93), .ZN(new_n384));
  NOR2_X1   g198(.A1(G475), .A2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n339), .A2(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G146), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n339), .B2(G140), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n387), .A2(KEYINPUT76), .A3(G125), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(G146), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT89), .A2(G143), .ZN(new_n398));
  NOR2_X1   g212(.A1(G237), .A2(G953), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(G214), .ZN(new_n400));
  INV_X1    g214(.A(G237), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n190), .A3(G214), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(KEYINPUT89), .A2(G143), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT89), .A2(G143), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n400), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n397), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n195), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n411), .A2(G214), .A3(new_n399), .A4(new_n398), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n404), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n414), .A2(KEYINPUT90), .A3(KEYINPUT18), .A4(G131), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n396), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n339), .A2(G140), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT76), .B1(new_n387), .B2(G125), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n392), .A2(new_n339), .A3(G140), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT16), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n425), .A2(KEYINPUT77), .A3(G146), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT77), .B1(new_n425), .B2(G146), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(KEYINPUT65), .A2(G131), .ZN(new_n429));
  NOR2_X1   g243(.A1(KEYINPUT65), .A2(G131), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n412), .A2(new_n431), .A3(new_n413), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n412), .B2(new_n413), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT91), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n258), .B1(new_n435), .B2(new_n400), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT91), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n412), .A2(new_n413), .A3(new_n431), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n388), .A2(new_n389), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n193), .B(new_n441), .C1(new_n423), .C2(new_n440), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n417), .B1(new_n428), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G113), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(new_n215), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n432), .A2(new_n433), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n420), .B(new_n193), .C1(new_n423), .C2(new_n424), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n425), .A2(G146), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n438), .A2(new_n450), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n446), .B(KEYINPUT92), .Z(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n417), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n386), .B1(new_n448), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n384), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n385), .B(KEYINPUT94), .Z(new_n462));
  INV_X1    g276(.A(KEYINPUT77), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n419), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n193), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n425), .A2(KEYINPUT77), .A3(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n436), .A2(new_n438), .ZN(new_n468));
  INV_X1    g282(.A(new_n441), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n395), .B2(KEYINPUT19), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n468), .A2(KEYINPUT91), .B1(new_n470), .B2(new_n193), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n471), .A3(new_n439), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n446), .B1(new_n472), .B2(new_n417), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n456), .A2(new_n417), .A3(new_n457), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n460), .B(new_n462), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT95), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n454), .B1(new_n449), .B2(new_n450), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n453), .A2(new_n452), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n416), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n444), .A2(new_n447), .B1(new_n480), .B2(new_n457), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n481), .C2(new_n386), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n434), .A2(new_n439), .A3(new_n442), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n416), .B1(new_n483), .B2(new_n467), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n458), .B1(new_n484), .B2(new_n446), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n485), .A2(KEYINPUT95), .A3(new_n460), .A4(new_n462), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n461), .A2(new_n477), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n446), .B1(new_n456), .B2(new_n417), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n188), .B1(new_n474), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT96), .B(G475), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G952), .ZN(new_n493));
  AOI211_X1 g307(.A(G953), .B(new_n493), .C1(G234), .C2(G237), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT21), .B(G898), .Z(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n188), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT99), .ZN(new_n499));
  INV_X1    g313(.A(G217), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n381), .A2(new_n500), .A3(G953), .ZN(new_n501));
  XNOR2_X1  g315(.A(G116), .B(G122), .ZN(new_n502));
  INV_X1    g316(.A(G122), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G116), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT14), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n502), .A2(new_n505), .A3(G107), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n213), .B1(new_n504), .B2(KEYINPUT14), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n502), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n243), .A2(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n195), .A2(G128), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n251), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n251), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n506), .A2(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT13), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n195), .A2(KEYINPUT97), .A3(KEYINPUT13), .A4(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(new_n516), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n517), .A2(new_n509), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G134), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n502), .A2(G107), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT98), .A4(new_n251), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT98), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n511), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n502), .A2(G107), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n523), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n501), .B(new_n514), .C1(new_n522), .C2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n502), .B(new_n213), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n521), .A2(new_n524), .A3(new_n526), .A4(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n501), .B1(new_n532), .B2(new_n514), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n188), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n536), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n514), .B1(new_n522), .B2(new_n528), .ZN(new_n539));
  INV_X1    g353(.A(new_n501), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n529), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n542), .B2(new_n188), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n499), .B1(new_n537), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n534), .A2(new_n536), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n188), .A3(new_n538), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(KEYINPUT99), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n498), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n487), .A2(new_n492), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n383), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G234), .ZN(new_n552));
  OAI21_X1  g366(.A(G217), .B1(new_n552), .B2(G902), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n553), .B(KEYINPUT74), .Z(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n391), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n243), .A2(G119), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n304), .A2(G128), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT23), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n243), .A2(G119), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT23), .ZN(new_n562));
  AOI211_X1 g376(.A(G110), .B(new_n557), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT24), .B(G110), .Z(new_n564));
  INV_X1    g378(.A(KEYINPUT75), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n561), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n558), .A2(KEYINPUT75), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n556), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n426), .B2(new_n427), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n572));
  INV_X1    g386(.A(G110), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n557), .B1(new_n560), .B2(new_n562), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n453), .B2(new_n452), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT78), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n569), .B1(new_n465), .B2(new_n466), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n576), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n585), .A3(new_n188), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT25), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n582), .A2(new_n585), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n555), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n582), .A2(new_n585), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n552), .B2(G217), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OR3_X1    g408(.A1(new_n590), .A2(KEYINPUT79), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT79), .B1(new_n590), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT30), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT66), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n257), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n254), .A2(G134), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n251), .A2(KEYINPUT66), .A3(G137), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n259), .B1(new_n603), .B2(new_n260), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n207), .B2(new_n209), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n231), .A2(new_n262), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n231), .A2(new_n262), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n608), .B(KEYINPUT30), .C1(new_n279), .C2(new_n604), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n348), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT26), .B(G101), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n399), .A2(G210), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g429(.A(new_n348), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n608), .B(new_n616), .C1(new_n279), .C2(new_n604), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n610), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  OR2_X1    g432(.A1(KEYINPUT71), .A2(KEYINPUT31), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n605), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n621), .A2(KEYINPUT28), .A3(new_n616), .A4(new_n608), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT28), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n348), .B1(new_n605), .B2(new_n606), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n615), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT71), .B(KEYINPUT31), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n610), .A2(new_n615), .A3(new_n617), .A4(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n620), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(G472), .A2(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT32), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n631), .A2(KEYINPUT32), .A3(new_n632), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G472), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT72), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n625), .A2(new_n639), .A3(new_n617), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n621), .A2(KEYINPUT72), .A3(new_n616), .A4(new_n608), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(KEYINPUT28), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n624), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT73), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT73), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n644), .A2(KEYINPUT29), .A3(new_n615), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n610), .A2(new_n617), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT29), .B1(new_n648), .B2(new_n627), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n626), .A2(new_n627), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n638), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n597), .B1(new_n637), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n551), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  INV_X1    g470(.A(new_n633), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n638), .B1(new_n631), .B2(new_n188), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n597), .A2(new_n659), .A3(new_n382), .A4(new_n296), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n298), .B(new_n498), .C1(new_n370), .C2(new_n379), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n487), .A2(new_n492), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT33), .B1(new_n501), .B2(KEYINPUT100), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n542), .B(new_n665), .Z(new_n666));
  NOR2_X1   g480(.A1(new_n535), .A2(G902), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n666), .A2(new_n667), .B1(new_n535), .B2(new_n534), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n663), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  AOI211_X1 g484(.A(KEYINPUT101), .B(new_n668), .C1(new_n487), .C2(new_n492), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  AND3_X1   g489(.A1(new_n544), .A2(new_n492), .A3(new_n547), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT20), .B1(new_n448), .B2(new_n458), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n385), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n461), .A2(new_n482), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n662), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT35), .B(G107), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NAND2_X1  g497(.A1(new_n571), .A2(new_n577), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n583), .A2(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n590), .B1(new_n592), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n551), .A2(new_n659), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  AND3_X1   g505(.A1(new_n631), .A2(KEYINPUT32), .A3(new_n632), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT32), .B1(new_n631), .B2(new_n632), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n646), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n645), .B1(new_n642), .B2(new_n624), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n615), .A2(KEYINPUT29), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n649), .A2(new_n650), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n188), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n687), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n355), .A2(new_n369), .A3(new_n300), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n299), .B1(new_n375), .B2(new_n378), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n297), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(G900), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n497), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n494), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n676), .A2(new_n679), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n703), .B1(new_n706), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n382), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n250), .A2(new_n265), .A3(new_n262), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n265), .B1(new_n250), .B2(new_n262), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n272), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n287), .ZN(new_n717));
  INV_X1    g531(.A(new_n288), .ZN(new_n718));
  AOI21_X1  g532(.A(G902), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n290), .B1(new_n719), .B2(new_n187), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n713), .B1(new_n720), .B2(new_n295), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n676), .A2(new_n679), .A3(new_n710), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(KEYINPUT102), .A3(new_n380), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n702), .A2(new_n712), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  NOR2_X1   g539(.A1(new_n704), .A2(new_n705), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT38), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n544), .A2(new_n547), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n664), .A2(new_n728), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n727), .A2(new_n298), .A3(new_n688), .A4(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n710), .B(KEYINPUT39), .Z(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(KEYINPUT40), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(KEYINPUT40), .ZN(new_n735));
  AOI21_X1  g549(.A(G902), .B1(new_n648), .B2(new_n615), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n640), .A2(new_n641), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(new_n615), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G472), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n694), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n730), .A2(new_n734), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G143), .ZN(G45));
  INV_X1    g556(.A(new_n710), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n743), .B(new_n668), .C1(new_n487), .C2(new_n492), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n702), .A2(new_n380), .A3(new_n721), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G146), .ZN(G48));
  AOI21_X1  g560(.A(new_n288), .B1(new_n716), .B2(new_n287), .ZN(new_n747));
  OAI21_X1  g561(.A(G469), .B1(new_n747), .B2(G902), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n289), .A3(new_n382), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n653), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n498), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n297), .B(new_n751), .C1(new_n704), .C2(new_n705), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n670), .A2(new_n671), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n492), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n485), .A2(new_n385), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT93), .B1(new_n757), .B2(KEYINPUT20), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n384), .B(new_n460), .C1(new_n485), .C2(new_n385), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT95), .B1(new_n677), .B2(new_n462), .ZN(new_n761));
  INV_X1    g575(.A(new_n462), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n481), .A2(new_n476), .A3(KEYINPUT20), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n756), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT101), .B1(new_n765), .B2(new_n668), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n664), .A2(new_n663), .A3(new_n669), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n661), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n748), .A2(new_n289), .A3(new_n382), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n769), .B(new_n597), .C1(new_n637), .C2(new_n652), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT103), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n755), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT41), .B(G113), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT104), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n772), .B(new_n774), .ZN(G15));
  NAND2_X1  g589(.A1(new_n661), .A2(new_n680), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n306), .ZN(G18));
  NAND3_X1  g592(.A1(new_n769), .A2(new_n380), .A3(new_n549), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n688), .B1(new_n637), .B2(new_n652), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n304), .ZN(G21));
  NOR3_X1   g596(.A1(new_n729), .A2(new_n752), .A3(new_n749), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n627), .B1(new_n695), .B2(new_n696), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n620), .A2(new_n630), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n658), .B1(new_n787), .B2(new_n632), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n588), .A2(new_n589), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n554), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n593), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n784), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n632), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n785), .B2(new_n786), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n795), .A2(KEYINPUT105), .A3(new_n658), .A4(new_n791), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n783), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT106), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT106), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n783), .B(new_n799), .C1(new_n793), .C2(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G122), .ZN(G24));
  NOR2_X1   g616(.A1(new_n749), .A2(new_n706), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n795), .A2(new_n687), .A3(new_n658), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n744), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G125), .ZN(G27));
  NAND3_X1  g620(.A1(new_n370), .A2(new_n297), .A3(new_n379), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n294), .A2(KEYINPUT107), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n294), .A2(KEYINPUT107), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n292), .A3(G469), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n289), .A2(new_n811), .A3(new_n291), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n812), .A3(new_n382), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n653), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n664), .A2(new_n669), .A3(new_n710), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT42), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n713), .B1(new_n720), .B2(new_n811), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n744), .A3(new_n808), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n637), .A2(new_n652), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT108), .B1(new_n820), .B2(new_n791), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n694), .A2(new_n701), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n792), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n819), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT42), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n817), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(new_n260), .ZN(G33));
  NAND2_X1  g642(.A1(new_n814), .A2(new_n722), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G134), .ZN(G36));
  NAND2_X1  g644(.A1(new_n292), .A2(new_n294), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT45), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n187), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n809), .A2(KEYINPUT45), .A3(new_n292), .A4(new_n810), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n290), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(KEYINPUT46), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n835), .A2(KEYINPUT46), .B1(new_n187), .B2(new_n719), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n713), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(new_n732), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n659), .A2(new_n687), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n765), .A2(new_n669), .ZN(new_n841));
  NOR2_X1   g655(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n840), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT44), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n807), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n839), .B(new_n848), .C1(new_n847), .C2(new_n846), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G137), .ZN(G39));
  XOR2_X1   g664(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n838), .A2(new_n852), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n822), .A2(new_n815), .A3(new_n597), .A4(new_n807), .ZN(new_n854));
  NOR2_X1   g668(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n853), .B(new_n854), .C1(new_n838), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(G140), .ZN(G42));
  NOR2_X1   g671(.A1(new_n843), .A2(new_n845), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n709), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n749), .A2(new_n807), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n821), .A2(new_n824), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(KEYINPUT119), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n865));
  INV_X1    g679(.A(new_n863), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(KEYINPUT48), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT48), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n865), .B(new_n869), .C1(new_n861), .C2(new_n866), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  INV_X1    g685(.A(new_n740), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n597), .A2(new_n872), .A3(new_n494), .A4(new_n860), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n493), .B(G953), .C1(new_n873), .C2(new_n672), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n793), .A2(new_n796), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n859), .A2(new_n803), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n871), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n874), .A2(new_n871), .A3(new_n876), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n868), .B(new_n870), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n727), .A2(new_n298), .A3(new_n769), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n859), .A2(new_n875), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n880), .B(new_n881), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n882), .B(KEYINPUT116), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n880), .A2(new_n881), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n887), .A2(new_n875), .A3(new_n859), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n853), .B1(new_n838), .B2(new_n855), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n748), .A2(new_n289), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n713), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n875), .A3(new_n808), .A4(new_n859), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n664), .A2(new_n669), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n862), .A2(new_n804), .B1(new_n873), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT51), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n890), .A2(new_n895), .A3(new_n900), .A4(new_n897), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n879), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n712), .A2(new_n723), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n296), .A2(new_n382), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n780), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n383), .A2(new_n815), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n903), .A2(new_n905), .B1(new_n702), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n729), .A2(new_n706), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n688), .A2(new_n743), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(new_n740), .A3(new_n818), .A4(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n907), .A2(KEYINPUT115), .A3(new_n805), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT52), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n724), .A2(new_n745), .A3(new_n910), .A4(new_n805), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n770), .A2(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n755), .B2(new_n771), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n918), .A2(new_n801), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n537), .A2(new_n543), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n664), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n660), .A2(new_n661), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n689), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT112), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n661), .A2(new_n924), .A3(new_n664), .A4(new_n669), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n664), .A2(new_n669), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT112), .B1(new_n926), .B2(new_n752), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n660), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n655), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT113), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n928), .A2(new_n655), .A3(KEYINPUT113), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n679), .A2(new_n492), .A3(new_n920), .A4(new_n710), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n807), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n702), .A2(new_n721), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT114), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT114), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n702), .A2(new_n721), .A3(new_n938), .A4(new_n935), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n804), .A2(new_n818), .A3(new_n744), .A4(new_n808), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n937), .A2(new_n829), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n827), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n916), .A2(new_n919), .A3(new_n933), .A4(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT53), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n912), .B1(new_n911), .B2(new_n915), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n913), .A2(KEYINPUT52), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n916), .A2(new_n947), .ZN(new_n948));
  AND4_X1   g762(.A1(new_n829), .A2(new_n937), .A3(new_n939), .A4(new_n940), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n813), .A2(new_n815), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n823), .B1(new_n822), .B2(new_n792), .ZN(new_n951));
  AOI211_X1 g765(.A(KEYINPUT108), .B(new_n791), .C1(new_n694), .C2(new_n701), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n953), .A2(KEYINPUT42), .B1(new_n814), .B2(new_n816), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n949), .A2(new_n954), .A3(new_n918), .A4(new_n801), .ZN(new_n955));
  INV_X1    g769(.A(new_n932), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT113), .B1(new_n928), .B2(new_n655), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n689), .B(new_n922), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT53), .B1(new_n948), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT54), .B1(new_n946), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n948), .A2(new_n959), .A3(KEYINPUT53), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT54), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n902), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(G952), .B2(G953), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n892), .B(KEYINPUT49), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n841), .A2(new_n791), .A3(new_n298), .A4(new_n713), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n968), .A2(new_n969), .A3(new_n872), .A4(new_n727), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT111), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(G75));
  NOR2_X1   g786(.A1(new_n376), .A2(new_n377), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(new_n358), .ZN(new_n974));
  XOR2_X1   g788(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n975));
  XOR2_X1   g789(.A(new_n974), .B(new_n975), .Z(new_n976));
  INV_X1    g790(.A(G210), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n977), .B(new_n188), .C1(new_n962), .C2(new_n963), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT121), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n979), .A2(KEYINPUT56), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n976), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n188), .B1(new_n962), .B2(new_n963), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(G210), .ZN(new_n984));
  INV_X1    g798(.A(new_n976), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(new_n980), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n190), .A2(G952), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n982), .A2(new_n986), .A3(new_n988), .ZN(G51));
  XNOR2_X1  g803(.A(new_n290), .B(KEYINPUT57), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n964), .B1(new_n962), .B2(new_n963), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n747), .B(KEYINPUT122), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n983), .A2(new_n834), .A3(new_n833), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n987), .B1(new_n995), .B2(new_n996), .ZN(G54));
  AND2_X1   g811(.A1(KEYINPUT58), .A2(G475), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n983), .A2(new_n485), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n485), .B1(new_n983), .B2(new_n998), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n999), .A2(new_n1000), .A3(new_n987), .ZN(G60));
  NAND2_X1  g815(.A1(G478), .A2(G902), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT59), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n666), .B(new_n1003), .C1(new_n991), .C2(new_n992), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n988), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n961), .A2(new_n965), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n666), .B1(new_n1006), .B2(new_n1003), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1005), .A2(new_n1007), .ZN(G63));
  NAND2_X1  g822(.A1(new_n962), .A2(new_n963), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G217), .A2(G902), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT60), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1009), .A2(new_n686), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1011), .B1(new_n962), .B2(new_n963), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1013), .B(new_n988), .C1(new_n591), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(KEYINPUT61), .B1(new_n1013), .B2(KEYINPUT123), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1018));
  INV_X1    g832(.A(new_n591), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n987), .B1(new_n1014), .B2(new_n686), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT123), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n1014), .B2(new_n686), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1020), .B(new_n1021), .C1(new_n1023), .C2(KEYINPUT61), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1017), .A2(new_n1024), .ZN(G66));
  AOI21_X1  g839(.A(new_n190), .B1(new_n342), .B2(new_n495), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n919), .A2(new_n933), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(new_n1027), .B2(new_n190), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n973), .B1(G898), .B2(new_n190), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1029), .B(KEYINPUT124), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1028), .B(new_n1030), .ZN(G69));
  NAND2_X1  g845(.A1(new_n607), .A2(new_n609), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(new_n470), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n921), .B1(new_n664), .B2(new_n669), .ZN(new_n1034));
  OR4_X1    g848(.A1(new_n653), .A2(new_n1034), .A3(new_n733), .A4(new_n807), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n849), .A2(new_n856), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n741), .A2(new_n805), .A3(new_n907), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT62), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n741), .A2(KEYINPUT62), .A3(new_n805), .A4(new_n907), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1033), .B1(new_n1041), .B2(G953), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n190), .A2(G900), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1043), .B(KEYINPUT126), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n849), .A2(new_n856), .ZN(new_n1045));
  AND4_X1   g859(.A1(new_n732), .A2(new_n838), .A3(new_n863), .A4(new_n908), .ZN(new_n1046));
  XNOR2_X1  g860(.A(new_n1046), .B(KEYINPUT127), .ZN(new_n1047));
  AND4_X1   g861(.A1(new_n805), .A2(new_n954), .A3(new_n829), .A4(new_n907), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1044), .B1(new_n1049), .B2(new_n190), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1042), .B1(new_n1050), .B2(new_n1033), .ZN(new_n1051));
  OAI21_X1  g865(.A(KEYINPUT125), .B1(new_n1050), .B2(new_n1033), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1053));
  INV_X1    g867(.A(new_n1053), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  OAI221_X1 g869(.A(new_n1042), .B1(KEYINPUT125), .B2(new_n1053), .C1(new_n1050), .C2(new_n1033), .ZN(new_n1056));
  AND2_X1   g870(.A1(new_n1055), .A2(new_n1056), .ZN(G72));
  NAND2_X1  g871(.A1(G472), .A2(G902), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT63), .Z(new_n1059));
  NAND2_X1  g873(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1060), .A2(new_n1035), .A3(new_n1045), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1059), .B1(new_n1061), .B2(new_n1027), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n1062), .A2(new_n615), .A3(new_n648), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1059), .B1(new_n1049), .B2(new_n1027), .ZN(new_n1064));
  NAND4_X1  g878(.A1(new_n1064), .A2(new_n627), .A3(new_n617), .A4(new_n610), .ZN(new_n1065));
  NAND3_X1  g879(.A1(new_n1063), .A2(new_n1065), .A3(new_n988), .ZN(new_n1066));
  OR2_X1    g880(.A1(new_n946), .A2(new_n960), .ZN(new_n1067));
  INV_X1    g881(.A(new_n1059), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n648), .A2(new_n627), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1068), .B1(new_n1069), .B2(new_n618), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1066), .B1(new_n1067), .B2(new_n1070), .ZN(G57));
endmodule


