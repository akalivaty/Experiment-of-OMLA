//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT0), .B(G128), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT64), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n187), .A2(KEYINPUT0), .A3(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n203), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G134), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n205), .A2(new_n210), .A3(new_n213), .A4(new_n207), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n189), .A2(new_n198), .A3(KEYINPUT65), .A4(new_n199), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n202), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n202), .A2(new_n215), .A3(new_n219), .A4(new_n216), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n192), .B(G146), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n190), .A3(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(new_n227), .A3(new_n224), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n187), .A2(new_n229), .A3(G128), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n204), .B2(new_n209), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n214), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n221), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n235), .A2(KEYINPUT68), .A3(new_n214), .A4(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n218), .A2(new_n220), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT69), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT70), .B1(new_n242), .B2(G116), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT2), .B(G113), .Z(new_n250));
  XOR2_X1   g064(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n238), .A2(new_n252), .A3(new_n239), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n231), .A2(new_n233), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n200), .B(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n254), .B1(new_n256), .B2(new_n215), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT30), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n241), .A2(new_n251), .A3(new_n253), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n257), .A2(KEYINPUT72), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n266));
  INV_X1    g080(.A(G237), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n266), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n259), .A2(new_n265), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n265), .A4(new_n273), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(KEYINPUT31), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n261), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n263), .A2(new_n264), .B1(new_n251), .B2(new_n238), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n286), .B2(KEYINPUT28), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(new_n273), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n288), .B1(new_n278), .B2(new_n280), .ZN(new_n294));
  INV_X1    g108(.A(new_n291), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n283), .B(new_n273), .C1(new_n285), .C2(new_n282), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n273), .B1(new_n259), .B2(new_n265), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n265), .B1(new_n260), .B2(new_n257), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n284), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n272), .A2(new_n299), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n300), .A2(new_n297), .A3(new_n301), .ZN(new_n308));
  OAI21_X1  g122(.A(G472), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n292), .A2(new_n296), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n190), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT78), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  OR3_X1    g129(.A1(new_n315), .A2(KEYINPUT16), .A3(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(new_n190), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G119), .B(G128), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT76), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT24), .B(G110), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(G119), .B2(new_n222), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n242), .A2(KEYINPUT23), .A3(G128), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n326), .A2(new_n327), .B1(G119), .B2(new_n222), .ZN(new_n328));
  OAI22_X1  g142(.A1(new_n324), .A2(KEYINPUT77), .B1(G110), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n319), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n318), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n317), .A2(new_n190), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(G110), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n334), .B(new_n335), .C1(new_n321), .C2(new_n323), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G137), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(KEYINPUT79), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G902), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n331), .A2(new_n336), .A3(new_n340), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(KEYINPUT80), .B2(KEYINPUT25), .ZN(new_n347));
  INV_X1    g161(.A(G217), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(G234), .B2(new_n344), .ZN(new_n349));
  NOR2_X1   g163(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n349), .A2(G902), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n343), .A2(new_n354), .A3(new_n345), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n343), .B2(new_n345), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(KEYINPUT82), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n352), .B2(new_n357), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n267), .A2(new_n268), .A3(G214), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(G143), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(G131), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(new_n318), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n311), .B(KEYINPUT92), .ZN(new_n368));
  MUX2_X1   g182(.A(new_n311), .B(new_n368), .S(KEYINPUT19), .Z(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n369), .B2(G146), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT18), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n365), .B1(new_n371), .B2(new_n213), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n365), .A2(new_n213), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n368), .A2(G146), .ZN(new_n374));
  OAI221_X1 g188(.A(new_n372), .B1(new_n373), .B2(new_n371), .C1(new_n374), .C2(new_n313), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT93), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n370), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n370), .B2(new_n375), .ZN(new_n379));
  XNOR2_X1  g193(.A(G113), .B(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT94), .B(G104), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n378), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT17), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n366), .A2(new_n385), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n373), .A2(new_n385), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n333), .A4(new_n332), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n388), .A2(new_n375), .A3(new_n383), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G475), .A2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT20), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(new_n391), .C1(new_n384), .C2(new_n389), .ZN(new_n395));
  INV_X1    g209(.A(G475), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n383), .B1(new_n388), .B2(new_n375), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n344), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT95), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n393), .A2(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT13), .B1(new_n222), .B2(G143), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n203), .ZN(new_n404));
  XNOR2_X1  g218(.A(G128), .B(G143), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G122), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G116), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n245), .A2(G122), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G107), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT97), .B1(new_n409), .B2(KEYINPUT14), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(KEYINPUT14), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n409), .A2(KEYINPUT97), .A3(KEYINPUT14), .ZN(new_n419));
  OAI21_X1  g233(.A(G107), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n405), .A2(G134), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n405), .A2(G134), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n411), .B2(new_n410), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT9), .B(G234), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n427), .A2(new_n348), .A3(G953), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n425), .A2(KEYINPUT98), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n429), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n415), .A2(new_n424), .A3(new_n428), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT98), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n434), .A3(new_n344), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(KEYINPUT99), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT99), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n431), .A2(new_n434), .A3(new_n440), .A4(new_n344), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n438), .B1(new_n442), .B2(new_n437), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n268), .A2(G952), .ZN(new_n444));
  NAND2_X1  g258(.A1(G234), .A2(G237), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT21), .B(G898), .Z(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(G902), .A3(G953), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n402), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G104), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G107), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT3), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n411), .A2(G104), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n451), .A2(G107), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(G101), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n453), .A2(new_n456), .B1(new_n451), .B2(G107), .ZN(new_n462));
  INV_X1    g276(.A(G101), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(KEYINPUT4), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n459), .A2(new_n460), .A3(new_n466), .A4(G101), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n251), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n458), .A2(new_n454), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n463), .B1(new_n452), .B2(KEYINPUT85), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n462), .A2(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n247), .A2(KEYINPUT5), .A3(new_n248), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(G113), .C1(KEYINPUT5), .C2(new_n248), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n250), .A2(new_n247), .A3(new_n248), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(G110), .B(G122), .Z(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(KEYINPUT90), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n472), .B1(new_n475), .B2(new_n474), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI22_X1  g296(.A1(new_n476), .A2(KEYINPUT90), .B1(KEYINPUT8), .B2(new_n477), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n477), .A2(KEYINPUT8), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n200), .A2(G125), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(G125), .B2(new_n235), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT89), .B(G224), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n268), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n268), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT7), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n491), .A2(KEYINPUT7), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n468), .A2(new_n476), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n477), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT6), .A3(new_n479), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n489), .B(new_n492), .Z(new_n500));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n501), .A3(new_n477), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n495), .A2(new_n496), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n496), .B1(new_n495), .B2(new_n503), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n506));
  OR3_X1    g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  OAI21_X1  g322(.A(G214), .B1(G237), .B2(G902), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G221), .B1(new_n427), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(G469), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n225), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n225), .A2(new_n513), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n230), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n472), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n235), .B2(new_n472), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n215), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT12), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n521), .A3(new_n215), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n256), .A2(new_n467), .A3(new_n465), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n472), .A2(KEYINPUT10), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n526));
  AOI22_X1  g340(.A1(new_n235), .A2(new_n525), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n524), .A2(new_n527), .A3(new_n214), .A4(new_n212), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n527), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n215), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n528), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n268), .A2(G227), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT83), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G140), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  MUX2_X1   g351(.A(new_n529), .B(new_n533), .S(new_n537), .Z(new_n538));
  AOI21_X1  g352(.A(new_n512), .B1(new_n538), .B2(new_n344), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT88), .B(G469), .Z(new_n540));
  AND4_X1   g354(.A1(new_n528), .A2(new_n520), .A3(new_n522), .A4(new_n537), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n531), .B2(new_n528), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n344), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n511), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n450), .A2(new_n510), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n310), .A2(new_n363), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT100), .B(G101), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(G3));
  NAND2_X1  g363(.A1(new_n290), .A2(new_n291), .ZN(new_n550));
  OAI21_X1  g364(.A(G472), .B1(new_n294), .B2(G902), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n509), .B1(new_n504), .B2(new_n505), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT101), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT101), .B(new_n509), .C1(new_n504), .C2(new_n505), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(G478), .B1(new_n439), .B2(new_n441), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n428), .B(KEYINPUT102), .Z(new_n561));
  AOI21_X1  g375(.A(KEYINPUT103), .B1(new_n425), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n433), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n425), .A2(KEYINPUT103), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT33), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n568));
  INV_X1    g382(.A(new_n434), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n568), .B1(new_n569), .B2(new_n430), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(G478), .A3(new_n344), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n402), .B1(new_n560), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n558), .A2(new_n573), .A3(new_n449), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n362), .A2(new_n545), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n553), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT34), .B(G104), .Z(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(G6));
  NAND2_X1  g394(.A1(new_n393), .A2(new_n395), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n401), .A2(new_n400), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n443), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n558), .A2(new_n449), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n553), .A2(new_n575), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G107), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT106), .B(KEYINPUT35), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G9));
  NOR2_X1   g403(.A1(new_n450), .A2(new_n510), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n337), .A2(KEYINPUT107), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n337), .A2(KEYINPUT107), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n353), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n352), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n545), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n590), .A2(new_n600), .A3(new_n550), .A4(new_n551), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT37), .B(G110), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G12));
  INV_X1    g417(.A(new_n545), .ZN(new_n604));
  AND4_X1   g418(.A1(new_n310), .A2(new_n604), .A3(new_n558), .A4(new_n598), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n446), .B1(G900), .B2(new_n448), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n584), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G128), .ZN(G30));
  XOR2_X1   g424(.A(new_n606), .B(KEYINPUT39), .Z(new_n611));
  NOR2_X1   g425(.A1(new_n545), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n613), .A2(KEYINPUT40), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(KEYINPUT40), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n402), .A2(new_n443), .ZN(new_n616));
  AND4_X1   g430(.A1(new_n509), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n344), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n276), .A2(new_n277), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n303), .B2(new_n272), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT108), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n296), .A3(new_n292), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n507), .A2(new_n508), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT38), .Z(new_n627));
  NAND4_X1  g441(.A1(new_n617), .A2(new_n599), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G143), .ZN(G45));
  NAND4_X1  g443(.A1(new_n310), .A2(new_n604), .A3(new_n558), .A4(new_n598), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n573), .A2(new_n606), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n190), .ZN(G48));
  INV_X1    g447(.A(new_n541), .ZN(new_n634));
  INV_X1    g448(.A(new_n542), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n543), .B(new_n511), .C1(new_n636), .C2(new_n512), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n310), .A2(new_n574), .A3(new_n363), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT41), .B(G113), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G15));
  NAND4_X1  g455(.A1(new_n310), .A2(new_n585), .A3(new_n363), .A4(new_n638), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G116), .ZN(G18));
  NAND3_X1  g457(.A1(new_n556), .A2(new_n638), .A3(new_n557), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n556), .A2(new_n638), .A3(KEYINPUT109), .A4(new_n557), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n450), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n310), .A3(new_n598), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G119), .ZN(G21));
  OR2_X1    g464(.A1(new_n304), .A2(new_n273), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n295), .B1(new_n281), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n290), .A2(new_n344), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT110), .B(G472), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n449), .ZN(new_n656));
  NOR4_X1   g470(.A1(new_n644), .A2(new_n656), .A3(new_n402), .A4(new_n443), .ZN(new_n657));
  INV_X1    g471(.A(new_n358), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G122), .ZN(G24));
  NAND2_X1  g474(.A1(new_n646), .A2(new_n647), .ZN(new_n661));
  INV_X1    g475(.A(new_n631), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n655), .A2(new_n661), .A3(new_n662), .A4(new_n598), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G125), .ZN(G27));
  AOI21_X1  g478(.A(KEYINPUT32), .B1(new_n290), .B2(new_n291), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n294), .A2(new_n293), .A3(new_n295), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT112), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT113), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT112), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n296), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n292), .B2(new_n296), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT112), .B1(new_n550), .B2(new_n293), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT113), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n671), .A2(new_n674), .A3(new_n309), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n538), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n676), .B1(new_n533), .B2(new_n537), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n677), .A2(new_n512), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n543), .B1(new_n512), .B2(new_n344), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n511), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n509), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n507), .B2(new_n508), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n631), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n675), .A2(new_n658), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n687));
  INV_X1    g501(.A(new_n310), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n362), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n681), .A2(new_n684), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n631), .A2(KEYINPUT42), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G131), .ZN(G33));
  NAND3_X1  g508(.A1(new_n689), .A2(new_n608), .A3(new_n690), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G134), .ZN(G36));
  AOI21_X1  g510(.A(new_n583), .B1(new_n560), .B2(new_n572), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT43), .Z(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n553), .A3(new_n599), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n684), .B1(new_n699), .B2(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(KEYINPUT44), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n512), .A2(new_n344), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n703));
  OR3_X1    g517(.A1(new_n677), .A2(new_n703), .A3(new_n678), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n512), .B1(new_n538), .B2(new_n703), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n543), .B1(new_n706), .B2(KEYINPUT46), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n511), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(new_n611), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n208), .ZN(G39));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n709), .B(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n631), .A2(new_n363), .A3(new_n684), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n688), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G140), .ZN(G42));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n698), .A2(new_n446), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n658), .A3(new_n655), .ZN(new_n720));
  NOR4_X1   g534(.A1(new_n720), .A2(new_n509), .A3(new_n627), .A4(new_n637), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT50), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n684), .A2(new_n446), .A3(new_n637), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n362), .ZN(new_n725));
  INV_X1    g539(.A(new_n625), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AOI211_X1 g542(.A(new_n436), .B(G902), .C1(new_n567), .C2(new_n570), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n583), .A2(new_n559), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n655), .A2(new_n598), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n698), .A2(new_n724), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n728), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n722), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n720), .A2(new_n684), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n543), .B1(new_n636), .B2(new_n512), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(new_n511), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT119), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n735), .B1(new_n714), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT120), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n718), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n737), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n714), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n718), .B1(new_n743), .B2(new_n735), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n722), .A2(new_n744), .A3(new_n733), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n583), .B1(new_n729), .B2(new_n559), .ZN(new_n746));
  INV_X1    g560(.A(new_n661), .ZN(new_n747));
  OAI221_X1 g561(.A(new_n444), .B1(new_n746), .B2(new_n727), .C1(new_n720), .C2(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT121), .Z(new_n749));
  AND3_X1   g563(.A1(new_n741), .A2(new_n745), .A3(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n639), .A2(new_n642), .A3(new_n649), .A4(new_n659), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n507), .A2(new_n449), .A3(new_n508), .A4(new_n509), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n442), .A2(new_n437), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n402), .B1(new_n753), .B2(new_n438), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n752), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n575), .A3(new_n550), .A4(new_n551), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n547), .A2(new_n601), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT114), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n547), .A2(new_n759), .A3(new_n601), .A4(new_n756), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n751), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n402), .A2(new_n683), .A3(new_n443), .A4(new_n606), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n310), .A2(new_n762), .A3(new_n604), .A4(new_n598), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n731), .A2(new_n662), .A3(new_n690), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n695), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n687), .A2(new_n761), .A3(new_n765), .A4(new_n692), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n663), .B1(new_n630), .B2(new_n607), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n632), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n606), .B(KEYINPUT115), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n511), .B(new_n769), .C1(new_n679), .C2(new_n680), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n558), .A2(new_n616), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n625), .A2(new_n772), .A3(new_n599), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n768), .A2(KEYINPUT52), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(new_n768), .B2(new_n773), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(KEYINPUT116), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n605), .A2(new_n662), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n609), .A2(new_n777), .A3(new_n663), .A4(new_n773), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n625), .A2(new_n772), .A3(new_n599), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n767), .A2(new_n632), .A3(new_n782), .A4(new_n779), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n766), .B1(new_n776), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT117), .B1(new_n785), .B2(KEYINPUT53), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n687), .A2(new_n692), .A3(new_n761), .A4(new_n765), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n783), .B1(new_n780), .B2(new_n781), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n778), .A2(KEYINPUT116), .A3(new_n779), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT118), .B1(new_n780), .B2(new_n774), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n766), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n780), .A2(KEYINPUT118), .A3(new_n774), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n786), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT54), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n775), .B2(new_n783), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n787), .A2(new_n796), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n792), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n785), .A2(KEYINPUT53), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n675), .A2(new_n658), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n732), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT48), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n750), .A2(new_n799), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(G952), .B2(G953), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n658), .A2(new_n511), .A3(new_n509), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(KEYINPUT49), .B2(new_n736), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n697), .C1(KEYINPUT49), .C2(new_n736), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(new_n627), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n811), .B1(new_n625), .B2(new_n815), .ZN(G75));
  AOI21_X1  g630(.A(new_n344), .B1(new_n803), .B2(new_n804), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(G210), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n499), .A2(new_n502), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(new_n500), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT55), .Z(new_n822));
  AND3_X1   g636(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n818), .B2(new_n819), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n268), .A2(G952), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(G51));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n795), .B2(new_n796), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n792), .B(new_n766), .C1(new_n776), .C2(new_n784), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT54), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n806), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n702), .B(KEYINPUT57), .Z(new_n832));
  OAI22_X1  g646(.A1(new_n831), .A2(new_n832), .B1(new_n542), .B2(new_n541), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n817), .A2(new_n704), .A3(new_n705), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n825), .B1(new_n833), .B2(new_n834), .ZN(G54));
  INV_X1    g649(.A(new_n825), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n817), .A2(KEYINPUT58), .A3(G475), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n836), .B1(new_n837), .B2(new_n390), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n390), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n839), .A2(KEYINPUT122), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(KEYINPUT122), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(G60));
  NAND2_X1  g656(.A1(G478), .A2(G902), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT59), .Z(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n567), .B2(new_n570), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n825), .B1(new_n830), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n799), .B2(new_n806), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n571), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT123), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n846), .B(new_n850), .C1(new_n847), .C2(new_n571), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(G63));
  NAND2_X1  g666(.A1(G217), .A2(G902), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT60), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n803), .B2(new_n804), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n825), .B1(new_n855), .B2(new_n596), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n355), .A2(new_n356), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n858), .B2(new_n855), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g674(.A(new_n268), .B1(new_n447), .B2(new_n490), .ZN(new_n861));
  INV_X1    g675(.A(new_n761), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n862), .B2(new_n268), .ZN(new_n863));
  INV_X1    g677(.A(G898), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n820), .B1(new_n864), .B2(G953), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n863), .B(new_n865), .ZN(G69));
  NAND3_X1  g680(.A1(new_n241), .A2(new_n253), .A3(new_n258), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT124), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(new_n369), .ZN(new_n869));
  INV_X1    g683(.A(new_n716), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n573), .A2(new_n584), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT125), .Z(new_n872));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n613), .A3(new_n684), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n711), .B(new_n870), .C1(new_n689), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n628), .A2(new_n768), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT62), .Z(new_n876));
  AND2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n869), .B1(new_n877), .B2(G953), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n268), .A2(G900), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT126), .Z(new_n880));
  NAND3_X1  g694(.A1(new_n807), .A2(new_n558), .A3(new_n616), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n881), .A2(new_n701), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(new_n710), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n716), .A2(new_n695), .A3(new_n768), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n693), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n880), .B1(new_n885), .B2(new_n268), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n878), .B1(new_n869), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n268), .B1(G227), .B2(G900), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(G72));
  XNOR2_X1  g703(.A(new_n619), .B(KEYINPUT63), .ZN(new_n890));
  INV_X1    g704(.A(new_n620), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n798), .B(new_n890), .C1(new_n891), .C2(new_n301), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT127), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n874), .A2(new_n761), .A3(new_n876), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n272), .B1(new_n894), .B2(new_n890), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n259), .A2(new_n265), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n883), .A2(new_n884), .A3(new_n693), .A4(new_n761), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n890), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n274), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n836), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n893), .A2(new_n900), .ZN(G57));
endmodule


