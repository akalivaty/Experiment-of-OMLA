//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT92), .Z(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT82), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT83), .B(G148gat), .Z(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT84), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(G148gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT82), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n212), .B(new_n213), .C1(new_n208), .C2(new_n207), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n210), .A2(new_n214), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n215), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT80), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n218), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n215), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n222), .A2(KEYINPUT81), .A3(new_n223), .A4(new_n225), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n208), .A2(G148gat), .ZN(new_n230));
  OAI22_X1  g029(.A1(new_n205), .A2(new_n230), .B1(new_n221), .B2(new_n216), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n220), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT86), .B(KEYINPUT3), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G211gat), .B(G218gat), .Z(new_n239));
  XOR2_X1   g038(.A(G197gat), .B(G204gat), .Z(new_n240));
  AOI21_X1  g039(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n241));
  OR3_X1    g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT75), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT75), .B1(new_n242), .B2(new_n243), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n243), .A2(KEYINPUT93), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT93), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n237), .B(new_n251), .C1(new_n244), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n235), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n210), .A2(new_n214), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n219), .A2(new_n215), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n232), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n203), .B1(new_n250), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g060(.A(new_n244), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(KEYINPUT29), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n202), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n248), .A2(KEYINPUT76), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n246), .B2(new_n247), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n265), .B1(new_n269), .B2(new_n238), .ZN(new_n270));
  OAI21_X1  g069(.A(G22gat), .B1(new_n260), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n236), .A2(new_n237), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n268), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n264), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G22gat), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n238), .A2(new_n249), .B1(new_n258), .B2(new_n254), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n274), .B(new_n275), .C1(new_n276), .C2(new_n203), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n271), .A2(KEYINPUT94), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n276), .B2(new_n203), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT94), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n280), .A3(G22gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(G78gat), .B(G106gat), .ZN(new_n282));
  INV_X1    g081(.A(G50gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT91), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT95), .B(G22gat), .C1(new_n260), .C2(new_n270), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(new_n286), .A3(new_n277), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT95), .B1(new_n279), .B2(G22gat), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n278), .A2(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n299), .A2(KEYINPUT65), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(KEYINPUT65), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n296), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G183gat), .B(G190gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n294), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(KEYINPUT66), .B(new_n294), .C1(new_n302), .C2(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(new_n306), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n297), .B(KEYINPUT67), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n300), .A2(new_n301), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n296), .A2(KEYINPUT25), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n311), .A2(new_n313), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(new_n310), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n319));
  INV_X1    g118(.A(G183gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT27), .B1(new_n320), .B2(KEYINPUT68), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT68), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  AND4_X1   g124(.A1(new_n319), .A2(new_n321), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n319), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  OR3_X1    g127(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT69), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n320), .A2(new_n325), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n314), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT26), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n312), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n330), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT69), .B1(new_n326), .B2(new_n328), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n329), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT71), .B(KEYINPUT1), .Z(new_n340));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n343), .A2(new_n342), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(KEYINPUT1), .ZN(new_n346));
  OAI22_X1  g145(.A1(new_n344), .A2(new_n345), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G227gat), .ZN(new_n350));
  INV_X1    g149(.A(G233gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n318), .A2(new_n338), .A3(new_n347), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n352), .A4(new_n353), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n293), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G15gat), .B(G43gat), .Z(new_n363));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n353), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n350), .B2(new_n351), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n368), .B(KEYINPUT34), .Z(new_n369));
  AOI21_X1  g168(.A(KEYINPUT33), .B1(new_n356), .B2(new_n357), .ZN(new_n370));
  INV_X1    g169(.A(new_n365), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n358), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n366), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n292), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n375));
  AND2_X1   g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n339), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n339), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n248), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n376), .B1(new_n339), .B2(new_n237), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n269), .B1(new_n382), .B2(new_n377), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT78), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT30), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n381), .B2(new_n383), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n375), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n381), .A2(new_n383), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n388), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n391), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(KEYINPUT79), .A3(new_n389), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT0), .ZN(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  XOR2_X1   g202(.A(KEYINPUT88), .B(KEYINPUT6), .Z(new_n404));
  AOI21_X1  g203(.A(new_n348), .B1(new_n234), .B2(new_n235), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n406), .B(KEYINPUT3), .C1(new_n220), .C2(new_n233), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n257), .A2(new_n411), .A3(new_n348), .A4(new_n232), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n234), .A2(KEYINPUT87), .A3(new_n411), .A4(new_n348), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n257), .A2(new_n348), .A3(new_n232), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT4), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n410), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n419), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n348), .B1(new_n257), .B2(new_n232), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n220), .A2(new_n233), .A3(new_n347), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(new_n220), .B2(new_n233), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT85), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n408), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n421), .B1(new_n430), .B2(new_n405), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT5), .B1(new_n417), .B2(new_n412), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n403), .B(new_n404), .C1(new_n427), .C2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n403), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n425), .B1(new_n431), .B2(new_n418), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n410), .A2(new_n419), .A3(new_n432), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n427), .A2(new_n403), .A3(new_n433), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n404), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT89), .A4(new_n404), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n399), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n358), .A2(new_n370), .A3(new_n371), .ZN(new_n445));
  AOI221_X4 g244(.A(new_n293), .B1(KEYINPUT33), .B2(new_n365), .C1(new_n356), .C2(new_n357), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT73), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n366), .A2(new_n448), .A3(new_n372), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n369), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT74), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT74), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n453), .B(new_n369), .C1(new_n447), .C2(new_n449), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n374), .B(new_n444), .C1(new_n452), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  INV_X1    g255(.A(new_n373), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n369), .B1(new_n366), .B2(new_n372), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n292), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n396), .A2(new_n397), .A3(new_n389), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n440), .B1(new_n404), .B2(new_n438), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n456), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n417), .A2(new_n412), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n419), .B1(new_n410), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n435), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n422), .A2(new_n423), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT39), .B1(new_n474), .B2(new_n421), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n477), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n463), .A3(new_n438), .A4(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n388), .B1(new_n393), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n481), .B2(new_n393), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT38), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n269), .A2(new_n382), .A3(new_n377), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n380), .A2(new_n248), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT37), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n394), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n292), .B(new_n480), .C1(new_n490), .C2(new_n465), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n444), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n461), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n457), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n445), .A2(KEYINPUT73), .A3(new_n446), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n448), .B1(new_n366), .B2(new_n372), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n451), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n453), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n450), .A2(KEYINPUT74), .A3(new_n451), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n459), .A2(KEYINPUT36), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n494), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n492), .B1(new_n505), .B2(KEYINPUT96), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n496), .B1(new_n452), .B2(new_n454), .ZN(new_n507));
  INV_X1    g306(.A(new_n504), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n507), .A2(new_n508), .B1(new_n461), .B2(new_n493), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n469), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT16), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n514), .A2(G1gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT101), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT101), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(G8gat), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT102), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT103), .B(G8gat), .Z(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G43gat), .B(G50gat), .Z(new_n528));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G43gat), .B(G50gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT97), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  OAI221_X1 g334(.A(new_n533), .B1(KEYINPUT15), .B2(new_n531), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  OR3_X1    g335(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT99), .Z(new_n540));
  OR2_X1    g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n538), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n537), .B2(KEYINPUT98), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(KEYINPUT98), .B2(new_n537), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n534), .B2(new_n535), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n545), .A2(KEYINPUT15), .A3(new_n530), .A4(new_n532), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n527), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n547), .A2(KEYINPUT100), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT100), .B1(new_n547), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n527), .B1(new_n550), .B2(new_n547), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n513), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI221_X1 g357(.A(new_n527), .B1(new_n550), .B2(new_n547), .C1(new_n551), .C2(new_n552), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(KEYINPUT18), .A3(new_n556), .A4(new_n549), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n527), .A2(new_n548), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n549), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n556), .B(KEYINPUT13), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G197gat), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT11), .B(G169gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT12), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n558), .A2(new_n572), .A3(new_n560), .A4(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n512), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G99gat), .B(G106gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT106), .ZN(new_n591));
  OAI221_X1 g390(.A(new_n591), .B1(new_n550), .B2(new_n547), .C1(new_n551), .C2(new_n552), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT107), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n547), .A2(new_n590), .B1(KEYINPUT41), .B2(new_n577), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n592), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n581), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n580), .A3(new_n597), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  INV_X1    g403(.A(G64gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(G57gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(G57gat), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(KEYINPUT104), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(KEYINPUT104), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  OR2_X1    g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT9), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n607), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT9), .B1(new_n615), .B2(new_n606), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n610), .A3(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n527), .B1(new_n604), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n604), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G127gat), .B(G155gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT105), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n624), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n621), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n603), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n590), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n618), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n590), .A2(new_n614), .A3(new_n617), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(KEYINPUT108), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT108), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n640), .A3(new_n618), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT10), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n635), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT109), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n639), .A2(G230gat), .A3(G233gat), .A4(new_n641), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n647), .A2(new_n648), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n645), .A2(KEYINPUT110), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n645), .A2(KEYINPUT110), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n656), .A2(new_n648), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n653), .B1(new_n657), .B2(new_n651), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n634), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n442), .A2(KEYINPUT111), .A3(new_n443), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT111), .B1(new_n442), .B2(new_n443), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n576), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g463(.A1(new_n576), .A2(new_n463), .A3(new_n659), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(KEYINPUT112), .A3(G8gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(G8gat), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT112), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n665), .A2(KEYINPUT42), .A3(new_n671), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n666), .B(new_n669), .C1(new_n674), .C2(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(G15gat), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n576), .A2(new_n677), .A3(new_n459), .A4(new_n659), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n576), .A2(new_n659), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n507), .A2(new_n508), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n678), .B1(new_n682), .B2(new_n677), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n461), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n658), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n632), .ZN(new_n688));
  INV_X1    g487(.A(new_n603), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n576), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n662), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n691), .A2(G29gat), .A3(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n456), .A2(new_n468), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n491), .B1(new_n509), .B2(new_n510), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n505), .A2(KEYINPUT96), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n689), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n509), .A2(new_n491), .B1(new_n456), .B2(new_n468), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n702), .B2(new_n689), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n575), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n692), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n693), .A2(KEYINPUT45), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n694), .A2(new_n706), .A3(new_n707), .ZN(G1328gat));
  INV_X1    g507(.A(new_n691), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n710));
  AOI211_X1 g509(.A(G36gat), .B(new_n464), .C1(new_n710), .C2(KEYINPUT46), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n710), .B2(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n705), .B2(new_n464), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n710), .A2(KEYINPUT46), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n709), .A2(new_n715), .A3(new_n711), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n460), .A2(G43gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT115), .B1(new_n705), .B2(new_n680), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n705), .A2(KEYINPUT115), .A3(new_n680), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n719), .ZN(new_n725));
  OAI21_X1  g524(.A(G43gat), .B1(new_n705), .B2(new_n680), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n724), .A2(new_n729), .ZN(G1330gat));
  NOR2_X1   g529(.A1(new_n705), .A2(new_n292), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n461), .A2(new_n283), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n731), .A2(new_n283), .B1(new_n691), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI221_X1 g534(.A(KEYINPUT48), .B1(new_n691), .B2(new_n732), .C1(new_n731), .C2(new_n283), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1331gat));
  NOR4_X1   g536(.A1(new_n702), .A2(new_n574), .A3(new_n634), .A4(new_n687), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n662), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n463), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  NAND2_X1  g543(.A1(new_n738), .A2(new_n681), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n460), .A2(G71gat), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n745), .A2(G71gat), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n738), .A2(new_n461), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n702), .A2(new_n689), .ZN(new_n751));
  INV_X1    g550(.A(new_n632), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n574), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(KEYINPUT51), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(new_n753), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n751), .A2(KEYINPUT117), .A3(KEYINPUT51), .A4(new_n753), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n761), .A2(new_n585), .A3(new_n658), .A4(new_n662), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n687), .A2(new_n574), .A3(new_n752), .ZN(new_n763));
  INV_X1    g562(.A(new_n700), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n703), .B(new_n763), .C1(new_n512), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n701), .A2(new_n767), .A3(new_n703), .A4(new_n763), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n766), .A2(new_n662), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n762), .B1(new_n769), .B2(new_n585), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n687), .A2(G92gat), .A3(new_n464), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n761), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  OAI21_X1  g572(.A(G92gat), .B1(new_n765), .B2(new_n464), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n766), .A2(new_n463), .A3(new_n768), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n754), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n776), .A2(G92gat), .B1(new_n777), .B2(new_n771), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(new_n773), .ZN(G1337gat));
  NAND3_X1  g578(.A1(new_n766), .A2(new_n681), .A3(new_n768), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n766), .A2(KEYINPUT118), .A3(new_n768), .A4(new_n681), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(G99gat), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n460), .A2(new_n687), .A3(G99gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n761), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1338gat));
  NOR3_X1   g586(.A1(new_n687), .A2(G106gat), .A3(new_n292), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT119), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n761), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n765), .B2(new_n292), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n766), .A2(new_n461), .A3(new_n768), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n795), .A2(G106gat), .B1(new_n777), .B2(new_n790), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(new_n792), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n654), .A2(new_n798), .A3(new_n655), .ZN(new_n799));
  INV_X1    g598(.A(new_n651), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n642), .A2(new_n635), .A3(new_n644), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT120), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n652), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n804), .A2(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n808), .A2(new_n810), .A3(new_n574), .A4(new_n653), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n556), .B1(new_n559), .B2(new_n549), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n562), .A2(new_n563), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n569), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n573), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n658), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n603), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n810), .A2(new_n653), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n603), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n809), .B2(new_n801), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n632), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n659), .A2(new_n575), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n662), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n463), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n292), .A2(new_n373), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n501), .B2(new_n502), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n574), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n462), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n574), .A2(G113gat), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(G1340gat));
  AOI21_X1  g634(.A(G120gat), .B1(new_n830), .B2(new_n658), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n658), .A2(G120gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n832), .B2(new_n632), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n632), .A2(G127gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n829), .B2(new_n840), .ZN(G1342gat));
  OR2_X1    g640(.A1(new_n689), .A2(G134gat), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n829), .A2(KEYINPUT56), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n832), .B2(new_n689), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT56), .B1(new_n829), .B2(new_n842), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NOR3_X1   g645(.A1(new_n681), .A2(new_n692), .A3(new_n463), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n461), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(new_n821), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n817), .B2(KEYINPUT121), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n851), .B(new_n603), .C1(new_n811), .C2(new_n816), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n632), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n848), .B1(new_n853), .B2(new_n823), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT57), .B1(new_n824), .B2(new_n461), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n574), .B(new_n847), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n680), .A2(new_n461), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n575), .A2(G141gat), .A3(new_n463), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n824), .A2(new_n662), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT58), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT58), .B1(new_n856), .B2(G141gat), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n825), .B2(new_n858), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n824), .A2(KEYINPUT122), .A3(new_n662), .A4(new_n859), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n860), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n863), .A2(new_n872), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n847), .A2(new_n658), .ZN(new_n874));
  INV_X1    g673(.A(new_n855), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n876), .B(new_n292), .C1(new_n822), .C2(new_n823), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT59), .B1(new_n879), .B2(new_n204), .ZN(new_n880));
  INV_X1    g679(.A(new_n207), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(KEYINPUT59), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n847), .B1(new_n854), .B2(new_n855), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n687), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n866), .A2(new_n867), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n464), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n658), .A2(new_n881), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(G1345gat));
  OAI21_X1  g688(.A(G155gat), .B1(new_n883), .B2(new_n632), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n752), .A2(new_n217), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n887), .B2(new_n891), .ZN(G1346gat));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n464), .A3(new_n603), .ZN(new_n893));
  INV_X1    g692(.A(new_n883), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n689), .A2(new_n218), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n893), .A2(new_n218), .B1(new_n894), .B2(new_n895), .ZN(G1347gat));
  AOI21_X1  g695(.A(new_n662), .B1(new_n822), .B2(new_n823), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n462), .A3(new_n463), .ZN(new_n898));
  INV_X1    g697(.A(G169gat), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n575), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n828), .A3(new_n463), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n574), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n900), .B1(new_n899), .B2(new_n903), .ZN(G1348gat));
  INV_X1    g703(.A(G176gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n898), .A2(new_n905), .A3(new_n687), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n901), .B2(new_n687), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(G1349gat));
  NAND2_X1  g710(.A1(new_n752), .A2(new_n327), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n901), .A2(KEYINPUT125), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(new_n901), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n898), .B2(new_n632), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n898), .B2(new_n689), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT61), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n902), .A2(new_n325), .A3(new_n603), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n875), .A2(new_n878), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n681), .A2(new_n464), .A3(new_n662), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n926), .A2(G197gat), .A3(new_n574), .A4(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(G197gat), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n858), .A2(new_n464), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n897), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n933), .B2(new_n575), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n928), .A2(new_n934), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n687), .A2(G204gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n933), .A2(KEYINPUT62), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n658), .B(new_n927), .C1(new_n855), .C2(new_n877), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G204gat), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT62), .B1(new_n933), .B2(new_n937), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n938), .A2(new_n940), .A3(new_n941), .A4(KEYINPUT127), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1353gat));
  OR3_X1    g745(.A1(new_n933), .A2(G211gat), .A3(new_n632), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n926), .A2(new_n752), .A3(new_n927), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  NAND3_X1  g750(.A1(new_n926), .A2(new_n603), .A3(new_n927), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G218gat), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n689), .A2(G218gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n933), .B2(new_n954), .ZN(G1355gat));
endmodule


