//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1322, new_n1323, new_n1324, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n210), .A2(G20), .A3(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n205), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n208), .B(new_n213), .C1(new_n220), .C2(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XOR2_X1   g0022(.A(G250), .B(G257), .Z(new_n223));
  XNOR2_X1  g0023(.A(G264), .B(G270), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT65), .B(KEYINPUT66), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n227), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  NOR2_X1   g0040(.A1(G20), .A2(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G150), .ZN(new_n242));
  INV_X1    g0042(.A(G20), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT8), .B(G58), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(G33), .ZN(new_n245));
  OAI221_X1 g0045(.A(new_n242), .B1(new_n201), .B2(new_n243), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n211), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n253), .A2(new_n250), .A3(G13), .A4(G20), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n248), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n243), .A2(G1), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n257), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(KEYINPUT68), .A3(G50), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n255), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n252), .A2(new_n254), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n258), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n249), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT73), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n273), .B(new_n274), .C1(new_n202), .C2(new_n271), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n211), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n280), .A2(new_n250), .A3(G274), .A4(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n278), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT72), .B(G200), .Z(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n288), .B1(new_n275), .B2(new_n277), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n270), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n295), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n297), .A2(KEYINPUT74), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n269), .B(new_n296), .C1(new_n298), .C2(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n269), .A2(new_n296), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT10), .B1(new_n297), .B2(KEYINPUT74), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n266), .C1(G169), .C2(new_n293), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n299), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT17), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n244), .A2(new_n257), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n264), .A2(new_n244), .B1(new_n255), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT77), .ZN(new_n310));
  INV_X1    g0110(.A(G68), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT3), .ZN(new_n312));
  INV_X1    g0112(.A(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n243), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT7), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n314), .A2(KEYINPUT7), .A3(new_n243), .A4(new_n315), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n311), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G58), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n311), .ZN(new_n322));
  NOR2_X1   g0122(.A1(G58), .A2(G68), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n241), .A2(G159), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n310), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT7), .B1(new_n330), .B2(new_n243), .ZN(new_n331));
  INV_X1    g0131(.A(new_n319), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n325), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(KEYINPUT77), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n324), .A2(new_n325), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n320), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n248), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n309), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(G223), .A2(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n285), .A2(G1698), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n343), .C1(new_n328), .C2(new_n329), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G87), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n277), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n280), .A2(G232), .A3(new_n286), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n284), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT78), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT78), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n280), .B1(new_n344), .B2(new_n345), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n284), .A2(new_n348), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n352), .A2(new_n353), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n355), .A2(new_n356), .B1(new_n294), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n307), .B1(new_n341), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n355), .A2(new_n361), .B1(new_n303), .B2(new_n357), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n341), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n309), .ZN(new_n364));
  INV_X1    g0164(.A(new_n248), .ZN(new_n365));
  INV_X1    g0165(.A(new_n338), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n333), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n337), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n327), .A2(new_n335), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT78), .B1(new_n347), .B2(new_n349), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n352), .A2(new_n353), .A3(new_n351), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n361), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n357), .A2(new_n303), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT18), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n356), .B1(new_n371), .B2(new_n372), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n357), .A2(new_n294), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(KEYINPUT17), .A3(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n359), .A2(new_n363), .A3(new_n376), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n229), .A2(new_n272), .ZN(new_n382));
  INV_X1    g0182(.A(G238), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n271), .ZN(new_n386));
  INV_X1    g0186(.A(G107), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n330), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(new_n277), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n280), .A2(G244), .A3(new_n286), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n284), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n294), .ZN(new_n392));
  INV_X1    g0192(.A(new_n291), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n391), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT15), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(G87), .ZN(new_n396));
  INV_X1    g0196(.A(G87), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT69), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n245), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n395), .A2(G87), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT69), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g0205(.A(KEYINPUT8), .B(G58), .Z(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n241), .B1(G20), .B2(G77), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n248), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT70), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n257), .A2(new_n202), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n263), .A2(new_n365), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n252), .A2(new_n202), .A3(new_n254), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n365), .B1(new_n405), .B2(new_n407), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n413), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT70), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n415), .A2(KEYINPUT71), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT71), .B1(new_n415), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n394), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(new_n418), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n277), .B1(new_n271), .B2(G107), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n382), .A2(new_n384), .B1(new_n314), .B2(new_n315), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n284), .A2(new_n390), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n361), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n389), .A2(new_n303), .A3(new_n284), .A4(new_n390), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n306), .A2(new_n381), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n241), .A2(G50), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n434), .B1(new_n243), .B2(G68), .C1(new_n202), .C2(new_n245), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n248), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT11), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n255), .A2(G68), .A3(new_n260), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n263), .A2(G68), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G97), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G226), .A2(G1698), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n229), .B2(G1698), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(new_n271), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT75), .B1(new_n448), .B2(new_n280), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n285), .A2(new_n272), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n229), .A2(G1698), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n328), .C2(new_n329), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n280), .B1(new_n452), .B2(new_n444), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT75), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n284), .B1(new_n383), .B2(new_n287), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n443), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI211_X1 g0259(.A(KEYINPUT13), .B(new_n457), .C1(new_n449), .C2(new_n455), .ZN(new_n460));
  OAI21_X1  g0260(.A(G200), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n453), .A2(new_n454), .ZN(new_n462));
  AOI211_X1 g0262(.A(KEYINPUT75), .B(new_n280), .C1(new_n452), .C2(new_n444), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT13), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(new_n443), .A3(new_n458), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(G190), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n442), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT76), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n361), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT14), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(G169), .B1(new_n459), .B2(new_n460), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT76), .A3(KEYINPUT14), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n472), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n465), .A2(G179), .A3(new_n466), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n473), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n442), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n433), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G264), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT82), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n271), .A2(new_n484), .A3(G264), .A4(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n330), .A2(G303), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n271), .A2(G257), .A3(new_n272), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n277), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n250), .A2(G45), .ZN(new_n490));
  OR2_X1    g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(G274), .A4(new_n280), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n282), .A2(G1), .ZN(new_n496));
  INV_X1    g0296(.A(new_n492), .ZN(new_n497));
  NOR2_X1   g0297(.A1(KEYINPUT5), .A2(G41), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(G274), .B1(new_n276), .B2(new_n211), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT79), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n493), .A2(new_n277), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n495), .A2(new_n501), .B1(new_n502), .B2(G270), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n489), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n264), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n250), .A2(G33), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n255), .A2(G116), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  INV_X1    g0309(.A(G97), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n509), .B(new_n243), .C1(G33), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(G20), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n248), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT20), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n506), .B(new_n508), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n504), .A2(KEYINPUT21), .A3(G169), .A4(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n517), .A2(G179), .A3(new_n489), .A4(new_n503), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n361), .B1(new_n489), .B2(new_n503), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT21), .B1(new_n521), .B2(new_n517), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n517), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n489), .A2(new_n503), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n356), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n356), .B1(new_n489), .B2(new_n503), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT83), .B1(new_n528), .B2(new_n517), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(G190), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n243), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n387), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n400), .A2(G116), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n243), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n537), .A2(KEYINPUT22), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(KEYINPUT22), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(KEYINPUT24), .B(new_n536), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n248), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n263), .A2(G107), .A3(new_n365), .A4(new_n507), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT25), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n252), .A2(new_n546), .A3(new_n387), .A4(new_n254), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n252), .A2(new_n387), .A3(new_n254), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT25), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT84), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n545), .A2(new_n549), .A3(new_n552), .A4(new_n547), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n544), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(new_n272), .C1(new_n328), .C2(new_n329), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G294), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n277), .A2(new_n559), .B1(new_n502), .B2(G264), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n495), .A2(new_n501), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G169), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(G179), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n555), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n560), .A2(new_n294), .A3(new_n561), .ZN(new_n567));
  AOI21_X1  g0367(.A(G200), .B1(new_n560), .B2(new_n561), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n544), .B(new_n554), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n272), .C1(new_n328), .C2(new_n329), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n277), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT80), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n282), .B2(G1), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n250), .A2(KEYINPUT80), .A3(G45), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n280), .A2(new_n577), .A3(G250), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n280), .A2(G274), .A3(new_n496), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(G169), .B1(new_n575), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n277), .B2(new_n574), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n303), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n404), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n403), .B1(new_n401), .B2(new_n402), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n255), .A3(new_n507), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n243), .B1(new_n444), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G97), .A2(G107), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n397), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n243), .B(G68), .C1(new_n328), .C2(new_n329), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n590), .B1(new_n245), .B2(new_n510), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n248), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n254), .B(new_n252), .C1(new_n586), .C2(new_n587), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n589), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n255), .A2(G87), .A3(new_n507), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT81), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT81), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n255), .A2(new_n604), .A3(G87), .A4(new_n507), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n601), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n575), .A2(new_n582), .A3(new_n294), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n584), .B2(new_n393), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n585), .A2(new_n600), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G244), .B(new_n272), .C1(new_n328), .C2(new_n329), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT4), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n509), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n277), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n495), .A2(new_n501), .B1(new_n502), .B2(G257), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n361), .ZN(new_n619));
  OAI21_X1  g0419(.A(G107), .B1(new_n331), .B2(new_n332), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT6), .ZN(new_n621));
  AND2_X1   g0421(.A1(G97), .A2(G107), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n592), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n387), .A2(KEYINPUT6), .A3(G97), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n625), .A2(G20), .B1(G77), .B2(new_n241), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n248), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n263), .A2(G97), .A3(new_n365), .A4(new_n507), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n252), .A2(new_n510), .A3(new_n254), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n616), .A2(new_n617), .A3(new_n303), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n619), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n627), .B2(new_n248), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n616), .A2(new_n294), .A3(new_n617), .ZN(new_n637));
  AOI21_X1  g0437(.A(G200), .B1(new_n616), .B2(new_n617), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n609), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  NOR4_X1   g0440(.A1(new_n481), .A2(new_n532), .A3(new_n570), .A4(new_n640), .ZN(G372));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n606), .A2(new_n608), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n584), .A2(new_n303), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n600), .B(new_n644), .C1(G169), .C2(new_n584), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n646), .B2(new_n635), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n616), .A2(new_n303), .A3(new_n617), .ZN(new_n648));
  AOI21_X1  g0448(.A(G169), .B1(new_n616), .B2(new_n617), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n648), .A2(new_n649), .A3(new_n636), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n609), .A2(new_n650), .A3(KEYINPUT26), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n647), .A2(new_n651), .B1(new_n600), .B2(new_n585), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT85), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n520), .B2(new_n522), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n521), .A2(new_n517), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(KEYINPUT85), .A3(new_n519), .A4(new_n518), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n361), .B1(new_n560), .B2(new_n561), .ZN(new_n659));
  INV_X1    g0459(.A(new_n562), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(G179), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n365), .B1(new_n540), .B2(new_n541), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n662), .A2(new_n543), .B1(new_n551), .B2(new_n553), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT86), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT86), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n555), .A2(new_n565), .A3(new_n665), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n654), .A2(new_n658), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n609), .A2(new_n569), .A3(new_n635), .A4(new_n639), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n652), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n481), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n468), .A2(new_n359), .A3(new_n380), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n478), .A2(new_n479), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n431), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n363), .A2(new_n376), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n299), .B(new_n302), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n305), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(G369));
  NAND3_X1  g0481(.A1(new_n250), .A2(new_n243), .A3(G13), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n524), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n654), .A2(new_n658), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n532), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n566), .A2(new_n688), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n554), .A2(new_n544), .B1(new_n563), .B2(new_n564), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n687), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT88), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n566), .A2(new_n569), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n555), .A2(new_n687), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n694), .A2(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n664), .A2(new_n666), .A3(new_n688), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n696), .A2(new_n697), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n523), .A2(new_n687), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(G399));
  NAND3_X1  g0512(.A1(new_n592), .A2(new_n397), .A3(new_n505), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT89), .Z(new_n714));
  NAND2_X1  g0514(.A1(new_n206), .A2(new_n281), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n714), .A2(new_n250), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n210), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT28), .Z(new_n719));
  INV_X1    g0519(.A(KEYINPUT93), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n489), .A2(G179), .A3(new_n503), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n616), .A2(new_n617), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n559), .A2(new_n277), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n502), .A2(G264), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n575), .A3(new_n725), .A4(new_n582), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT90), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT90), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n560), .A2(new_n584), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT91), .B1(new_n723), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n489), .A2(new_n503), .A3(G179), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n618), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT91), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n729), .A4(new_n727), .ZN(new_n735));
  XOR2_X1   g0535(.A(KEYINPUT92), .B(KEYINPUT30), .Z(new_n736));
  NAND3_X1  g0536(.A1(new_n731), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n584), .A2(G179), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n504), .A2(new_n618), .A3(new_n738), .A4(new_n562), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n721), .A2(new_n727), .A3(new_n722), .A4(new_n729), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n688), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n720), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NOR4_X1   g0545(.A1(new_n532), .A2(new_n640), .A3(new_n570), .A4(new_n687), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n687), .ZN(new_n748));
  INV_X1    g0548(.A(new_n744), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n737), .B2(new_n741), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n748), .A2(new_n743), .B1(new_n750), .B2(new_n720), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n646), .A2(new_n635), .A3(new_n642), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT26), .B1(new_n609), .B2(new_n650), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n645), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n695), .A2(new_n520), .A3(new_n522), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n668), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n688), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT29), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n669), .A2(new_n761), .A3(new_n688), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n719), .B1(new_n765), .B2(G1), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT94), .ZN(G364));
  NAND2_X1  g0567(.A1(new_n243), .A2(G13), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n250), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n716), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n691), .B2(G330), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n691), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n271), .A2(new_n206), .ZN(new_n775));
  INV_X1    g0575(.A(G355), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n776), .B1(G116), .B2(new_n206), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n236), .A2(new_n282), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n330), .A2(new_n206), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n282), .B2(new_n210), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n211), .B1(G20), .B2(new_n361), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n772), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n294), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n243), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n510), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n243), .A2(new_n303), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n792), .A2(G190), .A3(new_n356), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n271), .B1(new_n794), .B2(new_n202), .C1(new_n321), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n792), .A2(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G190), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n791), .B(new_n796), .C1(G68), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(new_n294), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n243), .A2(G179), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n793), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n806));
  OAI22_X1  g0606(.A1(new_n801), .A2(new_n258), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n393), .A2(G190), .A3(new_n802), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G87), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n393), .A2(new_n294), .A3(new_n802), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G107), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n799), .A2(new_n808), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n798), .ZN(new_n816));
  OR2_X1    g0616(.A1(KEYINPUT33), .A2(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(KEYINPUT33), .A2(G317), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G326), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n801), .A2(new_n820), .B1(new_n821), .B2(new_n790), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n813), .A2(G283), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  INV_X1    g0625(.A(G329), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n794), .A2(new_n825), .B1(new_n803), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n795), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n271), .B(new_n827), .C1(G322), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n810), .A2(G303), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n823), .A2(new_n824), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n815), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n788), .B1(new_n832), .B2(new_n785), .ZN(new_n833));
  INV_X1    g0633(.A(new_n784), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n691), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n774), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  AOI211_X1 g0637(.A(KEYINPUT98), .B(new_n429), .C1(new_n415), .C2(new_n418), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT98), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n422), .B2(new_n430), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n410), .B1(new_n409), .B2(new_n414), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT70), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n687), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT99), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT99), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n422), .A2(new_n846), .A3(new_n687), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n841), .A2(new_n848), .A3(new_n421), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n431), .B2(new_n688), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n670), .B2(new_n687), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n687), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n669), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n772), .B1(new_n855), .B2(new_n753), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n753), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n785), .A2(new_n782), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n330), .B1(new_n809), .B2(new_n387), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT96), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n816), .A2(new_n862), .B1(new_n510), .B2(new_n790), .ZN(new_n863));
  INV_X1    g0663(.A(new_n794), .ZN(new_n864));
  INV_X1    g0664(.A(new_n803), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G116), .A2(new_n864), .B1(new_n865), .B2(G311), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n866), .B1(new_n821), .B2(new_n795), .C1(new_n397), .C2(new_n812), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n863), .B(new_n867), .C1(G303), .C2(new_n800), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n828), .A2(G143), .B1(new_n864), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(G150), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n869), .B1(new_n816), .B2(new_n870), .C1(new_n871), .C2(new_n801), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT34), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n813), .A2(G68), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n810), .A2(G50), .ZN(new_n875));
  INV_X1    g0675(.A(new_n790), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(G58), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n330), .B1(new_n865), .B2(G132), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n874), .A2(new_n875), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n861), .A2(new_n868), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n785), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n772), .B1(G77), .B2(new_n859), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT97), .Z(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n783), .B2(new_n850), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n857), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(G384));
  NOR2_X1   g0686(.A1(new_n841), .A2(new_n687), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n669), .B2(new_n853), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT101), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n442), .A2(new_n688), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n674), .A2(new_n468), .A3(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n479), .B(new_n687), .C1(new_n478), .C2(new_n469), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n894), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n469), .B(new_n891), .C1(new_n478), .C2(new_n479), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT101), .B1(new_n899), .B2(new_n888), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT102), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n320), .B2(new_n338), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n333), .A2(KEYINPUT102), .A3(new_n366), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n337), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n248), .A3(new_n369), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n685), .B1(new_n905), .B2(new_n309), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n381), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n340), .B1(new_n327), .B2(new_n335), .ZN(new_n908));
  INV_X1    g0708(.A(new_n685), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n908), .A2(new_n364), .B1(new_n362), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n370), .A2(new_n379), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n905), .A2(new_n309), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n375), .A2(new_n685), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(new_n370), .B2(new_n379), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n913), .B1(new_n916), .B2(new_n911), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n907), .A2(new_n917), .A3(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT103), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT103), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n907), .A2(new_n917), .A3(new_n920), .A4(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n907), .A2(new_n917), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n919), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n896), .A2(new_n900), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n478), .A2(new_n479), .A3(new_n688), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n309), .A2(new_n905), .B1(new_n375), .B2(new_n685), .ZN(new_n929));
  INV_X1    g0729(.A(new_n912), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT37), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(new_n913), .B1(new_n381), .B2(new_n906), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n921), .B1(KEYINPUT38), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n920), .B1(new_n932), .B2(KEYINPUT38), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT39), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n368), .A2(new_n369), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n375), .A2(new_n685), .B1(new_n937), .B2(new_n309), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT37), .B1(new_n938), .B2(KEYINPUT104), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n910), .A2(new_n912), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n910), .A2(KEYINPUT104), .A3(KEYINPUT37), .A4(new_n912), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n370), .A2(new_n685), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT105), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n370), .A2(KEYINPUT17), .A3(new_n379), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT17), .B1(new_n370), .B2(new_n379), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n359), .A2(KEYINPUT105), .A3(new_n380), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n676), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n943), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n936), .B(new_n918), .C1(new_n951), .C2(KEYINPUT38), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n928), .B1(new_n935), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n676), .A2(new_n909), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n927), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n763), .A2(new_n481), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n679), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n955), .B(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n918), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n950), .A2(new_n944), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT104), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n910), .A2(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n962), .A2(KEYINPUT37), .B1(new_n912), .B2(new_n910), .ZN(new_n963));
  INV_X1    g0763(.A(new_n942), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n959), .B1(new_n966), .B2(new_n923), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n640), .A2(new_n570), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n968), .A2(new_n531), .A3(new_n523), .A4(new_n688), .ZN(new_n969));
  INV_X1    g0769(.A(new_n750), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n688), .B1(new_n737), .B2(new_n741), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n970), .C1(KEYINPUT31), .C2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n895), .A2(new_n972), .A3(new_n850), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT40), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n746), .A2(new_n750), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n748), .A2(new_n743), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n851), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT40), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n925), .A2(new_n977), .A3(new_n978), .A4(new_n895), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n972), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n481), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n980), .A2(new_n982), .ZN(new_n985));
  INV_X1    g0785(.A(G330), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n958), .A2(new_n988), .B1(G1), .B2(new_n768), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n958), .B2(new_n988), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n211), .A2(new_n243), .A3(new_n505), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n625), .B(KEYINPUT100), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT35), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT36), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n210), .B(G77), .C1(new_n321), .C2(new_n311), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n258), .A2(G68), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n250), .B(G13), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n990), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT106), .Z(G367));
  AND3_X1   g0803(.A1(new_n227), .A2(new_n206), .A3(new_n330), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n588), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n786), .B1(new_n1005), .B2(new_n206), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n772), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n821), .A2(new_n816), .B1(new_n801), .B2(new_n825), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G107), .B2(new_n876), .ZN(new_n1009));
  INV_X1    g0809(.A(G303), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n330), .B1(new_n795), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n794), .A2(new_n862), .B1(new_n803), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(new_n813), .C2(G97), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT46), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n809), .B2(new_n505), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n810), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1009), .A2(new_n1014), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n790), .A2(new_n311), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n804), .B2(new_n816), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G143), .B2(new_n800), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n330), .B1(new_n813), .B2(G77), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT111), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n795), .A2(new_n870), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT112), .B(G137), .Z(new_n1026));
  OAI22_X1  g0826(.A1(new_n1026), .A2(new_n803), .B1(new_n794), .B2(new_n258), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(new_n810), .C2(G58), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1022), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1023), .A2(KEYINPUT111), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1018), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1007), .B1(new_n1032), .B2(new_n785), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n609), .B1(new_n606), .B2(new_n688), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n645), .A2(new_n606), .A3(new_n688), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1033), .B1(new_n834), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT113), .Z(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n715), .B(KEYINPUT41), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n702), .A2(KEYINPUT110), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n648), .A2(new_n649), .A3(new_n636), .A4(new_n688), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(KEYINPUT107), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n635), .B(new_n639), .C1(new_n636), .C2(new_n688), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(KEYINPUT107), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT109), .B1(new_n711), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT109), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n710), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n701), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1050), .B(new_n1051), .C1(new_n1053), .C2(new_n705), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1049), .A2(new_n1054), .A3(KEYINPUT44), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n709), .A2(new_n710), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(new_n704), .A3(new_n1048), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n711), .A2(KEYINPUT45), .A3(new_n1048), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT44), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1042), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT44), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1067), .A2(new_n1041), .A3(new_n1061), .A4(new_n1055), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n701), .A2(new_n1052), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1070), .A2(new_n692), .A3(new_n1053), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1056), .A2(new_n1069), .B1(new_n691), .B2(G330), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n764), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1064), .A2(new_n1068), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1040), .B1(new_n1076), .B2(new_n765), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n771), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1048), .A2(new_n709), .A3(new_n710), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT108), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT108), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1053), .A2(new_n1081), .A3(new_n1048), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT42), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT42), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1080), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n635), .B1(new_n1051), .B2(new_n566), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n688), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1036), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT43), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1036), .A2(KEYINPUT43), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n703), .A2(new_n1051), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1083), .A2(KEYINPUT42), .B1(new_n688), .B2(new_n1087), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1096), .A2(new_n1091), .A3(new_n1090), .A4(new_n1086), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1039), .B1(new_n1078), .B2(new_n1100), .ZN(G387));
  NAND2_X1  g0901(.A1(new_n1074), .A2(new_n764), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n765), .A2(new_n1073), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n716), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n714), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1105), .A2(new_n775), .B1(G107), .B2(new_n206), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n232), .A2(G45), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT114), .Z(new_n1108));
  AOI211_X1 g0908(.A(G45), .B(new_n714), .C1(G68), .C2(G77), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n244), .A2(G50), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT50), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n779), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1106), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n772), .B1(new_n1113), .B2(new_n787), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n828), .A2(G317), .B1(new_n864), .B2(G303), .ZN(new_n1115));
  INV_X1    g0915(.A(G322), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1115), .B1(new_n816), .B2(new_n825), .C1(new_n1116), .C2(new_n801), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT48), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n810), .A2(G294), .B1(G283), .B2(new_n876), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT49), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n330), .B1(new_n820), .B2(new_n803), .C1(new_n812), .C2(new_n505), .ZN(new_n1126));
  OR3_X1    g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n330), .B1(new_n865), .B2(G150), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n258), .B2(new_n795), .C1(new_n311), .C2(new_n794), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n588), .A2(new_n876), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n510), .B2(new_n812), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n804), .A2(new_n801), .B1(new_n816), .B2(new_n244), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n809), .A2(new_n202), .ZN(new_n1133));
  OR4_X1    g0933(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n881), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1114), .B(new_n1135), .C1(new_n701), .C2(new_n784), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1073), .B2(new_n771), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1104), .A2(new_n1137), .ZN(G393));
  NAND4_X1  g0938(.A1(new_n1067), .A2(new_n703), .A3(new_n1061), .A4(new_n1055), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT115), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1142), .A2(KEYINPUT115), .A3(new_n703), .A4(new_n1067), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1067), .A2(new_n1061), .A3(new_n1055), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n702), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1103), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1103), .B1(new_n1144), .B2(new_n1042), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n715), .B1(new_n1148), .B2(new_n1068), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .A4(new_n771), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n786), .B1(new_n510), .B2(new_n206), .C1(new_n239), .C2(new_n779), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n772), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT116), .Z(new_n1154));
  OAI21_X1  g0954(.A(new_n814), .B1(new_n862), .B2(new_n809), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n330), .B1(new_n803), .B2(new_n1116), .C1(new_n821), .C2(new_n794), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n816), .A2(new_n1010), .B1(new_n505), .B2(new_n790), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n801), .A2(new_n1012), .B1(new_n825), .B2(new_n795), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT52), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n801), .A2(new_n870), .B1(new_n804), .B2(new_n795), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT51), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n790), .A2(new_n202), .ZN(new_n1163));
  INV_X1    g0963(.A(G143), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n271), .B1(new_n803), .B2(new_n1164), .C1(new_n244), .C2(new_n794), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G50), .C2(new_n798), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G68), .A2(new_n810), .B1(new_n813), .B2(G87), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1158), .A2(new_n1160), .B1(new_n1162), .B2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1154), .B1(new_n1169), .B2(new_n881), .C1(new_n1048), .C2(new_n834), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1151), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1150), .A2(new_n1171), .ZN(G390));
  AOI21_X1  g0972(.A(KEYINPUT38), .B1(new_n960), .B2(new_n965), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n928), .B1(new_n1173), .B2(new_n959), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n841), .A2(new_n421), .A3(new_n848), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1176), .B(new_n688), .C1(new_n756), .C2(new_n758), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n887), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT117), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(KEYINPUT117), .A3(new_n1178), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n895), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1175), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n928), .B1(new_n899), .B2(new_n888), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n935), .A2(new_n1184), .A3(new_n952), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n986), .B1(new_n747), .B2(new_n751), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n850), .A3(new_n895), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n972), .A2(G330), .A3(new_n850), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(new_n899), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1189), .A2(new_n1193), .A3(new_n770), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n935), .A2(new_n952), .A3(new_n782), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n772), .B1(new_n406), .B2(new_n859), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n800), .A2(G128), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n816), .B2(new_n1026), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G159), .B2(new_n876), .ZN(new_n1199));
  INV_X1    g0999(.A(G132), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n795), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT54), .B(G143), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n271), .B1(new_n794), .B2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(G125), .C2(new_n865), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1199), .B(new_n1204), .C1(new_n258), .C2(new_n812), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n810), .A2(G150), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT53), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1163), .B1(G283), .B2(new_n800), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n387), .B2(new_n816), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n795), .A2(new_n505), .B1(new_n803), .B2(new_n821), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n271), .B(new_n1210), .C1(G97), .C2(new_n864), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n811), .A3(new_n874), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1205), .A2(new_n1207), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1196), .B1(new_n1213), .B2(new_n785), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1194), .B1(new_n1195), .B2(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n935), .A2(new_n1184), .A3(new_n952), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1177), .A2(KEYINPUT117), .A3(new_n1178), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(new_n1179), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1174), .B1(new_n1218), .B2(new_n895), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1191), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n895), .B1(new_n1186), .B2(new_n850), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n889), .B1(new_n1221), .B2(new_n1191), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1190), .A2(new_n899), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1187), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n981), .A2(new_n481), .A3(new_n986), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n956), .A2(new_n1227), .A3(new_n679), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1220), .A2(new_n1226), .A3(new_n1188), .A4(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(KEYINPUT118), .A3(new_n716), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT118), .B1(new_n1229), .B2(new_n716), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1215), .B1(new_n1233), .B2(new_n1234), .ZN(G378));
  AOI22_X1  g1035(.A1(new_n798), .A2(G132), .B1(new_n864), .B2(G137), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT120), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G125), .A2(new_n800), .B1(new_n828), .B2(G128), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n870), .B2(new_n790), .C1(new_n809), .C2(new_n1202), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n813), .A2(G159), .ZN(new_n1243));
  AOI211_X1 g1043(.A(G33), .B(G41), .C1(new_n865), .C2(G124), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT59), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n1240), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n813), .A2(G58), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1005), .B2(new_n794), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1020), .B1(new_n816), .B2(new_n510), .C1(new_n505), .C2(new_n801), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n271), .A2(G41), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n862), .B2(new_n803), .C1(new_n387), .C2(new_n795), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1252), .A4(new_n1133), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n258), .B1(G33), .B2(G41), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1253), .A2(KEYINPUT58), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT119), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1247), .B(new_n1256), .C1(KEYINPUT58), .C2(new_n1253), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n772), .B1(G50), .B2(new_n859), .C1(new_n1257), .C2(new_n881), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n306), .A2(new_n266), .A3(new_n909), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n266), .A2(new_n909), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n299), .A2(new_n302), .A3(new_n305), .A4(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1258), .B1(new_n782), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n980), .A2(G330), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1265), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1265), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n980), .A2(G330), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n955), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n953), .A2(new_n954), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n926), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1269), .B1(new_n980), .B2(G330), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n986), .B(new_n1265), .C1(new_n974), .C2(new_n979), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1266), .B1(new_n1277), .B2(new_n771), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1229), .A2(new_n1228), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(KEYINPUT57), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n716), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1278), .B1(new_n1281), .B2(new_n1282), .ZN(G375));
  AND2_X1   g1083(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1228), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1040), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1231), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n899), .A2(new_n782), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n772), .B1(G68), .B2(new_n859), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n505), .A2(new_n816), .B1(new_n801), .B2(new_n821), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n330), .B1(new_n803), .B2(new_n1010), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n795), .A2(new_n862), .B1(new_n794), .B2(new_n387), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n813), .A2(G77), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n810), .A2(G97), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1130), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1248), .A2(new_n271), .ZN(new_n1298));
  XOR2_X1   g1098(.A(new_n1298), .B(KEYINPUT121), .Z(new_n1299));
  AOI22_X1  g1099(.A1(G150), .A2(new_n864), .B1(new_n865), .B2(G128), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n795), .B2(new_n1026), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(G159), .B2(new_n810), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(G50), .A2(new_n876), .B1(new_n800), .B2(G132), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1302), .B(new_n1303), .C1(new_n816), .C2(new_n1202), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1297), .B1(new_n1299), .B2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1290), .B1(new_n1305), .B2(new_n785), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1226), .A2(new_n771), .B1(new_n1289), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1288), .A2(new_n1307), .ZN(G381));
  INV_X1    g1108(.A(G375), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1309), .A2(KEYINPUT122), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(KEYINPUT122), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n764), .B1(new_n1148), .B2(new_n1068), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n770), .B1(new_n1312), .B2(new_n1040), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1038), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(G378), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1151), .A2(new_n1170), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1318));
  NOR4_X1   g1118(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1319));
  AND4_X1   g1119(.A1(new_n1315), .A2(new_n1316), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1310), .A2(new_n1311), .A3(new_n1320), .ZN(G407));
  NAND2_X1  g1121(.A1(new_n686), .A2(G213), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1310), .A2(new_n1316), .A3(new_n1311), .A4(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1324), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1125(.A1(new_n1323), .A2(G2897), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1284), .A2(KEYINPUT60), .A3(new_n1285), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1328), .A2(new_n716), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1231), .A2(KEYINPUT60), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1286), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(G384), .B1(new_n1332), .B2(new_n1307), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1307), .ZN(new_n1334));
  AOI211_X1 g1134(.A(new_n885), .B(new_n1334), .C1(new_n1329), .C2(new_n1331), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1327), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1328), .A2(new_n716), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1337), .B1(new_n1286), .B2(new_n1330), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n885), .B1(new_n1338), .B2(new_n1334), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1332), .A2(G384), .A3(new_n1307), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1326), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1336), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  OAI211_X1 g1143(.A(G378), .B(new_n1278), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1277), .A2(new_n1287), .A3(new_n1279), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1278), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1234), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(new_n1232), .A3(new_n1230), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(new_n1348), .A3(new_n1215), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1344), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1322), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT61), .B1(new_n1343), .B2(new_n1351), .ZN(new_n1352));
  XOR2_X1   g1152(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1353));
  NOR2_X1   g1153(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1353), .B1(new_n1351), .B2(new_n1355), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(G393), .B(new_n836), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(G387), .A2(new_n1318), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1314), .B1(new_n1077), .B2(new_n771), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(G390), .A2(KEYINPUT124), .A3(new_n1359), .A4(new_n1039), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1358), .A2(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(KEYINPUT124), .B1(new_n1315), .B2(G390), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1357), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1357), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1364), .B1(G387), .B2(new_n1318), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1315), .A2(G390), .ZN(new_n1366));
  NOR3_X1   g1166(.A1(new_n1365), .A2(new_n1366), .A3(KEYINPUT125), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT125), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1357), .B1(new_n1315), .B2(G390), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1368), .B1(new_n1369), .B2(new_n1358), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1363), .B1(new_n1367), .B2(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1323), .B1(new_n1344), .B2(new_n1349), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1372), .A2(KEYINPUT63), .A3(new_n1354), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1352), .A2(new_n1356), .A3(new_n1371), .A4(new_n1373), .ZN(new_n1374));
  XOR2_X1   g1174(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1375));
  AND3_X1   g1175(.A1(new_n1372), .A2(new_n1354), .A3(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT61), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1377), .B1(new_n1372), .B2(new_n1342), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1379), .B1(new_n1372), .B2(new_n1354), .ZN(new_n1380));
  NOR3_X1   g1180(.A1(new_n1376), .A2(new_n1378), .A3(new_n1380), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1374), .B1(new_n1381), .B2(new_n1371), .ZN(G405));
  NAND2_X1  g1182(.A1(new_n1354), .A2(KEYINPUT127), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(G375), .A2(new_n1316), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1383), .A2(new_n1384), .A3(new_n1344), .ZN(new_n1385));
  OAI21_X1  g1185(.A(KEYINPUT125), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1369), .A2(new_n1368), .A3(new_n1358), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1388));
  NOR2_X1   g1188(.A1(new_n1354), .A2(KEYINPUT127), .ZN(new_n1389));
  INV_X1    g1189(.A(new_n1389), .ZN(new_n1390));
  AND3_X1   g1190(.A1(new_n1388), .A2(new_n1363), .A3(new_n1390), .ZN(new_n1391));
  AOI21_X1  g1191(.A(new_n1390), .B1(new_n1388), .B2(new_n1363), .ZN(new_n1392));
  OAI21_X1  g1192(.A(new_n1385), .B1(new_n1391), .B2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1371), .A2(new_n1389), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1385), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1388), .A2(new_n1363), .A3(new_n1390), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1394), .A2(new_n1395), .A3(new_n1396), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1393), .A2(new_n1397), .ZN(G402));
endmodule


