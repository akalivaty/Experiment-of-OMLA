//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT74), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G116), .B(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G116), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n197), .A2(new_n204), .A3(KEYINPUT71), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT71), .B1(new_n197), .B2(new_n204), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT64), .A2(G143), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT64), .A2(G143), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n209), .B1(new_n212), .B2(new_n208), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT0), .B(G128), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT65), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT64), .A2(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n217), .B1(new_n222), .B2(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT0), .A3(G128), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n208), .A3(new_n221), .ZN(new_n225));
  INV_X1    g039(.A(new_n209), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  INV_X1    g042(.A(new_n214), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n215), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT66), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G134), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT11), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n233), .A3(G134), .ZN(new_n238));
  AOI211_X1 g052(.A(G131), .B(new_n234), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(G137), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n215), .A2(new_n224), .A3(new_n246), .A4(new_n230), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n232), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n233), .A2(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n234), .B2(KEYINPUT67), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n242), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(G131), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n241), .A2(new_n240), .A3(new_n242), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n258), .B(KEYINPUT1), .C1(new_n219), .C2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n262), .B2(new_n213), .ZN(new_n263));
  OAI21_X1  g077(.A(G146), .B1(new_n210), .B2(new_n211), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(G128), .A4(new_n216), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n227), .B(KEYINPUT70), .C1(new_n261), .C2(new_n260), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n256), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n207), .B1(new_n248), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n205), .A2(new_n206), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n202), .A2(new_n203), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n195), .A2(new_n196), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n197), .A2(new_n204), .A3(KEYINPUT71), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT73), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n255), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(KEYINPUT65), .B(new_n214), .C1(new_n225), .C2(new_n226), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n237), .B1(G134), .B2(new_n233), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n235), .A2(KEYINPUT11), .A3(G137), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n242), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n254), .A3(KEYINPUT72), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n239), .B2(new_n243), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n285), .A2(new_n224), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n280), .A2(new_n282), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT28), .B1(new_n271), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n280), .A2(new_n282), .A3(new_n293), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G237), .ZN(new_n300));
  INV_X1    g114(.A(G953), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(G210), .ZN(new_n302));
  INV_X1    g116(.A(G101), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n190), .B1(new_n299), .B2(new_n307), .ZN(new_n308));
  AOI211_X1 g122(.A(KEYINPUT74), .B(new_n306), .C1(new_n295), .C2(new_n298), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT30), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n248), .A2(new_n311), .A3(new_n270), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n268), .A2(new_n281), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n292), .A2(new_n290), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(new_n231), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT30), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n207), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n294), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n306), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT31), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(KEYINPUT31), .A3(new_n306), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI211_X1 g138(.A(KEYINPUT75), .B(new_n189), .C1(new_n310), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n248), .A2(new_n270), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n318), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n297), .B1(new_n328), .B2(new_n296), .ZN(new_n329));
  INV_X1    g143(.A(new_n298), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n307), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n299), .A2(new_n190), .A3(new_n307), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT31), .B1(new_n319), .B2(new_n306), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n319), .A2(KEYINPUT31), .A3(new_n306), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n332), .B(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n326), .B1(new_n336), .B2(new_n188), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n187), .B1(new_n325), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n319), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT29), .B1(new_n339), .B2(new_n307), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n307), .B2(new_n299), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n280), .B1(new_n282), .B2(new_n293), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n294), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n330), .B1(new_n343), .B2(KEYINPUT28), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT29), .A3(new_n306), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  INV_X1    g160(.A(G902), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT29), .A4(new_n306), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n341), .A2(new_n346), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n189), .B1(new_n310), .B2(new_n324), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n350), .A2(G472), .B1(new_n351), .B2(KEYINPUT32), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G214), .B1(G237), .B2(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G224), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT7), .B1(new_n356), .B2(G953), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n231), .A2(G125), .ZN(new_n359));
  INV_X1    g173(.A(G125), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n263), .A2(new_n360), .A3(new_n266), .A4(new_n267), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n361), .A3(new_n358), .ZN(new_n365));
  INV_X1    g179(.A(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G107), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(G107), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n366), .B2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G104), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n371), .A2(new_n374), .A3(new_n303), .A4(new_n367), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT85), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n196), .A2(KEYINPUT5), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(KEYINPUT5), .B2(new_n199), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n197), .B1(new_n380), .B2(new_n191), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n378), .B(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(G110), .B(G122), .Z(new_n383));
  XOR2_X1   g197(.A(new_n383), .B(KEYINPUT8), .Z(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n364), .A2(KEYINPUT87), .A3(new_n365), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n362), .A2(new_n363), .ZN(new_n387));
  AOI211_X1 g201(.A(KEYINPUT86), .B(new_n358), .C1(new_n359), .C2(new_n361), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n365), .B(new_n385), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n371), .A2(new_n374), .A3(new_n367), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n375), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(G101), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n207), .A2(new_n397), .B1(new_n381), .B2(new_n376), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n398), .A2(new_n383), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n386), .A2(new_n391), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(KEYINPUT84), .A3(new_n383), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n402), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n359), .A2(new_n361), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n356), .A2(G953), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n400), .A2(new_n347), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G210), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n400), .A2(new_n347), .A3(new_n411), .A4(new_n409), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n355), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G475), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n360), .A2(KEYINPUT16), .A3(G140), .ZN(new_n417));
  OR2_X1    g231(.A1(G125), .A2(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(G125), .A2(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n421), .A2(G146), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(G146), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n219), .A2(new_n300), .A3(new_n301), .A4(G214), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n300), .A2(new_n301), .A3(G214), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(G131), .B(new_n425), .C1(new_n427), .C2(new_n222), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT88), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n212), .A2(new_n426), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n430), .A2(new_n431), .A3(G131), .A4(new_n425), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n432), .A3(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n432), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n425), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n240), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n424), .B(new_n433), .C1(new_n437), .C2(KEYINPUT17), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n366), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n435), .B1(new_n441), .B2(new_n240), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n420), .B(new_n208), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n442), .B(new_n443), .C1(new_n441), .C2(new_n428), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n438), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT19), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT89), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n446), .A2(KEYINPUT89), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n420), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n418), .A2(KEYINPUT89), .A3(new_n446), .A4(new_n419), .ZN(new_n450));
  AOI21_X1  g264(.A(G146), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n452));
  OR3_X1    g266(.A1(new_n422), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n422), .B2(new_n451), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n437), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n440), .B1(new_n455), .B2(new_n444), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n416), .B(new_n347), .C1(new_n445), .C2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n440), .B1(new_n438), .B2(new_n444), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n347), .B1(new_n445), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G475), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(new_n444), .ZN(new_n463));
  INV_X1    g277(.A(new_n440), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n438), .A2(new_n440), .A3(new_n444), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n467), .A2(KEYINPUT20), .A3(new_n416), .A4(new_n347), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n459), .A2(new_n462), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n222), .A2(G128), .ZN(new_n470));
  INV_X1    g284(.A(G128), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G143), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(KEYINPUT13), .A3(new_n472), .ZN(new_n473));
  OR3_X1    g287(.A1(new_n212), .A2(KEYINPUT13), .A3(new_n471), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(G134), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n235), .A3(new_n472), .ZN(new_n478));
  XNOR2_X1  g292(.A(G116), .B(G122), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(new_n373), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT91), .A4(G134), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n470), .A2(new_n472), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G134), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n484), .A2(new_n478), .B1(new_n373), .B2(new_n479), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n200), .A2(KEYINPUT14), .A3(G122), .ZN(new_n486));
  INV_X1    g300(.A(new_n479), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(KEYINPUT14), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n373), .B2(new_n488), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT9), .B(G234), .Z(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(G217), .A3(new_n301), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n482), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n482), .B2(new_n489), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n347), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G478), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n469), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(G952), .A3(new_n301), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT21), .B(G898), .Z(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(G902), .A3(G953), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n415), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G217), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(G234), .B2(new_n347), .ZN(new_n508));
  INV_X1    g322(.A(new_n422), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n420), .A2(new_n208), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n471), .A2(G119), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n198), .A2(G128), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT24), .B(G110), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT78), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n198), .B2(G128), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n471), .A2(KEYINPUT23), .A3(G119), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(G110), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n509), .B(new_n510), .C1(new_n516), .C2(new_n521), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT77), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n520), .A2(new_n524), .A3(G110), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n520), .B2(G110), .ZN(new_n526));
  OAI221_X1 g340(.A(new_n523), .B1(new_n525), .B2(new_n526), .C1(new_n422), .C2(new_n423), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G137), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n301), .A2(G221), .A3(G234), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n529), .B(new_n530), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n527), .A3(new_n531), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n347), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n535), .A2(new_n537), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT79), .B1(new_n535), .B2(new_n537), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n508), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n534), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT80), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n508), .A2(G902), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G469), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n268), .A2(KEYINPUT10), .A3(new_n377), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n285), .A2(new_n396), .A3(new_n394), .A4(new_n224), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n471), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n266), .B1(new_n550), .B2(new_n223), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n377), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n548), .A2(new_n549), .A3(new_n314), .A4(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT83), .ZN(new_n556));
  XNOR2_X1  g370(.A(G110), .B(G140), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT82), .ZN(new_n558));
  INV_X1    g372(.A(G227), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G953), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n558), .B(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n555), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n556), .B1(new_n555), .B2(new_n561), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n263), .A2(new_n376), .A3(new_n266), .A4(new_n267), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n552), .ZN(new_n565));
  INV_X1    g379(.A(new_n314), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT12), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n568), .B(new_n244), .C1(new_n564), .C2(new_n552), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n562), .A2(new_n563), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n548), .A2(new_n549), .A3(new_n554), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n566), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n561), .B1(new_n573), .B2(new_n555), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n547), .B(new_n347), .C1(new_n571), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(G469), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n561), .ZN(new_n577));
  INV_X1    g391(.A(new_n555), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n555), .A3(new_n561), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(G469), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G221), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n490), .B2(new_n347), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT81), .Z(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n353), .A2(new_n506), .A3(new_n546), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n310), .B2(new_n324), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n336), .A2(new_n347), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT92), .ZN(new_n595));
  INV_X1    g409(.A(new_n337), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n351), .A2(new_n326), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n593), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n546), .A3(new_n587), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT93), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n413), .A2(new_n414), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n354), .ZN(new_n602));
  INV_X1    g416(.A(new_n505), .ZN(new_n603));
  INV_X1    g417(.A(new_n495), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n493), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT33), .B1(new_n494), .B2(new_n495), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(G478), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n497), .A2(new_n347), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n497), .B(new_n347), .C1(new_n494), .C2(new_n495), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n469), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n602), .A2(new_n603), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n600), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(new_n366), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  INV_X1    g433(.A(new_n469), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n499), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n415), .A2(new_n505), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n415), .A2(new_n625), .A3(new_n505), .A4(new_n622), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n600), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  OR2_X1    g443(.A1(new_n528), .A2(KEYINPUT96), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n528), .A2(KEYINPUT96), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n545), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n541), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n541), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n587), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n598), .A2(new_n506), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  OAI21_X1  g459(.A(new_n502), .B1(new_n504), .B2(G900), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n621), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT98), .B1(new_n602), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n415), .A2(new_n651), .A3(new_n648), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n353), .A2(new_n642), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XNOR2_X1  g468(.A(new_n601), .B(KEYINPUT38), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n646), .B(KEYINPUT39), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n587), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n469), .A2(new_n499), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n355), .B(new_n661), .C1(new_n658), .C2(KEYINPUT40), .ZN(new_n662));
  INV_X1    g476(.A(new_n636), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n319), .A2(new_n307), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n347), .B1(new_n343), .B2(new_n306), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n338), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n660), .A2(new_n662), .A3(new_n663), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n212), .ZN(G45));
  NAND3_X1  g484(.A1(new_n613), .A2(new_n469), .A3(new_n646), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n353), .A2(new_n415), .A3(new_n642), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n555), .A2(new_n561), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT83), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n567), .A2(new_n569), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n555), .A2(new_n556), .A3(new_n561), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n574), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n347), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n685), .A3(new_n347), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(G469), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n675), .B1(new_n687), .B2(new_n575), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n685), .B1(new_n682), .B2(new_n347), .ZN(new_n689));
  AOI211_X1 g503(.A(KEYINPUT99), .B(G902), .C1(new_n680), .C2(new_n681), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n690), .A3(new_n547), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(KEYINPUT100), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n688), .A2(new_n692), .A3(new_n584), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n353), .A2(new_n693), .A3(new_n546), .A4(new_n615), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND2_X1  g510(.A1(new_n353), .A2(new_n546), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n624), .A2(new_n626), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n688), .A2(new_n692), .ZN(new_n699));
  INV_X1    g513(.A(new_n584), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n200), .ZN(G18));
  NAND2_X1  g517(.A1(new_n500), .A2(new_n505), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n338), .B2(new_n352), .ZN(new_n705));
  INV_X1    g519(.A(new_n575), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT100), .B1(new_n691), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n687), .A2(new_n675), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n415), .A2(new_n707), .A3(new_n700), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n709), .A3(new_n640), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NAND2_X1  g525(.A1(new_n661), .A2(KEYINPUT101), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n469), .A2(new_n713), .A3(new_n499), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n415), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n603), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n594), .A2(G472), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n324), .B1(new_n306), .B2(new_n344), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n188), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n693), .A2(new_n717), .A3(new_n546), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND4_X1  g537(.A1(new_n707), .A2(new_n415), .A3(new_n700), .A4(new_n708), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n671), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n613), .A2(KEYINPUT102), .A3(new_n469), .A4(new_n646), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n718), .A3(new_n636), .A4(new_n720), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n360), .ZN(G27));
  XNOR2_X1  g545(.A(new_n576), .B(KEYINPUT103), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n575), .A2(new_n581), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n575), .A2(KEYINPUT104), .A3(new_n581), .A4(new_n732), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n735), .A2(new_n700), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n413), .A2(new_n354), .A3(new_n414), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n413), .A2(KEYINPUT105), .A3(new_n354), .A4(new_n414), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n546), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n743), .B1(new_n352), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n745), .A3(KEYINPUT42), .A4(new_n728), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n742), .A2(new_n353), .A3(new_n546), .A4(new_n728), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  INV_X1    g567(.A(new_n697), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n648), .A3(new_n742), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(new_n732), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n579), .A2(new_n580), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(G469), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(KEYINPUT107), .A3(G469), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n575), .B1(new_n764), .B2(KEYINPUT46), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n700), .B(new_n657), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n598), .A2(KEYINPUT108), .A3(new_n663), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n469), .A2(new_n612), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT43), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT108), .B1(new_n598), .B2(new_n663), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n767), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n740), .A2(new_n741), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n774), .B(new_n776), .C1(new_n773), .C2(new_n772), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  OAI21_X1  g592(.A(new_n700), .B1(new_n765), .B2(new_n766), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n775), .A2(new_n546), .A3(new_n671), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n338), .A3(new_n352), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  INV_X1    g598(.A(new_n502), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n770), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n693), .A2(new_n776), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT116), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n636), .A3(new_n721), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n701), .A2(new_n502), .A3(new_n775), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n668), .A2(new_n743), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n620), .A3(new_n612), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n787), .A2(new_n546), .A3(new_n721), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n355), .B1(KEYINPUT115), .B2(KEYINPUT50), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n655), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n693), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n699), .B(KEYINPUT109), .Z(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n585), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n776), .B(new_n795), .C1(new_n781), .C2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n794), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n789), .A2(new_n808), .A3(new_n745), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n789), .B2(new_n745), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT48), .ZN(new_n811));
  OR3_X1    g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n791), .A2(new_n792), .ZN(new_n813));
  OAI211_X1 g627(.A(G952), .B(new_n301), .C1(new_n813), .C2(new_n614), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n810), .B2(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n806), .A2(new_n807), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n735), .A2(new_n700), .A3(new_n736), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n716), .A2(new_n647), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n668), .A2(new_n819), .A3(new_n663), .ZN(new_n820));
  INV_X1    g634(.A(new_n729), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n709), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n653), .A2(new_n820), .A3(new_n673), .A4(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT112), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n602), .B(new_n641), .C1(new_n338), .C2(new_n352), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n730), .B1(new_n827), .B2(new_n672), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n653), .A4(new_n820), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n710), .A2(new_n588), .A3(new_n722), .A4(new_n643), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n614), .A2(KEYINPUT111), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n613), .A2(new_n837), .A3(new_n469), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n621), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n839), .A2(new_n415), .A3(new_n505), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n598), .A2(new_n840), .A3(new_n546), .A4(new_n587), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n694), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n835), .A2(new_n702), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n353), .A2(new_n500), .A3(new_n642), .A4(new_n646), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n821), .A2(new_n737), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n775), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n752), .A2(new_n843), .A3(new_n755), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT53), .B1(new_n834), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n752), .A2(new_n843), .A3(new_n755), .A4(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n830), .A2(new_n831), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n852));
  NOR3_X1   g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n834), .A2(new_n848), .A3(KEYINPUT53), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n855), .A2(KEYINPUT114), .A3(new_n856), .A4(new_n857), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n817), .A2(new_n854), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n795), .A2(new_n709), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n862), .A2(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n801), .A2(KEYINPUT49), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT110), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n656), .A2(new_n585), .A3(new_n769), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n801), .B2(KEYINPUT49), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n668), .A2(new_n355), .A3(new_n743), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n870), .ZN(G75));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n347), .B1(new_n855), .B2(new_n857), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT56), .B1(new_n873), .B2(G210), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n405), .B(new_n408), .Z(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT55), .Z(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n755), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n747), .A2(new_n749), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n883), .B2(new_n746), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n835), .A2(new_n846), .A3(new_n702), .A4(new_n842), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n832), .B1(new_n830), .B2(new_n831), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n857), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n890), .A2(G210), .A3(G902), .ZN(new_n891));
  OAI211_X1 g705(.A(KEYINPUT118), .B(new_n876), .C1(new_n891), .C2(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n878), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n301), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(G902), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT119), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n873), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n412), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n877), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n893), .A2(new_n895), .A3(new_n902), .ZN(G51));
  NAND2_X1  g717(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n858), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n732), .B(KEYINPUT57), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n682), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n897), .A2(new_n762), .A3(new_n763), .A4(new_n899), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n894), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND2_X1  g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT120), .Z(new_n912));
  NAND3_X1  g726(.A1(new_n897), .A2(new_n899), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n466), .A3(new_n465), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n897), .A2(new_n467), .A3(new_n899), .A4(new_n912), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n914), .A2(new_n895), .A3(new_n915), .ZN(G60));
  NAND2_X1  g730(.A1(new_n606), .A2(new_n607), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n860), .A2(new_n854), .A3(new_n861), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n609), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n905), .A2(new_n917), .A3(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n894), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT60), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n855), .B2(new_n857), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n895), .B1(new_n927), .B2(new_n544), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n633), .A2(new_n634), .ZN(new_n929));
  INV_X1    g743(.A(new_n926), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n890), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n932), .B2(KEYINPUT61), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n890), .A2(new_n929), .A3(new_n930), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n934), .B(new_n895), .C1(new_n544), .C2(new_n927), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(KEYINPUT123), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n936), .C1(new_n928), .C2(new_n931), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n935), .B2(new_n936), .ZN(new_n941));
  OAI22_X1  g755(.A1(new_n933), .A2(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G66));
  AOI21_X1  g756(.A(new_n301), .B1(new_n503), .B2(G224), .ZN(new_n943));
  INV_X1    g757(.A(new_n843), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n301), .ZN(new_n945));
  INV_X1    g759(.A(G898), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n405), .B1(new_n946), .B2(G953), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  NOR2_X1   g762(.A1(new_n301), .A2(G900), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n559), .B2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT127), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n449), .A2(new_n450), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n317), .B(new_n953), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n777), .A2(new_n783), .ZN(new_n956));
  INV_X1    g770(.A(new_n828), .ZN(new_n957));
  INV_X1    g771(.A(new_n653), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT124), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n828), .A2(new_n960), .A3(new_n653), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n669), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n775), .A2(new_n658), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n754), .A2(new_n839), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n963), .A2(new_n964), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n962), .B2(new_n965), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n956), .A2(new_n966), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n955), .B1(new_n971), .B2(new_n301), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n777), .A2(new_n783), .A3(new_n959), .A4(new_n961), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n745), .A2(new_n415), .A3(new_n715), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n884), .B1(new_n767), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n301), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n949), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n977), .A2(KEYINPUT126), .A3(new_n978), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n952), .B(new_n973), .C1(new_n983), .C2(new_n954), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n954), .B1(new_n981), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n951), .B1(new_n985), .B2(new_n972), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n971), .B2(new_n944), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n894), .B1(new_n990), .B2(new_n665), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n339), .A2(new_n306), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n974), .A2(new_n944), .A3(new_n976), .ZN(new_n993));
  INV_X1    g807(.A(new_n989), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n992), .A2(new_n665), .A3(new_n994), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n849), .B2(new_n853), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n991), .A2(new_n995), .A3(new_n997), .ZN(G57));
endmodule


