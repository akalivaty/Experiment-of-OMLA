

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G2105), .A2(n527), .ZN(n987) );
  OR2_X1 U554 ( .A1(n798), .A2(n797), .ZN(n520) );
  OR2_X1 U555 ( .A1(n789), .A2(n788), .ZN(n521) );
  NOR2_X1 U556 ( .A1(n752), .A2(n751), .ZN(n754) );
  INV_X1 U557 ( .A(KEYINPUT91), .ZN(n714) );
  AND2_X1 U558 ( .A1(n771), .A2(n770), .ZN(n772) );
  INV_X1 U559 ( .A(KEYINPUT64), .ZN(n779) );
  NAND2_X1 U560 ( .A1(G160), .A2(n713), .ZN(n725) );
  AND2_X1 U561 ( .A1(n799), .A2(n520), .ZN(n800) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n650) );
  NOR2_X1 U563 ( .A1(G651), .A2(n623), .ZN(n645) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n522), .Z(n985) );
  NAND2_X1 U566 ( .A1(G137), .A2(n985), .ZN(n523) );
  XNOR2_X1 U567 ( .A(n523), .B(KEYINPUT66), .ZN(n526) );
  INV_X1 U568 ( .A(G2104), .ZN(n527) );
  NAND2_X1 U569 ( .A1(G101), .A2(n987), .ZN(n524) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n524), .Z(n525) );
  NAND2_X1 U571 ( .A1(n526), .A2(n525), .ZN(n532) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n981) );
  NAND2_X1 U573 ( .A1(G113), .A2(n981), .ZN(n530) );
  NAND2_X1 U574 ( .A1(n527), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U575 ( .A(n528), .B(KEYINPUT65), .ZN(n982) );
  NAND2_X1 U576 ( .A1(G125), .A2(n982), .ZN(n529) );
  NAND2_X1 U577 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X2 U578 ( .A1(n532), .A2(n531), .ZN(G160) );
  NAND2_X1 U579 ( .A1(G90), .A2(n650), .ZN(n535) );
  XNOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .ZN(n533) );
  XNOR2_X1 U581 ( .A(n533), .B(KEYINPUT67), .ZN(n623) );
  INV_X1 U582 ( .A(G651), .ZN(n538) );
  NOR2_X1 U583 ( .A1(n623), .A2(n538), .ZN(n651) );
  NAND2_X1 U584 ( .A1(G77), .A2(n651), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n537) );
  XOR2_X1 U586 ( .A(KEYINPUT9), .B(KEYINPUT69), .Z(n536) );
  XNOR2_X1 U587 ( .A(n537), .B(n536), .ZN(n543) );
  NOR2_X1 U588 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n539), .Z(n646) );
  NAND2_X1 U590 ( .A1(G64), .A2(n646), .ZN(n541) );
  NAND2_X1 U591 ( .A1(G52), .A2(n645), .ZN(n540) );
  AND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(G301) );
  INV_X1 U594 ( .A(G301), .ZN(G171) );
  INV_X1 U595 ( .A(G57), .ZN(G237) );
  NAND2_X1 U596 ( .A1(G138), .A2(n985), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G102), .A2(n987), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G114), .A2(n981), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G126), .A2(n982), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(G164) );
  XOR2_X1 U603 ( .A(KEYINPUT4), .B(KEYINPUT76), .Z(n551) );
  NAND2_X1 U604 ( .A1(G89), .A2(n650), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U606 ( .A(KEYINPUT75), .B(n552), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n651), .A2(G76), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT5), .ZN(n560) );
  NAND2_X1 U610 ( .A1(G63), .A2(n646), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G51), .A2(n645), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U615 ( .A(n561), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G94), .A2(G452), .ZN(n562) );
  XOR2_X1 U618 ( .A(KEYINPUT70), .B(n562), .Z(G173) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n563) );
  XOR2_X1 U620 ( .A(n563), .B(KEYINPUT10), .Z(n823) );
  NAND2_X1 U621 ( .A1(n823), .A2(G567), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  XOR2_X1 U623 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n566) );
  NAND2_X1 U624 ( .A1(G56), .A2(n646), .ZN(n565) );
  XNOR2_X1 U625 ( .A(n566), .B(n565), .ZN(n576) );
  NAND2_X1 U626 ( .A1(G43), .A2(n645), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n567), .B(KEYINPUT73), .ZN(n574) );
  NAND2_X1 U628 ( .A1(G81), .A2(n650), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n568), .B(KEYINPUT72), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G68), .A2(n651), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT13), .B(n572), .Z(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n900) );
  INV_X1 U636 ( .A(G860), .ZN(n596) );
  OR2_X1 U637 ( .A1(n900), .A2(n596), .ZN(G153) );
  NAND2_X1 U638 ( .A1(G301), .A2(G868), .ZN(n577) );
  XNOR2_X1 U639 ( .A(n577), .B(KEYINPUT74), .ZN(n586) );
  INV_X1 U640 ( .A(G868), .ZN(n666) );
  NAND2_X1 U641 ( .A1(G92), .A2(n650), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G79), .A2(n651), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G66), .A2(n646), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G54), .A2(n645), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(n584), .B(KEYINPUT15), .Z(n896) );
  INV_X1 U649 ( .A(n896), .ZN(n1002) );
  NAND2_X1 U650 ( .A1(n666), .A2(n1002), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G65), .A2(n646), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G53), .A2(n645), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G91), .A2(n650), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G78), .A2(n651), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n724) );
  INV_X1 U659 ( .A(n724), .ZN(G299) );
  XOR2_X1 U660 ( .A(KEYINPUT77), .B(n666), .Z(n593) );
  NOR2_X1 U661 ( .A1(G286), .A2(n593), .ZN(n595) );
  NOR2_X1 U662 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U664 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n597), .A2(n896), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U667 ( .A1(n1002), .A2(n666), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT78), .B(n599), .Z(n600) );
  NOR2_X1 U669 ( .A1(G559), .A2(n600), .ZN(n602) );
  NOR2_X1 U670 ( .A1(G868), .A2(n900), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G135), .A2(n985), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G111), .A2(n981), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n987), .A2(G99), .ZN(n605) );
  XOR2_X1 U676 ( .A(KEYINPUT80), .B(n605), .Z(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT79), .B(KEYINPUT18), .Z(n609) );
  NAND2_X1 U679 ( .A1(G123), .A2(n982), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n612), .B(KEYINPUT81), .ZN(n996) );
  XOR2_X1 U683 ( .A(G2096), .B(n996), .Z(n613) );
  NOR2_X1 U684 ( .A1(G2100), .A2(n613), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT82), .B(n614), .Z(G156) );
  NAND2_X1 U686 ( .A1(n896), .A2(G559), .ZN(n662) );
  XNOR2_X1 U687 ( .A(n900), .B(n662), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n615), .A2(G860), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G67), .A2(n646), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G55), .A2(n645), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G93), .A2(n650), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G80), .A2(n651), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n665) );
  XOR2_X1 U696 ( .A(n622), .B(n665), .Z(G145) );
  NAND2_X1 U697 ( .A1(G87), .A2(n623), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n646), .A2(n626), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G49), .A2(n645), .ZN(n627) );
  XOR2_X1 U702 ( .A(KEYINPUT83), .B(n627), .Z(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U704 ( .A(KEYINPUT84), .B(n630), .ZN(G288) );
  NAND2_X1 U705 ( .A1(G88), .A2(n650), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G75), .A2(n651), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G62), .A2(n646), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G50), .A2(n645), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G73), .A2(n651), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n637), .Z(n642) );
  NAND2_X1 U714 ( .A1(G61), .A2(n646), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G86), .A2(n650), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U717 ( .A(KEYINPUT85), .B(n640), .Z(n641) );
  NOR2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(G48), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U721 ( .A1(n645), .A2(G47), .ZN(n648) );
  NAND2_X1 U722 ( .A1(n646), .A2(G60), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U724 ( .A(KEYINPUT68), .B(n649), .Z(n655) );
  NAND2_X1 U725 ( .A1(G85), .A2(n650), .ZN(n653) );
  NAND2_X1 U726 ( .A1(G72), .A2(n651), .ZN(n652) );
  AND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(G290) );
  XOR2_X1 U729 ( .A(KEYINPUT19), .B(G166), .Z(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(G305), .ZN(n657) );
  XOR2_X1 U731 ( .A(n665), .B(n657), .Z(n659) );
  XOR2_X1 U732 ( .A(n900), .B(G299), .Z(n658) );
  XNOR2_X1 U733 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U734 ( .A(G288), .B(n660), .Z(n661) );
  XNOR2_X1 U735 ( .A(n661), .B(G290), .ZN(n1001) );
  XNOR2_X1 U736 ( .A(n1001), .B(n662), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n663), .A2(G868), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n664), .B(KEYINPUT86), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U747 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n674) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U750 ( .A1(n675), .A2(G218), .ZN(n676) );
  NAND2_X1 U751 ( .A1(G96), .A2(n676), .ZN(n948) );
  NAND2_X1 U752 ( .A1(G2106), .A2(n948), .ZN(n680) );
  NAND2_X1 U753 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U754 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G108), .A2(n678), .ZN(n949) );
  NAND2_X1 U756 ( .A1(G567), .A2(n949), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n680), .A2(n679), .ZN(n950) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U759 ( .A1(n950), .A2(n681), .ZN(n826) );
  NAND2_X1 U760 ( .A1(n826), .A2(G36), .ZN(G176) );
  INV_X1 U761 ( .A(G166), .ZN(G303) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n682) );
  NOR2_X1 U764 ( .A1(n683), .A2(n682), .ZN(n818) );
  NAND2_X1 U765 ( .A1(G140), .A2(n985), .ZN(n685) );
  NAND2_X1 U766 ( .A1(G104), .A2(n987), .ZN(n684) );
  NAND2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U768 ( .A(KEYINPUT34), .B(n686), .ZN(n692) );
  NAND2_X1 U769 ( .A1(n982), .A2(G128), .ZN(n687) );
  XNOR2_X1 U770 ( .A(n687), .B(KEYINPUT88), .ZN(n689) );
  NAND2_X1 U771 ( .A1(G116), .A2(n981), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U773 ( .A(n690), .B(KEYINPUT35), .Z(n691) );
  NOR2_X1 U774 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U775 ( .A(KEYINPUT36), .B(n693), .Z(n694) );
  XNOR2_X1 U776 ( .A(KEYINPUT89), .B(n694), .ZN(n998) );
  XNOR2_X1 U777 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NOR2_X1 U778 ( .A1(n998), .A2(n816), .ZN(n842) );
  NAND2_X1 U779 ( .A1(n818), .A2(n842), .ZN(n813) );
  NAND2_X1 U780 ( .A1(G131), .A2(n985), .ZN(n696) );
  NAND2_X1 U781 ( .A1(G95), .A2(n987), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n700) );
  NAND2_X1 U783 ( .A1(G107), .A2(n981), .ZN(n698) );
  NAND2_X1 U784 ( .A1(G119), .A2(n982), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n698), .A2(n697), .ZN(n699) );
  OR2_X1 U786 ( .A1(n700), .A2(n699), .ZN(n976) );
  AND2_X1 U787 ( .A1(n976), .A2(G1991), .ZN(n709) );
  INV_X1 U788 ( .A(G1996), .ZN(n954) );
  NAND2_X1 U789 ( .A1(G105), .A2(n987), .ZN(n701) );
  XNOR2_X1 U790 ( .A(n701), .B(KEYINPUT38), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n985), .A2(G141), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U793 ( .A1(G117), .A2(n981), .ZN(n705) );
  NAND2_X1 U794 ( .A1(G129), .A2(n982), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n978) );
  NOR2_X1 U797 ( .A1(n954), .A2(n978), .ZN(n708) );
  NOR2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n836) );
  INV_X1 U799 ( .A(n836), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n710), .A2(n818), .ZN(n806) );
  NAND2_X1 U801 ( .A1(n813), .A2(n806), .ZN(n803) );
  INV_X1 U802 ( .A(G40), .ZN(n711) );
  OR2_X1 U803 ( .A1(G1384), .A2(n711), .ZN(n712) );
  NOR2_X1 U804 ( .A1(G164), .A2(n712), .ZN(n713) );
  BUF_X1 U805 ( .A(n725), .Z(n763) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n763), .ZN(n745) );
  NAND2_X1 U807 ( .A1(G8), .A2(n745), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n725), .A2(G8), .ZN(n797) );
  NOR2_X1 U809 ( .A1(G1966), .A2(n797), .ZN(n715) );
  XNOR2_X1 U810 ( .A(n715), .B(n714), .ZN(n758) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n876) );
  NOR2_X1 U812 ( .A1(n763), .A2(n876), .ZN(n717) );
  AND2_X1 U813 ( .A1(n763), .A2(G1961), .ZN(n716) );
  NOR2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n749) );
  NAND2_X1 U815 ( .A1(n749), .A2(G171), .ZN(n744) );
  INV_X1 U816 ( .A(n725), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n730), .A2(G2072), .ZN(n718) );
  XNOR2_X1 U818 ( .A(KEYINPUT27), .B(n718), .ZN(n721) );
  NAND2_X1 U819 ( .A1(G1956), .A2(n725), .ZN(n719) );
  XOR2_X1 U820 ( .A(KEYINPUT92), .B(n719), .Z(n720) );
  NOR2_X1 U821 ( .A1(n721), .A2(n720), .ZN(n723) );
  NOR2_X1 U822 ( .A1(n724), .A2(n723), .ZN(n722) );
  XOR2_X1 U823 ( .A(n722), .B(KEYINPUT28), .Z(n741) );
  NAND2_X1 U824 ( .A1(n724), .A2(n723), .ZN(n739) );
  NOR2_X1 U825 ( .A1(n725), .A2(n954), .ZN(n726) );
  XOR2_X1 U826 ( .A(n726), .B(KEYINPUT26), .Z(n728) );
  NAND2_X1 U827 ( .A1(n763), .A2(G1341), .ZN(n727) );
  NAND2_X1 U828 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U829 ( .A1(n900), .A2(n729), .ZN(n734) );
  NAND2_X1 U830 ( .A1(G1348), .A2(n763), .ZN(n732) );
  NAND2_X1 U831 ( .A1(G2067), .A2(n730), .ZN(n731) );
  NAND2_X1 U832 ( .A1(n732), .A2(n731), .ZN(n735) );
  NOR2_X1 U833 ( .A1(n1002), .A2(n735), .ZN(n733) );
  OR2_X1 U834 ( .A1(n734), .A2(n733), .ZN(n737) );
  NAND2_X1 U835 ( .A1(n1002), .A2(n735), .ZN(n736) );
  NAND2_X1 U836 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U837 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U838 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U839 ( .A(KEYINPUT29), .B(n742), .Z(n743) );
  NAND2_X1 U840 ( .A1(n744), .A2(n743), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n758), .A2(n745), .ZN(n746) );
  NAND2_X1 U842 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U843 ( .A(n747), .B(KEYINPUT30), .ZN(n748) );
  NOR2_X1 U844 ( .A1(n748), .A2(G168), .ZN(n752) );
  OR2_X1 U845 ( .A1(G171), .A2(n749), .ZN(n750) );
  XNOR2_X1 U846 ( .A(n750), .B(KEYINPUT93), .ZN(n751) );
  XOR2_X1 U847 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n753) );
  XNOR2_X1 U848 ( .A(n754), .B(n753), .ZN(n755) );
  NAND2_X1 U849 ( .A1(n756), .A2(n755), .ZN(n762) );
  XNOR2_X1 U850 ( .A(KEYINPUT95), .B(n762), .ZN(n757) );
  NOR2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n774) );
  AND2_X1 U853 ( .A1(G286), .A2(G8), .ZN(n761) );
  NAND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n771) );
  INV_X1 U855 ( .A(G8), .ZN(n769) );
  NOR2_X1 U856 ( .A1(G1971), .A2(n797), .ZN(n765) );
  NOR2_X1 U857 ( .A1(G2090), .A2(n763), .ZN(n764) );
  NOR2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U859 ( .A1(n766), .A2(G303), .ZN(n767) );
  XNOR2_X1 U860 ( .A(n767), .B(KEYINPUT96), .ZN(n768) );
  OR2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U862 ( .A(n772), .B(KEYINPUT32), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n792) );
  NOR2_X1 U864 ( .A1(G1971), .A2(G303), .ZN(n775) );
  NOR2_X1 U865 ( .A1(G288), .A2(G1976), .ZN(n907) );
  NOR2_X1 U866 ( .A1(n775), .A2(n907), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n792), .A2(n776), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G288), .A2(G1976), .ZN(n910) );
  NAND2_X1 U869 ( .A1(n777), .A2(n910), .ZN(n778) );
  NOR2_X1 U870 ( .A1(n778), .A2(n797), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n780), .B(n779), .ZN(n781) );
  INV_X1 U872 ( .A(KEYINPUT33), .ZN(n784) );
  AND2_X1 U873 ( .A1(n781), .A2(n784), .ZN(n789) );
  INV_X1 U874 ( .A(n797), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n782), .A2(n907), .ZN(n783) );
  NOR2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(KEYINPUT97), .ZN(n787) );
  XNOR2_X1 U878 ( .A(G1981), .B(G305), .ZN(n894) );
  INV_X1 U879 ( .A(n894), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U881 ( .A1(G2090), .A2(G303), .ZN(n790) );
  NAND2_X1 U882 ( .A1(G8), .A2(n790), .ZN(n791) );
  XNOR2_X1 U883 ( .A(n791), .B(KEYINPUT98), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n794), .A2(n797), .ZN(n799) );
  NOR2_X1 U886 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U887 ( .A(n795), .B(KEYINPUT90), .Z(n796) );
  XNOR2_X1 U888 ( .A(KEYINPUT24), .B(n796), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n521), .A2(n800), .ZN(n801) );
  XNOR2_X1 U890 ( .A(KEYINPUT99), .B(n801), .ZN(n802) );
  NOR2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n805) );
  XNOR2_X1 U892 ( .A(G1986), .B(G290), .ZN(n904) );
  NAND2_X1 U893 ( .A1(n904), .A2(n818), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n821) );
  INV_X1 U895 ( .A(n806), .ZN(n809) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n976), .ZN(n843) );
  NOR2_X1 U898 ( .A1(n807), .A2(n843), .ZN(n808) );
  NOR2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n811) );
  AND2_X1 U900 ( .A1(n978), .A2(n954), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n810), .B(KEYINPUT100), .ZN(n839) );
  NOR2_X1 U902 ( .A1(n811), .A2(n839), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U905 ( .A(KEYINPUT101), .B(n815), .Z(n817) );
  NAND2_X1 U906 ( .A1(n998), .A2(n816), .ZN(n864) );
  NAND2_X1 U907 ( .A1(n817), .A2(n864), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n822), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n823), .ZN(G217) );
  INV_X1 U912 ( .A(n823), .ZN(G223) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n825) );
  XNOR2_X1 U916 ( .A(KEYINPUT106), .B(n825), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(G188) );
  NAND2_X1 U919 ( .A1(n985), .A2(G136), .ZN(n834) );
  NAND2_X1 U920 ( .A1(G100), .A2(n987), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G112), .A2(n981), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n982), .A2(G124), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT44), .B(n830), .Z(n831) );
  NOR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT112), .B(n835), .Z(G162) );
  XNOR2_X1 U928 ( .A(G160), .B(G2084), .ZN(n837) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(n848) );
  XOR2_X1 U930 ( .A(G2090), .B(G162), .Z(n838) );
  NOR2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U932 ( .A(n840), .B(KEYINPUT51), .ZN(n841) );
  NOR2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n846) );
  NOR2_X1 U934 ( .A1(n843), .A2(n996), .ZN(n844) );
  XOR2_X1 U935 ( .A(KEYINPUT117), .B(n844), .Z(n845) );
  NAND2_X1 U936 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U937 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U938 ( .A(KEYINPUT118), .B(n849), .Z(n862) );
  NAND2_X1 U939 ( .A1(G115), .A2(n981), .ZN(n851) );
  NAND2_X1 U940 ( .A1(G127), .A2(n982), .ZN(n850) );
  NAND2_X1 U941 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U942 ( .A(n852), .B(KEYINPUT47), .ZN(n854) );
  NAND2_X1 U943 ( .A1(G103), .A2(n987), .ZN(n853) );
  NAND2_X1 U944 ( .A1(n854), .A2(n853), .ZN(n857) );
  NAND2_X1 U945 ( .A1(n985), .A2(G139), .ZN(n855) );
  XOR2_X1 U946 ( .A(KEYINPUT114), .B(n855), .Z(n856) );
  NOR2_X1 U947 ( .A1(n857), .A2(n856), .ZN(n973) );
  XOR2_X1 U948 ( .A(G2072), .B(n973), .Z(n859) );
  XOR2_X1 U949 ( .A(G164), .B(G2078), .Z(n858) );
  NOR2_X1 U950 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U951 ( .A(KEYINPUT50), .B(n860), .Z(n861) );
  NOR2_X1 U952 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U953 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U954 ( .A(n865), .B(KEYINPUT119), .ZN(n866) );
  XNOR2_X1 U955 ( .A(KEYINPUT52), .B(n866), .ZN(n867) );
  XOR2_X1 U956 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n889) );
  NAND2_X1 U957 ( .A1(n867), .A2(n889), .ZN(n868) );
  NAND2_X1 U958 ( .A1(n868), .A2(G29), .ZN(n869) );
  XOR2_X1 U959 ( .A(KEYINPUT121), .B(n869), .Z(n946) );
  XOR2_X1 U960 ( .A(G25), .B(G1991), .Z(n875) );
  XOR2_X1 U961 ( .A(G2067), .B(G26), .Z(n870) );
  NAND2_X1 U962 ( .A1(n870), .A2(G28), .ZN(n873) );
  XNOR2_X1 U963 ( .A(KEYINPUT122), .B(G2072), .ZN(n871) );
  XNOR2_X1 U964 ( .A(G33), .B(n871), .ZN(n872) );
  NOR2_X1 U965 ( .A1(n873), .A2(n872), .ZN(n874) );
  NAND2_X1 U966 ( .A1(n875), .A2(n874), .ZN(n881) );
  XOR2_X1 U967 ( .A(n876), .B(G27), .Z(n878) );
  XNOR2_X1 U968 ( .A(G1996), .B(G32), .ZN(n877) );
  NOR2_X1 U969 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U970 ( .A(n879), .B(KEYINPUT123), .ZN(n880) );
  NOR2_X1 U971 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U972 ( .A(KEYINPUT53), .B(n882), .Z(n885) );
  XOR2_X1 U973 ( .A(KEYINPUT54), .B(G34), .Z(n883) );
  XNOR2_X1 U974 ( .A(G2084), .B(n883), .ZN(n884) );
  NAND2_X1 U975 ( .A1(n885), .A2(n884), .ZN(n887) );
  XNOR2_X1 U976 ( .A(G35), .B(G2090), .ZN(n886) );
  NOR2_X1 U977 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U978 ( .A(n889), .B(n888), .Z(n891) );
  INV_X1 U979 ( .A(G29), .ZN(n890) );
  NAND2_X1 U980 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U981 ( .A1(n892), .A2(G11), .ZN(n944) );
  INV_X1 U982 ( .A(G16), .ZN(n940) );
  XOR2_X1 U983 ( .A(n940), .B(KEYINPUT56), .Z(n918) );
  XOR2_X1 U984 ( .A(G168), .B(G1966), .Z(n893) );
  NOR2_X1 U985 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U986 ( .A(KEYINPUT57), .B(n895), .Z(n916) );
  XOR2_X1 U987 ( .A(G171), .B(G1961), .Z(n898) );
  XOR2_X1 U988 ( .A(n896), .B(G1348), .Z(n897) );
  NOR2_X1 U989 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U990 ( .A(KEYINPUT124), .B(n899), .ZN(n906) );
  XOR2_X1 U991 ( .A(n900), .B(G1341), .Z(n902) );
  XOR2_X1 U992 ( .A(G299), .B(G1956), .Z(n901) );
  NAND2_X1 U993 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U994 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U995 ( .A1(n906), .A2(n905), .ZN(n914) );
  XOR2_X1 U996 ( .A(n907), .B(KEYINPUT125), .Z(n909) );
  XNOR2_X1 U997 ( .A(G303), .B(G1971), .ZN(n908) );
  NOR2_X1 U998 ( .A1(n909), .A2(n908), .ZN(n911) );
  NAND2_X1 U999 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1000 ( .A(KEYINPUT126), .B(n912), .ZN(n913) );
  NOR2_X1 U1001 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1002 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1003 ( .A1(n918), .A2(n917), .ZN(n942) );
  XOR2_X1 U1004 ( .A(G5), .B(G1961), .Z(n935) );
  XOR2_X1 U1005 ( .A(G1348), .B(KEYINPUT59), .Z(n919) );
  XNOR2_X1 U1006 ( .A(G4), .B(n919), .ZN(n921) );
  XNOR2_X1 U1007 ( .A(G20), .B(G1956), .ZN(n920) );
  NOR2_X1 U1008 ( .A1(n921), .A2(n920), .ZN(n925) );
  XNOR2_X1 U1009 ( .A(G1341), .B(G19), .ZN(n923) );
  XNOR2_X1 U1010 ( .A(G1981), .B(G6), .ZN(n922) );
  NOR2_X1 U1011 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1012 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1013 ( .A(n926), .B(KEYINPUT60), .ZN(n933) );
  XNOR2_X1 U1014 ( .A(G1971), .B(G22), .ZN(n928) );
  XNOR2_X1 U1015 ( .A(G23), .B(G1976), .ZN(n927) );
  NOR2_X1 U1016 ( .A1(n928), .A2(n927), .ZN(n930) );
  XOR2_X1 U1017 ( .A(G1986), .B(G24), .Z(n929) );
  NAND2_X1 U1018 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1019 ( .A(KEYINPUT58), .B(n931), .ZN(n932) );
  NOR2_X1 U1020 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1021 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1022 ( .A(G21), .B(G1966), .ZN(n936) );
  NOR2_X1 U1023 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1024 ( .A(KEYINPUT61), .B(n938), .ZN(n939) );
  NAND2_X1 U1025 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1026 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1027 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1028 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1029 ( .A(KEYINPUT62), .B(n947), .Z(G311) );
  XNOR2_X1 U1030 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1031 ( .A(G132), .ZN(G219) );
  INV_X1 U1032 ( .A(G120), .ZN(G236) );
  INV_X1 U1033 ( .A(G96), .ZN(G221) );
  INV_X1 U1034 ( .A(G82), .ZN(G220) );
  INV_X1 U1035 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1036 ( .A1(n949), .A2(n948), .ZN(G325) );
  INV_X1 U1037 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1038 ( .A(KEYINPUT107), .B(n950), .ZN(G319) );
  XOR2_X1 U1039 ( .A(KEYINPUT41), .B(G2474), .Z(n952) );
  XNOR2_X1 U1040 ( .A(G1956), .B(G1976), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(n952), .B(n951), .ZN(n953) );
  XOR2_X1 U1042 ( .A(n953), .B(G1971), .Z(n956) );
  XOR2_X1 U1043 ( .A(n954), .B(G1961), .Z(n955) );
  XNOR2_X1 U1044 ( .A(n956), .B(n955), .ZN(n960) );
  XOR2_X1 U1045 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n958) );
  XNOR2_X1 U1046 ( .A(G1986), .B(G1966), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(n958), .B(n957), .ZN(n959) );
  XOR2_X1 U1048 ( .A(n960), .B(n959), .Z(n962) );
  XNOR2_X1 U1049 ( .A(G1991), .B(G1981), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(n962), .B(n961), .ZN(G229) );
  XOR2_X1 U1051 ( .A(KEYINPUT43), .B(G2678), .Z(n964) );
  XNOR2_X1 U1052 ( .A(G2072), .B(G2090), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(n964), .B(n963), .ZN(n968) );
  XOR2_X1 U1054 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n966) );
  XNOR2_X1 U1055 ( .A(G2067), .B(KEYINPUT42), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n966), .B(n965), .ZN(n967) );
  XOR2_X1 U1057 ( .A(n968), .B(n967), .Z(n970) );
  XNOR2_X1 U1058 ( .A(G2096), .B(G2100), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(n970), .B(n969), .ZN(n972) );
  XOR2_X1 U1060 ( .A(G2084), .B(G2078), .Z(n971) );
  XNOR2_X1 U1061 ( .A(n972), .B(n971), .ZN(G227) );
  XOR2_X1 U1062 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n975) );
  XNOR2_X1 U1063 ( .A(G164), .B(n973), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n975), .B(n974), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(n977), .B(n976), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(G160), .B(n978), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(n980), .B(n979), .ZN(n994) );
  NAND2_X1 U1068 ( .A1(G118), .A2(n981), .ZN(n984) );
  NAND2_X1 U1069 ( .A1(G130), .A2(n982), .ZN(n983) );
  NAND2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n992) );
  NAND2_X1 U1071 ( .A1(n985), .A2(G142), .ZN(n986) );
  XOR2_X1 U1072 ( .A(KEYINPUT113), .B(n986), .Z(n989) );
  NAND2_X1 U1073 ( .A1(n987), .A2(G106), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1075 ( .A(n990), .B(KEYINPUT45), .Z(n991) );
  NOR2_X1 U1076 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1077 ( .A(n994), .B(n993), .Z(n995) );
  XOR2_X1 U1078 ( .A(n996), .B(n995), .Z(n997) );
  XNOR2_X1 U1079 ( .A(G162), .B(n997), .ZN(n999) );
  XNOR2_X1 U1080 ( .A(n999), .B(n998), .ZN(n1000) );
  NOR2_X1 U1081 ( .A1(G37), .A2(n1000), .ZN(G395) );
  XOR2_X1 U1082 ( .A(KEYINPUT115), .B(n1001), .Z(n1004) );
  XOR2_X1 U1083 ( .A(n1002), .B(G286), .Z(n1003) );
  XNOR2_X1 U1084 ( .A(n1004), .B(n1003), .ZN(n1005) );
  XOR2_X1 U1085 ( .A(n1005), .B(G171), .Z(n1006) );
  NOR2_X1 U1086 ( .A1(n1006), .A2(G37), .ZN(n1007) );
  XNOR2_X1 U1087 ( .A(n1007), .B(KEYINPUT116), .ZN(G397) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT103), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(n1008), .B(G2454), .ZN(n1018) );
  XOR2_X1 U1090 ( .A(KEYINPUT104), .B(G2446), .Z(n1010) );
  XNOR2_X1 U1091 ( .A(G2451), .B(G2430), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(n1010), .B(n1009), .ZN(n1014) );
  XOR2_X1 U1093 ( .A(KEYINPUT102), .B(G2438), .Z(n1012) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G2435), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(n1014), .B(n1013), .Z(n1016) );
  XNOR2_X1 U1097 ( .A(G2443), .B(G2427), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NAND2_X1 U1100 ( .A1(n1019), .A2(G14), .ZN(n1020) );
  XOR2_X1 U1101 ( .A(n1020), .B(KEYINPUT105), .Z(n1026) );
  NAND2_X1 U1102 ( .A1(G319), .A2(n1026), .ZN(n1023) );
  NOR2_X1 U1103 ( .A1(G229), .A2(G227), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(KEYINPUT49), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1105 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  NOR2_X1 U1106 ( .A1(G395), .A2(G397), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(G225) );
  INV_X1 U1108 ( .A(G225), .ZN(G308) );
  INV_X1 U1109 ( .A(n1026), .ZN(G401) );
  INV_X1 U1110 ( .A(G108), .ZN(G238) );
endmodule

