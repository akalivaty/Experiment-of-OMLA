//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n216), .A2(G1), .A3(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n213), .A2(G20), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n251), .A2(new_n253), .A3(G274), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G232), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G107), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n256), .A2(new_n258), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n218), .A2(new_n252), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n254), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n249), .A2(new_n250), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT68), .A2(G1), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n274), .A2(KEYINPUT69), .A3(new_n253), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT69), .B1(new_n274), .B2(new_n253), .ZN(new_n276));
  OAI21_X1  g0076(.A(G244), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G179), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G20), .A2(G77), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT15), .B(G87), .ZN(new_n282));
  INV_X1    g0082(.A(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n281), .B1(new_n282), .B2(new_n284), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n218), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(new_n207), .B2(new_n259), .ZN(new_n291));
  NAND4_X1  g0091(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n218), .B1(new_n291), .B2(new_n292), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT68), .A2(G1), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT68), .A2(G1), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(G77), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n271), .A2(G13), .A3(G20), .A4(new_n273), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n221), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n295), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n268), .A2(new_n277), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n280), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n263), .A2(new_n221), .ZN(new_n310));
  MUX2_X1   g0110(.A(G222), .B(G223), .S(G1698), .Z(new_n311));
  OAI211_X1 g0111(.A(new_n267), .B(new_n310), .C1(new_n263), .C2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G274), .ZN(new_n313));
  AND2_X1   g0113(.A1(G1), .A2(G13), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n252), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n251), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G226), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n274), .A2(new_n253), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT69), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n274), .A2(KEYINPUT69), .A3(new_n253), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n307), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n296), .A2(new_n300), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G50), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n203), .A2(G20), .ZN(new_n329));
  INV_X1    g0129(.A(G150), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n329), .B1(new_n330), .B2(new_n286), .C1(new_n284), .C2(new_n287), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n294), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n328), .B(new_n332), .C1(G50), .C2(new_n302), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n324), .A2(new_n279), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n326), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n333), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(KEYINPUT9), .B1(new_n324), .B2(G190), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n325), .A2(G200), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT10), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT10), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n309), .B(new_n336), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT72), .ZN(new_n346));
  INV_X1    g0146(.A(G68), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G20), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n348), .B1(new_n284), .B2(new_n221), .C1(new_n286), .C2(new_n202), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n294), .A2(new_n349), .A3(KEYINPUT11), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT11), .B1(new_n294), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n352), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT72), .A3(new_n350), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n327), .A2(G68), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  INV_X1    g0160(.A(G238), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n321), .B2(new_n322), .ZN(new_n362));
  NOR2_X1   g0162(.A1(G226), .A2(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(G232), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(G1698), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n255), .B1(G33), .B2(G97), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n316), .B1(new_n366), .B2(new_n266), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n362), .A2(new_n367), .A3(KEYINPUT13), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  OAI21_X1  g0169(.A(G238), .B1(new_n275), .B2(new_n276), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G226), .B2(G1698), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n371), .B1(new_n373), .B2(new_n263), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n254), .B1(new_n267), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n369), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n360), .B(G169), .C1(new_n368), .C2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT13), .B1(new_n362), .B2(new_n367), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n370), .A2(new_n369), .A3(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(G179), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n360), .B1(new_n382), .B2(G169), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n359), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n368), .A2(new_n376), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G200), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n378), .B2(new_n379), .ZN(new_n388));
  OR3_X1    g0188(.A1(new_n386), .A2(new_n359), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n305), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(KEYINPUT71), .C1(new_n278), .C2(new_n387), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT71), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n387), .B1(new_n268), .B2(new_n277), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n305), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n306), .A2(new_n385), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n345), .A2(new_n384), .A3(new_n389), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G223), .A2(G1698), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n318), .B2(G1698), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n261), .B2(G33), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n259), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(new_n403), .A3(new_n404), .A4(new_n262), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n266), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n316), .B1(new_n319), .B2(new_n364), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n387), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n299), .A2(new_n272), .B1(new_n314), .B2(new_n252), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n254), .B1(new_n410), .B2(G232), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n403), .A2(new_n404), .A3(new_n262), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n318), .A2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G223), .B2(G1698), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n406), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n267), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(new_n416), .A3(new_n385), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n409), .A2(new_n417), .A3(KEYINPUT75), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n411), .A2(new_n416), .A3(new_n419), .A4(new_n385), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n418), .A2(KEYINPUT76), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT76), .B1(new_n418), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n287), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n302), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n327), .B2(new_n424), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT7), .B1(new_n263), .B2(new_n283), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT7), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n428), .B(G20), .C1(new_n260), .C2(new_n262), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G58), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n347), .ZN(new_n432));
  OAI21_X1  g0232(.A(G20), .B1(new_n432), .B2(new_n201), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n285), .A2(G159), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT16), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n296), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n404), .A2(new_n262), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT73), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n428), .B(new_n283), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G68), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n428), .B1(new_n412), .B2(new_n283), .ZN(new_n444));
  OAI211_X1 g0244(.A(KEYINPUT16), .B(new_n436), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT74), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n428), .B1(new_n255), .B2(G20), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n283), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n347), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n438), .B1(new_n449), .B2(new_n435), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT74), .A4(new_n294), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n426), .B1(new_n446), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n399), .B1(new_n423), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n418), .A2(new_n420), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT76), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n418), .A2(KEYINPUT76), .A3(new_n420), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n426), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n445), .A2(new_n294), .A3(new_n450), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT74), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n463), .B2(new_n451), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n459), .A2(KEYINPUT17), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n411), .A2(new_n416), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n279), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(G169), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT18), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT18), .ZN(new_n470));
  INV_X1    g0270(.A(new_n468), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n453), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n454), .A2(new_n465), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n398), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n271), .A2(G33), .A3(new_n273), .ZN(new_n475));
  AND4_X1   g0275(.A1(new_n289), .A2(new_n293), .A3(new_n302), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G116), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT79), .A2(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT79), .A2(G116), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n303), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n259), .A2(G97), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(G33), .B2(G283), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n480), .A2(G20), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n294), .A2(KEYINPUT20), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT20), .B1(new_n294), .B2(new_n484), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n477), .B(new_n481), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n271), .A2(G45), .A3(new_n273), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G41), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(G270), .B(new_n253), .C1(new_n488), .C2(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n315), .A2(new_n299), .A3(new_n494), .A4(G45), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n263), .A2(G303), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n224), .A2(G1698), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(G257), .B2(G1698), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n412), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n267), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n307), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT21), .B1(new_n487), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G257), .A2(G1698), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n224), .B2(G1698), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n403), .A3(new_n404), .A4(new_n262), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n266), .B1(new_n506), .B2(new_n497), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n493), .A2(new_n495), .ZN(new_n508));
  OAI211_X1 g0308(.A(KEYINPUT21), .B(G169), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n496), .A2(G179), .A3(new_n501), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n487), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(KEYINPUT82), .A3(new_n487), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n503), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n517), .A2(new_n518), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g0320(.A(G97), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(KEYINPUT6), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n283), .B1(new_n221), .B2(new_n286), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n223), .B1(new_n447), .B2(new_n448), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n294), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n302), .A2(G97), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n476), .B2(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n403), .A2(new_n404), .A3(new_n262), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n222), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT4), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n260), .A2(new_n262), .A3(G250), .A4(G1698), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT4), .A2(G244), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n260), .A2(new_n262), .A3(new_n535), .A4(new_n257), .ZN(new_n536));
  INV_X1    g0336(.A(G283), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n534), .B(new_n536), .C1(new_n259), .C2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n267), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n253), .C1(new_n488), .C2(new_n492), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n495), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT78), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT78), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n543), .A3(new_n495), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n530), .B1(G200), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n539), .A2(new_n542), .A3(G190), .A4(new_n544), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n545), .A2(new_n307), .B1(new_n527), .B2(new_n529), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n539), .A2(new_n542), .A3(new_n279), .A4(new_n544), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n488), .A2(G250), .A3(new_n253), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n315), .A2(G45), .A3(new_n299), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n222), .A2(G1698), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(G238), .B2(G1698), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n412), .A2(new_n555), .B1(new_n480), .B2(new_n259), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n553), .B1(new_n267), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT80), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n279), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n267), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n551), .A2(new_n552), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(new_n279), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT80), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n307), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n559), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n518), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n371), .A2(new_n283), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n284), .A2(KEYINPUT19), .A3(new_n521), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n403), .A2(new_n404), .A3(new_n283), .A4(new_n262), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n347), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n294), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n303), .A2(new_n282), .ZN(new_n576));
  INV_X1    g0376(.A(new_n282), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n296), .A2(new_n302), .A3(new_n475), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n574), .A2(new_n294), .B1(new_n303), .B2(new_n282), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n564), .A2(G200), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n560), .A2(new_n561), .A3(G190), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n476), .A2(G87), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n586), .A2(new_n581), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n566), .A2(new_n584), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n487), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n507), .A2(new_n508), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G190), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n592), .C1(new_n387), .C2(new_n591), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n516), .A2(new_n550), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n283), .B(G33), .C1(new_n478), .C2(new_n479), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT23), .B1(new_n283), .B2(G107), .ZN(new_n597));
  OR3_X1    g0397(.A1(new_n283), .A2(KEYINPUT23), .A3(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n568), .A2(G20), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT22), .B1(new_n255), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(KEYINPUT22), .A2(G87), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n573), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n595), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NOR4_X1   g0406(.A1(new_n604), .A2(new_n599), .A3(new_n601), .A4(KEYINPUT24), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n294), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n223), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT25), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n302), .B2(G107), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n476), .A2(G107), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(G250), .A2(G1698), .ZN(new_n615));
  INV_X1    g0415(.A(G257), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(G1698), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n403), .A3(new_n404), .A4(new_n262), .ZN(new_n618));
  NAND2_X1  g0418(.A1(G33), .A2(G294), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n266), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(G264), .B(new_n253), .C1(new_n488), .C2(new_n492), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT83), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n616), .A2(G1698), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G250), .B2(G1698), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n619), .B1(new_n412), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n267), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT83), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n621), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n623), .A2(new_n495), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(KEYINPUT84), .A3(new_n387), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n621), .A3(new_n495), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(G190), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT84), .B1(new_n630), .B2(new_n387), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n614), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(G169), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n630), .B2(new_n279), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n613), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n594), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n474), .A2(new_n641), .ZN(G372));
  INV_X1    g0442(.A(KEYINPUT86), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n487), .A2(new_n502), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT21), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n487), .B2(new_n511), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT85), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n551), .A2(new_n552), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n551), .B2(new_n552), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n560), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n307), .B1(new_n557), .B2(new_n279), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(G200), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n584), .A2(new_n652), .B1(new_n588), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n647), .A2(new_n550), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n636), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n643), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n589), .A2(new_n549), .A3(new_n548), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n545), .A2(new_n307), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n549), .A3(new_n530), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT87), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n548), .A2(new_n663), .A3(new_n549), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n662), .A2(new_n654), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n659), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n584), .A2(new_n652), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n588), .A2(new_n653), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n545), .A2(G200), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n527), .A3(new_n529), .A4(new_n547), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n661), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(KEYINPUT86), .A3(new_n636), .A4(new_n647), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n657), .A2(new_n666), .A3(new_n667), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n474), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n423), .A2(new_n453), .A3(new_n399), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT17), .B1(new_n459), .B2(new_n464), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n280), .A2(new_n305), .A3(new_n308), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n384), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n389), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n472), .A2(new_n469), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n342), .A2(new_n344), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n336), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n676), .A2(new_n686), .ZN(G369));
  AND2_X1   g0487(.A1(new_n283), .A2(G13), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n299), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n487), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT89), .Z(new_n696));
  INV_X1    g0496(.A(KEYINPUT90), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n696), .A2(new_n697), .A3(new_n646), .ZN(new_n698));
  INV_X1    g0498(.A(new_n503), .ZN(new_n699));
  INV_X1    g0499(.A(new_n515), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT82), .B1(new_n511), .B2(new_n487), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n593), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n696), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n697), .B1(new_n696), .B2(new_n646), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n638), .A2(new_n613), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n630), .A2(new_n387), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT84), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n633), .A3(new_n631), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n707), .B1(new_n711), .B2(new_n614), .ZN(new_n712));
  INV_X1    g0512(.A(new_n694), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n614), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n694), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n706), .A2(new_n716), .A3(G330), .ZN(new_n717));
  INV_X1    g0517(.A(new_n516), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n718), .A3(new_n713), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n694), .B(KEYINPUT91), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n707), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n717), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n208), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n569), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT92), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(new_n730), .B1(new_n212), .B2(new_n727), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  NAND4_X1  g0533(.A1(new_n662), .A2(new_n654), .A3(KEYINPUT26), .A4(new_n664), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n588), .A2(new_n585), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n580), .A2(new_n583), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n559), .A2(new_n563), .A3(new_n565), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n661), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n734), .B1(new_n739), .B2(new_n658), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n516), .A2(new_n639), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n673), .A3(new_n636), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n742), .A3(new_n667), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n743), .A2(KEYINPUT94), .A3(new_n713), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT94), .B1(new_n743), .B2(new_n713), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT29), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n675), .A2(new_n721), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT29), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n507), .A2(new_n508), .A3(new_n279), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(new_n623), .A3(new_n629), .A4(new_n557), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n751), .B1(new_n753), .B2(new_n545), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n591), .A2(G179), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n630), .A2(new_n545), .A3(new_n755), .A4(new_n651), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(KEYINPUT93), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n623), .A2(new_n629), .ZN(new_n759));
  INV_X1    g0559(.A(new_n545), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n510), .A2(new_n564), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(KEYINPUT30), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(new_n757), .B2(KEYINPUT93), .ZN(new_n763));
  OAI211_X1 g0563(.A(KEYINPUT31), .B(new_n720), .C1(new_n758), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n754), .A2(new_n762), .A3(new_n756), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n694), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT31), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n738), .A2(new_n672), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n712), .A2(new_n703), .A3(new_n769), .A4(new_n721), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n764), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n750), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n733), .B1(new_n773), .B2(G1), .ZN(G364));
  INV_X1    g0574(.A(new_n706), .ZN(new_n775));
  INV_X1    g0575(.A(G330), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n706), .A2(G330), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n270), .B1(new_n688), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n726), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n777), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n289), .B1(G20), .B2(new_n307), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n255), .A2(G355), .A3(new_n208), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G116), .B2(new_n208), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n531), .A2(new_n725), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n250), .B2(new_n213), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n247), .A2(G45), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n781), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n283), .A2(new_n279), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OR3_X1    g0602(.A1(new_n802), .A2(new_n387), .A3(KEYINPUT98), .ZN(new_n803));
  OAI21_X1  g0603(.A(KEYINPUT98), .B1(new_n802), .B2(new_n387), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n803), .A2(G190), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n803), .A2(new_n385), .A3(new_n804), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G50), .A2(new_n806), .B1(new_n808), .B2(G68), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n385), .A2(G179), .A3(G200), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n283), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n521), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n263), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n283), .A2(G179), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(G190), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n568), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n814), .A2(new_n385), .A3(G200), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(G107), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G190), .A2(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G159), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT32), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n809), .A2(new_n813), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n801), .A2(G190), .A3(new_n387), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT96), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n801), .A2(new_n820), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n827), .A2(G58), .B1(G77), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT97), .ZN(new_n830));
  INV_X1    g0630(.A(G326), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n805), .A2(new_n831), .B1(new_n832), .B2(new_n811), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT99), .ZN(new_n834));
  INV_X1    g0634(.A(new_n821), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G311), .A2(new_n828), .B1(new_n835), .B2(G329), .ZN(new_n836));
  INV_X1    g0636(.A(G322), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n836), .B(new_n263), .C1(new_n837), .C2(new_n826), .ZN(new_n838));
  INV_X1    g0638(.A(G303), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n537), .A2(new_n817), .B1(new_n815), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(KEYINPUT33), .B(G317), .Z(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n807), .B2(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n825), .A2(new_n830), .B1(new_n834), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n800), .B1(new_n844), .B2(new_n787), .ZN(new_n845));
  INV_X1    g0645(.A(new_n790), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n706), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n783), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NOR2_X1   g0649(.A1(new_n713), .A2(new_n390), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n309), .B1(new_n397), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n680), .A2(new_n694), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT101), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n853), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT101), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n393), .A2(new_n305), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n395), .B1(new_n857), .B2(KEYINPUT71), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n850), .B1(new_n858), .B2(new_n394), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n855), .B(new_n856), .C1(new_n859), .C2(new_n309), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n747), .ZN(new_n863));
  INV_X1    g0663(.A(new_n861), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n675), .A2(new_n721), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n781), .B1(new_n866), .B2(new_n772), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n772), .B2(new_n866), .ZN(new_n868));
  INV_X1    g0668(.A(new_n787), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n789), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n781), .B1(new_n870), .B2(G77), .ZN(new_n871));
  INV_X1    g0671(.A(new_n828), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n263), .B1(new_n832), .B2(new_n826), .C1(new_n872), .C2(new_n480), .ZN(new_n873));
  INV_X1    g0673(.A(new_n815), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n812), .B(new_n873), .C1(G107), .C2(new_n874), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n875), .B1(new_n537), .B2(new_n807), .C1(new_n839), .C2(new_n805), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n818), .A2(G87), .ZN(new_n877));
  INV_X1    g0677(.A(G311), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n821), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT100), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n827), .A2(G143), .B1(G159), .B2(new_n828), .ZN(new_n881));
  INV_X1    g0681(.A(G137), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n881), .B1(new_n882), .B2(new_n805), .C1(new_n330), .C2(new_n807), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT34), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n811), .A2(new_n431), .B1(new_n817), .B2(new_n347), .ZN(new_n886));
  INV_X1    g0686(.A(G132), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n531), .B1(new_n887), .B2(new_n821), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n886), .B(new_n888), .C1(G50), .C2(new_n874), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n883), .B2(new_n884), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n876), .A2(new_n880), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n871), .B1(new_n891), .B2(new_n787), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n864), .B2(new_n789), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n868), .A2(new_n893), .ZN(G384));
  INV_X1    g0694(.A(G116), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n289), .A2(new_n283), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT35), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n524), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n897), .B2(new_n524), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT36), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n212), .A2(new_n221), .A3(new_n432), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n202), .A2(G68), .ZN(new_n902));
  AOI211_X1 g0702(.A(G13), .B(new_n299), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(G169), .B1(new_n368), .B2(new_n376), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT14), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n380), .A3(new_n377), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n359), .A3(new_n713), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n436), .B1(new_n443), .B2(new_n444), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n438), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n445), .A2(new_n294), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n426), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n692), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n473), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n464), .B1(new_n422), .B2(new_n421), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n913), .B1(new_n471), .B2(new_n914), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT37), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT103), .B1(new_n453), .B2(new_n914), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n464), .A2(new_n923), .A3(new_n692), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n453), .A2(new_n471), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT37), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n918), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n921), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n917), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n917), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT39), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n918), .A2(new_n926), .A3(new_n927), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n453), .A2(KEYINPUT103), .A3(new_n914), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n923), .B1(new_n464), .B2(new_n692), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n679), .B2(new_n683), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n918), .A2(new_n926), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n937), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n938), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n917), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n932), .A2(new_n933), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n933), .B1(new_n932), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n909), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n865), .A2(new_n855), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n359), .A2(new_n694), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n384), .A2(new_n389), .A3(new_n951), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n386), .A2(new_n359), .A3(new_n388), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n359), .B(new_n694), .C1(new_n907), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n930), .A2(new_n931), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n956), .A2(new_n957), .B1(new_n683), .B2(new_n914), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n746), .A2(new_n474), .A3(new_n749), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n686), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n960), .B(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(new_n854), .A3(new_n860), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n641), .A2(new_n721), .B1(new_n767), .B2(new_n766), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT105), .B1(new_n766), .B2(new_n767), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT105), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n765), .A2(new_n967), .A3(KEYINPUT31), .A4(new_n694), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n964), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT40), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(new_n930), .C2(new_n931), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n952), .A2(new_n954), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(new_n861), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n770), .A3(new_n768), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n945), .B2(new_n943), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n972), .B1(new_n977), .B2(new_n971), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n474), .A2(new_n975), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n776), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n979), .B2(new_n978), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n963), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n299), .B2(new_n688), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n963), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n904), .B1(new_n983), .B2(new_n984), .ZN(G367));
  AOI22_X1  g0785(.A1(new_n239), .A2(new_n795), .B1(new_n725), .B2(new_n577), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n782), .B1(new_n791), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n713), .B1(new_n581), .B2(new_n587), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(new_n584), .A3(new_n652), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n669), .B2(new_n988), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n874), .A2(KEYINPUT46), .A3(G116), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT111), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n815), .A2(new_n480), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n991), .A2(new_n992), .B1(KEYINPUT46), .B2(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n872), .A2(new_n537), .B1(new_n223), .B2(new_n811), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n992), .B2(new_n991), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n832), .B2(new_n807), .C1(new_n878), .C2(new_n805), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n994), .B(new_n997), .C1(G303), .C2(new_n827), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n817), .A2(new_n521), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n531), .B(new_n999), .C1(G317), .C2(new_n835), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT112), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(G143), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n805), .A2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n255), .B1(new_n330), .B2(new_n826), .C1(new_n872), .C2(new_n202), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n811), .A2(new_n347), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n817), .A2(new_n221), .ZN(new_n1007));
  NOR4_X1   g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n815), .A2(new_n431), .B1(new_n821), .B2(new_n882), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT113), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1009), .A2(KEYINPUT113), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G159), .C2(new_n808), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n998), .A2(new_n1002), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT47), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n787), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1013), .A2(KEYINPUT47), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n987), .B1(new_n846), .B2(new_n990), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n779), .B(KEYINPUT110), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n717), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n720), .A2(new_n530), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n550), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n720), .A2(new_n549), .A3(new_n548), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n719), .A2(new_n722), .A3(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT107), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT107), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1025), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT44), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n723), .B2(new_n1023), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n719), .A2(new_n722), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1023), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(KEYINPUT44), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT45), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1019), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1035), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1037), .A2(new_n717), .A3(new_n1033), .A4(new_n1027), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n719), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT108), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n718), .A2(new_n713), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n714), .A2(new_n715), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1044), .A2(new_n1041), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1042), .B1(new_n1045), .B2(new_n1040), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n778), .A2(KEYINPUT109), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1042), .C1(new_n1045), .C2(new_n1040), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n773), .B1(new_n1039), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n726), .B(KEYINPUT41), .Z(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1018), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n717), .A2(KEYINPUT106), .A3(new_n1031), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT106), .B1(new_n717), .B2(new_n1031), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1040), .A2(new_n1023), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n661), .B1(new_n1021), .B2(new_n639), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1063), .A2(KEYINPUT42), .B1(new_n721), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(KEYINPUT42), .B2(new_n1063), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1062), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1060), .A2(new_n1067), .A3(new_n1066), .A4(new_n1061), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1017), .B1(new_n1055), .B2(new_n1071), .ZN(G387));
  AOI21_X1  g0872(.A(new_n796), .B1(new_n236), .B2(G45), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n728), .ZN(new_n1074));
  AOI211_X1 g0874(.A(G45), .B(new_n1074), .C1(G68), .C2(G77), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT115), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n287), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT50), .B1(new_n287), .B2(G50), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1073), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1074), .A2(new_n208), .A3(new_n255), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(G107), .B2(new_n208), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT114), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n792), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n827), .A2(G317), .B1(G303), .B2(new_n828), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n878), .B2(new_n807), .C1(new_n837), .C2(new_n805), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n811), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1092), .A2(G283), .B1(new_n874), .B2(G294), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT49), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n412), .B1(new_n821), .B2(new_n831), .C1(new_n480), .C2(new_n817), .ZN(new_n1098));
  OR3_X1    g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n807), .A2(new_n287), .B1(new_n347), .B2(new_n872), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT116), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n531), .B1(new_n330), .B2(new_n821), .C1(new_n202), .C2(new_n826), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n815), .A2(new_n221), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n811), .A2(new_n282), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n1102), .A2(new_n999), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n822), .B2(new_n805), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1099), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n782), .B(new_n1086), .C1(new_n1107), .C2(new_n787), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT117), .Z(new_n1109));
  NAND3_X1  g0909(.A1(new_n714), .A2(new_n715), .A3(new_n790), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1109), .A2(new_n1110), .B1(new_n1111), .B2(new_n1018), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n727), .B1(new_n1111), .B2(new_n773), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n773), .B2(new_n1111), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(G393));
  NAND3_X1  g0916(.A1(new_n1036), .A2(new_n1038), .A3(new_n1018), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n791), .B1(new_n521), .B2(new_n208), .C1(new_n244), .C2(new_n796), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n781), .B1(new_n1118), .B2(KEYINPUT118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n826), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n806), .A2(G317), .B1(G311), .B2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT52), .Z(new_n1122));
  OAI221_X1 g0922(.A(new_n263), .B1(new_n817), .B2(new_n223), .C1(new_n872), .C2(new_n832), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n874), .A2(G283), .B1(new_n835), .B2(G322), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT119), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n480), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1123), .B(new_n1126), .C1(new_n1127), .C2(new_n1092), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n808), .A2(G303), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1122), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n805), .A2(new_n330), .B1(new_n822), .B2(new_n826), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT51), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n877), .B1(new_n347), .B2(new_n815), .C1(new_n221), .C2(new_n811), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n872), .A2(new_n287), .B1(new_n821), .B2(new_n1003), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1133), .A2(new_n412), .A3(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n1135), .C1(new_n202), .C2(new_n807), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n869), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1119), .B(new_n1137), .C1(KEYINPUT118), .C2(new_n1118), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1023), .B2(new_n846), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1111), .A2(new_n773), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1039), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1111), .A2(new_n773), .A3(new_n1038), .A4(new_n1036), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n726), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1117), .B(new_n1139), .C1(new_n1142), .C2(new_n1144), .ZN(G390));
  AOI21_X1  g0945(.A(new_n776), .B1(new_n965), .B2(new_n969), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n474), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n961), .A2(new_n686), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n975), .A2(G330), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n973), .B1(new_n862), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n771), .A2(new_n955), .A3(G330), .A4(new_n864), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n864), .B1(new_n744), .B2(new_n745), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n855), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n771), .A2(G330), .A3(new_n864), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1155), .A2(new_n973), .B1(new_n1146), .B2(new_n974), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n950), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1152), .A2(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT38), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n925), .B2(new_n928), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n473), .A2(new_n925), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n927), .B1(new_n940), .B2(new_n937), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n930), .A2(new_n1164), .A3(KEYINPUT39), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n915), .B1(new_n679), .B2(new_n683), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n934), .A2(new_n937), .B1(KEYINPUT37), .B2(new_n920), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n944), .B1(new_n1168), .B2(new_n945), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT104), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n932), .A2(new_n946), .A3(new_n933), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n956), .A2(new_n908), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n909), .B1(new_n943), .B2(new_n945), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n743), .A2(new_n713), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT94), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n743), .A2(KEYINPUT94), .A3(new_n713), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n853), .B1(new_n1179), .B2(new_n864), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1174), .B1(new_n1180), .B2(new_n973), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1173), .A2(new_n1181), .A3(new_n1151), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1146), .A2(new_n974), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1173), .B2(new_n1181), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1159), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1173), .A2(new_n1181), .A3(new_n1151), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n961), .A2(new_n686), .A3(new_n1147), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1180), .A2(new_n1151), .A3(new_n1150), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1174), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1154), .B2(new_n955), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n947), .A2(new_n948), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1172), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1186), .B(new_n1190), .C1(new_n1194), .C2(new_n1183), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1185), .A2(new_n1195), .A3(new_n726), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n263), .B1(new_n821), .B2(new_n832), .C1(new_n872), .C2(new_n521), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n816), .B(new_n1197), .C1(G68), .C2(new_n818), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n811), .A2(new_n221), .B1(new_n826), .B2(new_n895), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT120), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT120), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G107), .A2(new_n808), .B1(new_n806), .B2(G283), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G128), .A2(new_n806), .B1(new_n808), .B2(G137), .ZN(new_n1204));
  INV_X1    g1004(.A(G125), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n826), .A2(new_n887), .B1(new_n821), .B2(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT54), .B(G143), .Z(new_n1207));
  AOI211_X1 g1007(.A(new_n263), .B(new_n1206), .C1(new_n828), .C2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1092), .A2(G159), .B1(new_n818), .B2(G50), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n815), .A2(new_n330), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT53), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1204), .A2(new_n1208), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1203), .A2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n781), .B1(new_n424), .B2(new_n870), .C1(new_n1213), .C2(new_n869), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1193), .B2(new_n788), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1018), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1196), .A2(new_n1217), .ZN(G378));
  INV_X1    g1018(.A(new_n1018), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n685), .A2(new_n335), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n337), .A2(new_n692), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n685), .B(new_n335), .C1(new_n337), .C2(new_n692), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n970), .B1(new_n930), .B2(new_n1164), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT40), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n776), .B(new_n1229), .C1(new_n1231), .C2(new_n972), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1229), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n978), .B2(G330), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n908), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1232), .A2(new_n1234), .B1(new_n1235), .B2(new_n958), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT40), .B1(new_n1168), .B2(new_n945), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1230), .A2(KEYINPUT40), .B1(new_n1237), .B2(new_n970), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1229), .B1(new_n1238), .B2(new_n776), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n978), .A2(G330), .A3(new_n1233), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(new_n949), .A3(new_n1240), .A4(new_n959), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1219), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n781), .B1(new_n870), .B2(G50), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n531), .A2(G41), .ZN(new_n1244));
  AOI211_X1 g1044(.A(G50), .B(new_n1244), .C1(new_n259), .C2(new_n249), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1120), .A2(G107), .B1(new_n828), .B2(new_n577), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n537), .B2(new_n821), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1247), .A2(new_n1006), .A3(new_n1103), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n817), .A2(new_n431), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT121), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n808), .B2(G97), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n806), .A2(G116), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1248), .A2(new_n1251), .A3(new_n1244), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT58), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1245), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n811), .A2(new_n330), .ZN(new_n1256));
  INV_X1    g1056(.A(G128), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n872), .A2(new_n882), .B1(new_n826), .B2(new_n1257), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1256), .B(new_n1258), .C1(new_n874), .C2(new_n1207), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n1205), .B2(new_n805), .C1(new_n887), .C2(new_n807), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT59), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n818), .A2(G159), .ZN(new_n1262));
  AOI211_X1 g1062(.A(G33), .B(G41), .C1(new_n835), .C2(G124), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1260), .A2(KEYINPUT59), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1255), .B1(new_n1254), .B2(new_n1253), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1243), .B1(new_n1266), .B2(new_n787), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1233), .B2(new_n789), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT122), .Z(new_n1269));
  NOR2_X1   g1069(.A1(new_n1242), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1182), .A2(new_n1184), .A3(new_n1159), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n1187), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT57), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1195), .A2(new_n1148), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n727), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1271), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(G375));
  INV_X1    g1081(.A(new_n1158), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1187), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1054), .A3(new_n1159), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n781), .B1(new_n870), .B2(G68), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n263), .B1(new_n821), .B2(new_n839), .C1(new_n872), .C2(new_n223), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1007), .B(new_n1286), .C1(G97), .C2(new_n874), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1104), .B1(G283), .B2(new_n1120), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1289), .A2(KEYINPUT123), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(KEYINPUT123), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(G294), .A2(new_n806), .B1(new_n808), .B2(new_n1127), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1287), .A2(new_n1290), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1250), .B1(new_n808), .B2(new_n1207), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n887), .B2(new_n805), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1092), .A2(G50), .B1(G150), .B2(new_n828), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1296), .B(KEYINPUT124), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n531), .B1(new_n1257), .B2(new_n821), .C1(new_n822), .C2(new_n815), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(G137), .B2(new_n827), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1295), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1285), .B1(new_n1301), .B2(new_n787), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n955), .B2(new_n789), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1284), .B(new_n1303), .C1(new_n1219), .C2(new_n1282), .ZN(G381));
  AND3_X1   g1104(.A1(new_n1112), .A2(new_n1114), .A3(new_n848), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1117), .A2(new_n1139), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1144), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(new_n1141), .ZN(new_n1308));
  INV_X1    g1108(.A(G384), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1305), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1310), .A2(G381), .ZN(new_n1311));
  OR4_X1    g1111(.A1(G387), .A2(G375), .A3(new_n1311), .A4(G378), .ZN(G407));
  INV_X1    g1112(.A(G378), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n693), .A2(G213), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1280), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(G407), .A2(G213), .A3(new_n1316), .ZN(G409));
  NOR2_X1   g1117(.A1(G387), .A2(new_n1308), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1053), .B1(new_n1143), .B2(new_n773), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1070), .B(new_n1069), .C1(new_n1319), .C2(new_n1018), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G390), .B1(new_n1320), .B2(new_n1017), .ZN(new_n1321));
  OAI21_X1  g1121(.A(KEYINPUT126), .B1(new_n1318), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n848), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1305), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT126), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G387), .A2(new_n1308), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1320), .A2(new_n1017), .A3(G390), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1324), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1325), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1278), .B1(new_n1273), .B2(new_n1187), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n726), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1272), .ZN(new_n1335));
  OAI211_X1 g1135(.A(G378), .B(new_n1270), .C1(new_n1334), .C2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1277), .A2(new_n1054), .A3(new_n1272), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1270), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1313), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1303), .B1(new_n1282), .B2(new_n1219), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1159), .A2(KEYINPUT60), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1283), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1188), .A2(new_n1187), .A3(new_n1189), .A4(KEYINPUT60), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n726), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1342), .B1(new_n1344), .B2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1348), .A2(G384), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1346), .B1(new_n1283), .B2(new_n1343), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1350), .A2(new_n1309), .A3(new_n1342), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1340), .A2(new_n1341), .A3(new_n1314), .A4(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1315), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1355));
  OAI211_X1 g1155(.A(G2897), .B(new_n1315), .C1(new_n1349), .C2(new_n1351), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1348), .A2(G384), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1309), .B1(new_n1350), .B2(new_n1342), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1315), .A2(G2897), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1357), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1356), .A2(new_n1360), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1353), .B(new_n1354), .C1(new_n1355), .C2(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1341), .B1(new_n1355), .B2(new_n1352), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1332), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1364));
  AND2_X1   g1164(.A1(new_n1356), .A2(new_n1360), .ZN(new_n1365));
  AOI21_X1  g1165(.A(G378), .B1(new_n1270), .B2(new_n1337), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1366), .B1(G378), .B2(new_n1280), .ZN(new_n1367));
  OAI211_X1 g1167(.A(KEYINPUT125), .B(new_n1365), .C1(new_n1367), .C2(new_n1315), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT125), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1369), .B1(new_n1355), .B2(new_n1361), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1368), .A2(new_n1370), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1325), .A2(new_n1354), .A3(new_n1331), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1340), .A2(new_n1314), .A3(new_n1352), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT63), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1372), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT127), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1376), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1355), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1352), .ZN(new_n1378));
  NAND4_X1  g1178(.A1(new_n1371), .A2(new_n1375), .A3(new_n1377), .A4(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1364), .A2(new_n1379), .ZN(G405));
  NOR2_X1   g1180(.A1(new_n1280), .A2(G378), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1381), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1332), .A2(new_n1336), .A3(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1336), .ZN(new_n1384));
  OAI211_X1 g1184(.A(new_n1325), .B(new_n1331), .C1(new_n1384), .C2(new_n1381), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1383), .A2(new_n1385), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1386), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1383), .A2(new_n1352), .A3(new_n1385), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1387), .A2(new_n1388), .ZN(G402));
endmodule


