

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744;

  BUF_X1 U365 ( .A(n682), .Z(n674) );
  XNOR2_X1 U366 ( .A(n573), .B(n572), .ZN(n658) );
  XNOR2_X1 U367 ( .A(n344), .B(n568), .ZN(n633) );
  OR2_X1 U368 ( .A1(n569), .A2(n394), .ZN(n393) );
  NAND2_X1 U369 ( .A1(n564), .A2(n565), .ZN(n344) );
  BUF_X2 U370 ( .A(n515), .Z(n610) );
  OR2_X1 U371 ( .A1(n662), .A2(G902), .ZN(n382) );
  XNOR2_X1 U372 ( .A(G113), .B(n343), .ZN(n475) );
  BUF_X1 U373 ( .A(G143), .Z(n343) );
  NOR2_X2 U374 ( .A1(G953), .A2(G237), .ZN(n469) );
  NAND2_X1 U375 ( .A1(n342), .A2(n576), .ZN(n577) );
  NAND2_X1 U376 ( .A1(n578), .A2(KEYINPUT44), .ZN(n342) );
  XNOR2_X2 U377 ( .A(G146), .B(G125), .ZN(n452) );
  NOR2_X1 U378 ( .A1(n608), .A2(n607), .ZN(n605) );
  XNOR2_X2 U379 ( .A(n481), .B(n480), .ZN(n509) );
  XNOR2_X2 U380 ( .A(n610), .B(n516), .ZN(n563) );
  XNOR2_X2 U381 ( .A(n457), .B(G134), .ZN(n367) );
  XNOR2_X1 U382 ( .A(n393), .B(KEYINPUT22), .ZN(n558) );
  NOR2_X1 U383 ( .A1(n621), .A2(n620), .ZN(n491) );
  XNOR2_X1 U384 ( .A(n404), .B(G953), .ZN(n733) );
  OR2_X1 U385 ( .A1(n512), .A2(n544), .ZN(n703) );
  OR2_X1 U386 ( .A1(n517), .A2(n559), .ZN(n498) );
  XNOR2_X1 U387 ( .A(n358), .B(n347), .ZN(n544) );
  BUF_X1 U388 ( .A(n604), .Z(n345) );
  INV_X1 U389 ( .A(KEYINPUT81), .ZN(n398) );
  AND2_X1 U390 ( .A1(n377), .A2(n374), .ZN(n373) );
  OR2_X1 U391 ( .A1(n378), .A2(n383), .ZN(n372) );
  AND2_X1 U392 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U393 ( .A(n546), .B(n547), .ZN(n360) );
  AND2_X1 U394 ( .A1(n521), .A2(n520), .ZN(n531) );
  XNOR2_X1 U395 ( .A(n548), .B(KEYINPUT102), .ZN(n504) );
  NAND2_X1 U396 ( .A1(n379), .A2(n505), .ZN(n709) );
  NOR2_X1 U397 ( .A1(n544), .A2(n543), .ZN(n357) );
  AND2_X1 U398 ( .A1(n604), .A2(n605), .ZN(n565) );
  NAND2_X1 U399 ( .A1(n524), .A2(n605), .ZN(n428) );
  XNOR2_X1 U400 ( .A(n397), .B(n396), .ZN(n446) );
  XNOR2_X1 U401 ( .A(n398), .B(G110), .ZN(n397) );
  XNOR2_X1 U402 ( .A(G104), .B(G107), .ZN(n396) );
  NOR2_X1 U403 ( .A1(n633), .A2(n569), .ZN(n380) );
  NOR2_X1 U404 ( .A1(n569), .A2(n353), .ZN(n546) );
  XNOR2_X1 U405 ( .A(n357), .B(n545), .ZN(n569) );
  XNOR2_X1 U406 ( .A(n524), .B(KEYINPUT1), .ZN(n604) );
  NOR2_X1 U407 ( .A1(n732), .A2(KEYINPUT75), .ZN(n585) );
  NAND2_X2 U408 ( .A1(n373), .A2(n372), .ZN(n732) );
  XNOR2_X2 U409 ( .A(n729), .B(n403), .ZN(n434) );
  XNOR2_X2 U410 ( .A(n367), .B(n401), .ZN(n729) );
  OR2_X1 U411 ( .A1(n694), .A2(n366), .ZN(n361) );
  INV_X1 U412 ( .A(n622), .ZN(n365) );
  NAND2_X1 U413 ( .A1(n362), .A2(n352), .ZN(n351) );
  INV_X1 U414 ( .A(n360), .ZN(n352) );
  INV_X1 U415 ( .A(n712), .ZN(n384) );
  INV_X1 U416 ( .A(KEYINPUT76), .ZN(n383) );
  NOR2_X1 U417 ( .A1(n384), .A2(n383), .ZN(n376) );
  INV_X1 U418 ( .A(n655), .ZN(n375) );
  AND2_X1 U419 ( .A1(n364), .A2(n363), .ZN(n576) );
  INV_X1 U420 ( .A(n691), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n402), .B(G101), .ZN(n451) );
  INV_X1 U422 ( .A(KEYINPUT66), .ZN(n402) );
  XNOR2_X1 U423 ( .A(KEYINPUT68), .B(G137), .ZN(n400) );
  INV_X1 U424 ( .A(KEYINPUT39), .ZN(n465) );
  NOR2_X1 U425 ( .A1(n391), .A2(n465), .ZN(n386) );
  XNOR2_X1 U426 ( .A(n440), .B(n439), .ZN(n447) );
  XNOR2_X1 U427 ( .A(G116), .B(G113), .ZN(n439) );
  XNOR2_X1 U428 ( .A(n438), .B(G119), .ZN(n440) );
  INV_X1 U429 ( .A(KEYINPUT3), .ZN(n438) );
  XNOR2_X1 U430 ( .A(n418), .B(n369), .ZN(n482) );
  INV_X1 U431 ( .A(KEYINPUT8), .ZN(n369) );
  XOR2_X1 U432 ( .A(KEYINPUT95), .B(G107), .Z(n485) );
  NAND2_X1 U433 ( .A1(n360), .A2(KEYINPUT91), .ZN(n359) );
  XNOR2_X1 U434 ( .A(n533), .B(n464), .ZN(n618) );
  NAND2_X1 U435 ( .A1(G234), .A2(G237), .ZN(n429) );
  XNOR2_X1 U436 ( .A(n452), .B(KEYINPUT10), .ZN(n468) );
  XOR2_X1 U437 ( .A(KEYINPUT12), .B(KEYINPUT94), .Z(n471) );
  XNOR2_X1 U438 ( .A(G122), .B(G104), .ZN(n473) );
  XNOR2_X1 U439 ( .A(n451), .B(n450), .ZN(n455) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n450) );
  INV_X1 U441 ( .A(G237), .ZN(n442) );
  NOR2_X1 U442 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n446), .B(n395), .ZN(n449) );
  INV_X1 U444 ( .A(KEYINPUT16), .ZN(n395) );
  XNOR2_X1 U445 ( .A(G140), .B(KEYINPUT86), .ZN(n412) );
  XNOR2_X1 U446 ( .A(G119), .B(G128), .ZN(n410) );
  XNOR2_X1 U447 ( .A(n709), .B(KEYINPUT96), .ZN(n536) );
  NAND2_X1 U448 ( .A1(n388), .A2(n385), .ZN(n537) );
  NAND2_X1 U449 ( .A1(n387), .A2(n386), .ZN(n385) );
  NAND2_X1 U450 ( .A1(n565), .A2(n610), .ZN(n353) );
  NAND2_X1 U451 ( .A1(n551), .A2(n492), .ZN(n394) );
  INV_X1 U452 ( .A(KEYINPUT64), .ZN(n404) );
  XNOR2_X1 U453 ( .A(n370), .B(n368), .ZN(n670) );
  AND2_X1 U454 ( .A1(n482), .A2(G217), .ZN(n368) );
  XNOR2_X1 U455 ( .A(n486), .B(n483), .ZN(n371) );
  OR2_X1 U456 ( .A1(n733), .A2(G952), .ZN(n687) );
  INV_X1 U457 ( .A(n706), .ZN(n356) );
  XOR2_X1 U458 ( .A(n441), .B(n447), .Z(n346) );
  XOR2_X1 U459 ( .A(n511), .B(KEYINPUT65), .Z(n347) );
  AND2_X1 U460 ( .A1(n361), .A2(n365), .ZN(n348) );
  AND2_X1 U461 ( .A1(n384), .A2(n383), .ZN(n349) );
  AND2_X1 U462 ( .A1(n351), .A2(n348), .ZN(n350) );
  INV_X1 U463 ( .A(KEYINPUT91), .ZN(n366) );
  NAND2_X1 U464 ( .A1(n350), .A2(n359), .ZN(n364) );
  AND2_X1 U465 ( .A1(n614), .A2(n353), .ZN(n615) );
  XNOR2_X2 U466 ( .A(n354), .B(n399), .ZN(n457) );
  XNOR2_X2 U467 ( .A(KEYINPUT72), .B(G143), .ZN(n354) );
  AND2_X1 U468 ( .A1(n360), .A2(n355), .ZN(n710) );
  INV_X1 U469 ( .A(n709), .ZN(n355) );
  AND2_X1 U470 ( .A1(n360), .A2(n356), .ZN(n708) );
  NAND2_X1 U471 ( .A1(n533), .A2(n617), .ZN(n358) );
  AND2_X1 U472 ( .A1(n694), .A2(n366), .ZN(n362) );
  XNOR2_X1 U473 ( .A(n367), .B(n371), .ZN(n370) );
  XNOR2_X1 U474 ( .A(n380), .B(KEYINPUT34), .ZN(n571) );
  NAND2_X1 U475 ( .A1(n378), .A2(n349), .ZN(n377) );
  XNOR2_X1 U476 ( .A(n529), .B(KEYINPUT48), .ZN(n378) );
  INV_X1 U477 ( .A(n505), .ZN(n508) );
  NAND2_X1 U478 ( .A1(n536), .A2(n706), .ZN(n510) );
  INV_X1 U479 ( .A(n509), .ZN(n379) );
  XNOR2_X2 U480 ( .A(n382), .B(G472), .ZN(n515) );
  XNOR2_X1 U481 ( .A(n434), .B(n346), .ZN(n662) );
  INV_X1 U482 ( .A(n504), .ZN(n387) );
  NAND2_X1 U483 ( .A1(n391), .A2(n465), .ZN(n389) );
  NAND2_X1 U484 ( .A1(n504), .A2(n465), .ZN(n390) );
  NAND2_X1 U485 ( .A1(n445), .A2(n493), .ZN(n503) );
  NAND2_X1 U486 ( .A1(n445), .A2(n392), .ZN(n391) );
  AND2_X1 U487 ( .A1(n618), .A2(n493), .ZN(n392) );
  AND2_X2 U488 ( .A1(n595), .A2(n594), .ZN(n682) );
  NAND2_X1 U489 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U491 ( .A(KEYINPUT60), .ZN(n601) );
  XNOR2_X1 U492 ( .A(n654), .B(n653), .ZN(G75) );
  INV_X1 U493 ( .A(G128), .ZN(n399) );
  XNOR2_X1 U494 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n453) );
  XNOR2_X1 U495 ( .A(n453), .B(n400), .ZN(n401) );
  XNOR2_X1 U496 ( .A(n451), .B(G146), .ZN(n403) );
  XOR2_X1 U497 ( .A(G131), .B(G140), .Z(n466) );
  XOR2_X1 U498 ( .A(n466), .B(n446), .Z(n406) );
  NAND2_X1 U499 ( .A1(G227), .A2(n733), .ZN(n405) );
  XNOR2_X1 U500 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n434), .B(n407), .ZN(n675) );
  OR2_X2 U502 ( .A1(n675), .A2(G902), .ZN(n408) );
  XNOR2_X2 U503 ( .A(n408), .B(G469), .ZN(n524) );
  XNOR2_X1 U504 ( .A(KEYINPUT85), .B(KEYINPUT24), .ZN(n409) );
  XNOR2_X1 U505 ( .A(n409), .B(n468), .ZN(n417) );
  XOR2_X1 U506 ( .A(G110), .B(G137), .Z(n411) );
  XNOR2_X1 U507 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U508 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n413) );
  XNOR2_X1 U509 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U510 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U511 ( .A(n417), .B(n416), .ZN(n420) );
  NAND2_X1 U512 ( .A1(n733), .A2(G234), .ZN(n418) );
  NAND2_X1 U513 ( .A1(n482), .A2(G221), .ZN(n419) );
  XNOR2_X1 U514 ( .A(n420), .B(n419), .ZN(n667) );
  NOR2_X1 U515 ( .A1(G902), .A2(n667), .ZN(n425) );
  XNOR2_X1 U516 ( .A(G902), .B(KEYINPUT15), .ZN(n589) );
  NAND2_X1 U517 ( .A1(n589), .A2(G234), .ZN(n421) );
  XNOR2_X1 U518 ( .A(n421), .B(KEYINPUT20), .ZN(n426) );
  NAND2_X1 U519 ( .A1(G217), .A2(n426), .ZN(n423) );
  INV_X1 U520 ( .A(KEYINPUT25), .ZN(n422) );
  XNOR2_X2 U521 ( .A(n425), .B(n424), .ZN(n608) );
  NAND2_X1 U522 ( .A1(G221), .A2(n426), .ZN(n427) );
  XNOR2_X1 U523 ( .A(KEYINPUT21), .B(n427), .ZN(n607) );
  XNOR2_X2 U524 ( .A(n428), .B(KEYINPUT88), .ZN(n548) );
  XNOR2_X1 U525 ( .A(n429), .B(KEYINPUT14), .ZN(n431) );
  NAND2_X1 U526 ( .A1(G952), .A2(n431), .ZN(n430) );
  XNOR2_X1 U527 ( .A(KEYINPUT82), .B(n430), .ZN(n632) );
  NOR2_X1 U528 ( .A1(G953), .A2(n632), .ZN(n542) );
  NAND2_X1 U529 ( .A1(G902), .A2(n431), .ZN(n539) );
  OR2_X1 U530 ( .A1(n733), .A2(n539), .ZN(n432) );
  NOR2_X1 U531 ( .A1(G900), .A2(n432), .ZN(n433) );
  OR2_X1 U532 ( .A1(n542), .A2(n433), .ZN(n493) );
  NAND2_X1 U533 ( .A1(n469), .A2(G210), .ZN(n435) );
  XNOR2_X1 U534 ( .A(n435), .B(G131), .ZN(n437) );
  XNOR2_X1 U535 ( .A(KEYINPUT89), .B(KEYINPUT5), .ZN(n436) );
  XNOR2_X1 U536 ( .A(n437), .B(n436), .ZN(n441) );
  INV_X1 U537 ( .A(G902), .ZN(n487) );
  NAND2_X1 U538 ( .A1(n487), .A2(n442), .ZN(n461) );
  NAND2_X1 U539 ( .A1(n461), .A2(G214), .ZN(n617) );
  NAND2_X1 U540 ( .A1(n515), .A2(n617), .ZN(n444) );
  XNOR2_X1 U541 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U543 ( .A(n447), .B(G122), .ZN(n448) );
  XNOR2_X1 U544 ( .A(n449), .B(n448), .ZN(n721) );
  XNOR2_X1 U545 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U546 ( .A(n455), .B(n454), .ZN(n459) );
  NAND2_X1 U547 ( .A1(n733), .A2(G224), .ZN(n456) );
  XNOR2_X1 U548 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U549 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U550 ( .A(n721), .B(n460), .ZN(n684) );
  NAND2_X1 U551 ( .A1(n684), .A2(n589), .ZN(n463) );
  AND2_X1 U552 ( .A1(n461), .A2(G210), .ZN(n462) );
  XNOR2_X2 U553 ( .A(n463), .B(n462), .ZN(n533) );
  INV_X1 U554 ( .A(KEYINPUT38), .ZN(n464) );
  INV_X1 U555 ( .A(n466), .ZN(n467) );
  XNOR2_X1 U556 ( .A(n468), .B(n467), .ZN(n730) );
  NAND2_X1 U557 ( .A1(G214), .A2(n469), .ZN(n470) );
  XNOR2_X1 U558 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U559 ( .A(n472), .B(KEYINPUT93), .Z(n474) );
  XNOR2_X1 U560 ( .A(n474), .B(n473), .ZN(n478) );
  XOR2_X1 U561 ( .A(KEYINPUT11), .B(KEYINPUT92), .Z(n476) );
  XNOR2_X1 U562 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U563 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U564 ( .A(n730), .B(n479), .ZN(n597) );
  NAND2_X1 U565 ( .A1(n597), .A2(n487), .ZN(n481) );
  XOR2_X1 U566 ( .A(KEYINPUT13), .B(G475), .Z(n480) );
  XOR2_X1 U567 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n483) );
  XNOR2_X1 U568 ( .A(G116), .B(G122), .ZN(n484) );
  XNOR2_X1 U569 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U570 ( .A1(n670), .A2(n487), .ZN(n488) );
  XNOR2_X1 U571 ( .A(n488), .B(G478), .ZN(n505) );
  NAND2_X1 U572 ( .A1(n509), .A2(n508), .ZN(n706) );
  NOR2_X1 U573 ( .A1(n537), .A2(n706), .ZN(n490) );
  XNOR2_X1 U574 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U575 ( .A(n490), .B(n489), .ZN(n661) );
  NAND2_X1 U576 ( .A1(n618), .A2(n617), .ZN(n621) );
  NOR2_X1 U577 ( .A1(n509), .A2(n505), .ZN(n551) );
  INV_X1 U578 ( .A(n551), .ZN(n620) );
  XNOR2_X1 U579 ( .A(n491), .B(KEYINPUT41), .ZN(n603) );
  INV_X1 U580 ( .A(n607), .ZN(n492) );
  AND2_X1 U581 ( .A1(n493), .A2(n492), .ZN(n494) );
  NAND2_X1 U582 ( .A1(n608), .A2(n494), .ZN(n496) );
  INV_X1 U583 ( .A(KEYINPUT69), .ZN(n495) );
  XNOR2_X1 U584 ( .A(n496), .B(n495), .ZN(n517) );
  INV_X1 U585 ( .A(n515), .ZN(n559) );
  INV_X1 U586 ( .A(KEYINPUT28), .ZN(n497) );
  XNOR2_X1 U587 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U588 ( .A1(n499), .A2(n524), .ZN(n512) );
  NOR2_X1 U589 ( .A1(n603), .A2(n512), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n500), .B(KEYINPUT42), .ZN(n742) );
  NOR2_X1 U591 ( .A1(n661), .A2(n742), .ZN(n502) );
  XOR2_X1 U592 ( .A(KEYINPUT78), .B(KEYINPUT46), .Z(n501) );
  XNOR2_X1 U593 ( .A(n502), .B(n501), .ZN(n528) );
  OR2_X1 U594 ( .A1(n504), .A2(n503), .ZN(n507) );
  AND2_X1 U595 ( .A1(n505), .A2(n509), .ZN(n570) );
  NAND2_X1 U596 ( .A1(n570), .A2(n533), .ZN(n506) );
  NOR2_X1 U597 ( .A1(n507), .A2(n506), .ZN(n702) );
  XNOR2_X2 U598 ( .A(n510), .B(KEYINPUT97), .ZN(n622) );
  XNOR2_X1 U599 ( .A(KEYINPUT71), .B(KEYINPUT19), .ZN(n511) );
  NOR2_X1 U600 ( .A1(n622), .A2(n703), .ZN(n513) );
  XOR2_X1 U601 ( .A(KEYINPUT47), .B(n513), .Z(n514) );
  NOR2_X1 U602 ( .A1(n702), .A2(n514), .ZN(n526) );
  XNOR2_X1 U603 ( .A(KEYINPUT98), .B(KEYINPUT6), .ZN(n516) );
  OR2_X1 U604 ( .A1(n517), .A2(n563), .ZN(n518) );
  XNOR2_X1 U605 ( .A(n518), .B(KEYINPUT101), .ZN(n521) );
  INV_X1 U606 ( .A(n617), .ZN(n519) );
  NOR2_X1 U607 ( .A1(n706), .A2(n519), .ZN(n520) );
  NAND2_X1 U608 ( .A1(n531), .A2(n533), .ZN(n523) );
  XOR2_X1 U609 ( .A(KEYINPUT80), .B(KEYINPUT36), .Z(n522) );
  XNOR2_X1 U610 ( .A(n523), .B(n522), .ZN(n525) );
  NAND2_X1 U611 ( .A1(n525), .A2(n345), .ZN(n660) );
  NAND2_X1 U612 ( .A1(n526), .A2(n660), .ZN(n527) );
  NOR2_X1 U613 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U614 ( .A(n345), .ZN(n530) );
  NAND2_X1 U615 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U616 ( .A(n532), .B(KEYINPUT43), .ZN(n535) );
  INV_X1 U617 ( .A(n533), .ZN(n534) );
  AND2_X1 U618 ( .A1(n535), .A2(n534), .ZN(n712) );
  OR2_X1 U619 ( .A1(n537), .A2(n536), .ZN(n655) );
  INV_X1 U620 ( .A(n732), .ZN(n639) );
  NAND2_X1 U621 ( .A1(n639), .A2(KEYINPUT2), .ZN(n584) );
  XOR2_X1 U622 ( .A(KEYINPUT31), .B(KEYINPUT90), .Z(n547) );
  INV_X1 U623 ( .A(G953), .ZN(n715) );
  NOR2_X1 U624 ( .A1(n715), .A2(G898), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n538), .B(KEYINPUT83), .ZN(n724) );
  NOR2_X1 U626 ( .A1(n539), .A2(n724), .ZN(n540) );
  XNOR2_X1 U627 ( .A(n540), .B(KEYINPUT84), .ZN(n541) );
  NOR2_X1 U628 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U629 ( .A(KEYINPUT0), .ZN(n545) );
  INV_X1 U630 ( .A(n569), .ZN(n550) );
  NOR2_X1 U631 ( .A1(n548), .A2(n610), .ZN(n549) );
  NAND2_X1 U632 ( .A1(n550), .A2(n549), .ZN(n694) );
  INV_X1 U633 ( .A(n608), .ZN(n562) );
  NAND2_X1 U634 ( .A1(n563), .A2(n562), .ZN(n552) );
  OR2_X1 U635 ( .A1(n552), .A2(n345), .ZN(n553) );
  NOR2_X1 U636 ( .A1(n558), .A2(n553), .ZN(n691) );
  NAND2_X1 U637 ( .A1(n608), .A2(n345), .ZN(n554) );
  XNOR2_X1 U638 ( .A(KEYINPUT99), .B(n554), .ZN(n555) );
  NAND2_X1 U639 ( .A1(n555), .A2(n563), .ZN(n556) );
  NOR2_X1 U640 ( .A1(n558), .A2(n556), .ZN(n557) );
  XNOR2_X1 U641 ( .A(n557), .B(KEYINPUT32), .ZN(n743) );
  NOR2_X1 U642 ( .A1(n558), .A2(n345), .ZN(n560) );
  NAND2_X1 U643 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X2 U644 ( .A1(n562), .A2(n561), .ZN(n656) );
  NOR2_X1 U645 ( .A1(n743), .A2(n656), .ZN(n574) );
  INV_X1 U646 ( .A(n563), .ZN(n564) );
  XNOR2_X1 U647 ( .A(KEYINPUT100), .B(KEYINPUT33), .ZN(n567) );
  INV_X1 U648 ( .A(KEYINPUT70), .ZN(n566) );
  XNOR2_X1 U649 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U650 ( .A1(n571), .A2(n570), .ZN(n573) );
  INV_X1 U651 ( .A(KEYINPUT35), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n574), .A2(n658), .ZN(n578) );
  XNOR2_X1 U653 ( .A(n577), .B(KEYINPUT79), .ZN(n582) );
  INV_X1 U654 ( .A(n578), .ZN(n580) );
  INV_X1 U655 ( .A(KEYINPUT44), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X2 U658 ( .A(n583), .B(KEYINPUT45), .ZN(n714) );
  INV_X1 U659 ( .A(n714), .ZN(n646) );
  NOR2_X2 U660 ( .A1(n584), .A2(n646), .ZN(n643) );
  INV_X1 U661 ( .A(n643), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n585), .A2(n714), .ZN(n586) );
  INV_X1 U663 ( .A(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U664 ( .A1(n586), .A2(n644), .ZN(n588) );
  INV_X1 U665 ( .A(n589), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n732), .A2(n589), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n590), .A2(n714), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n591), .A2(KEYINPUT75), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n682), .A2(G475), .ZN(n599) );
  XNOR2_X1 U671 ( .A(KEYINPUT117), .B(KEYINPUT59), .ZN(n596) );
  XNOR2_X1 U672 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n600), .A2(n687), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(n601), .ZN(G60) );
  NOR2_X1 U676 ( .A1(n605), .A2(n345), .ZN(n606) );
  XOR2_X1 U677 ( .A(KEYINPUT50), .B(n606), .Z(n613) );
  NAND2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n609), .B(KEYINPUT49), .ZN(n611) );
  NOR2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U682 ( .A(KEYINPUT51), .B(n615), .Z(n616) );
  NOR2_X1 U683 ( .A1(n603), .A2(n616), .ZN(n628) );
  NOR2_X1 U684 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U685 ( .A1(n620), .A2(n619), .ZN(n624) );
  NOR2_X1 U686 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U687 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U688 ( .A1(n633), .A2(n625), .ZN(n626) );
  XNOR2_X1 U689 ( .A(n626), .B(KEYINPUT112), .ZN(n627) );
  NOR2_X1 U690 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U691 ( .A(n629), .B(KEYINPUT113), .Z(n630) );
  XNOR2_X1 U692 ( .A(KEYINPUT52), .B(n630), .ZN(n631) );
  NOR2_X1 U693 ( .A1(n632), .A2(n631), .ZN(n635) );
  NOR2_X1 U694 ( .A1(n603), .A2(n633), .ZN(n634) );
  NOR2_X1 U695 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U696 ( .A(n636), .B(KEYINPUT114), .ZN(n637) );
  NAND2_X1 U697 ( .A1(n637), .A2(n715), .ZN(n651) );
  NAND2_X1 U698 ( .A1(KEYINPUT73), .A2(n644), .ZN(n641) );
  NOR2_X1 U699 ( .A1(KEYINPUT73), .A2(n644), .ZN(n638) );
  NOR2_X1 U700 ( .A1(n639), .A2(n638), .ZN(n640) );
  AND2_X1 U701 ( .A1(n641), .A2(n640), .ZN(n642) );
  OR2_X1 U702 ( .A1(n643), .A2(n642), .ZN(n649) );
  XOR2_X1 U703 ( .A(KEYINPUT73), .B(n644), .Z(n645) );
  NAND2_X1 U704 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U705 ( .A(KEYINPUT74), .B(n647), .Z(n648) );
  NOR2_X1 U706 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U707 ( .A1(n651), .A2(n650), .ZN(n654) );
  INV_X1 U708 ( .A(KEYINPUT53), .ZN(n652) );
  XNOR2_X1 U709 ( .A(n652), .B(KEYINPUT115), .ZN(n653) );
  XNOR2_X1 U710 ( .A(n655), .B(G134), .ZN(G36) );
  XOR2_X1 U711 ( .A(G110), .B(n656), .Z(G12) );
  XNOR2_X1 U712 ( .A(G122), .B(KEYINPUT124), .ZN(n657) );
  XNOR2_X1 U713 ( .A(n658), .B(n657), .ZN(G24) );
  XOR2_X1 U714 ( .A(G125), .B(KEYINPUT37), .Z(n659) );
  XNOR2_X1 U715 ( .A(n660), .B(n659), .ZN(G27) );
  XOR2_X1 U716 ( .A(n661), .B(G131), .Z(G33) );
  NAND2_X1 U717 ( .A1(n682), .A2(G472), .ZN(n664) );
  XOR2_X1 U718 ( .A(KEYINPUT62), .B(n662), .Z(n663) );
  XNOR2_X1 U719 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U720 ( .A1(n665), .A2(n687), .ZN(n666) );
  XNOR2_X1 U721 ( .A(n666), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U722 ( .A1(n674), .A2(G217), .ZN(n668) );
  XNOR2_X1 U723 ( .A(n668), .B(n667), .ZN(n669) );
  INV_X1 U724 ( .A(n687), .ZN(n680) );
  NOR2_X1 U725 ( .A1(n669), .A2(n680), .ZN(G66) );
  NAND2_X1 U726 ( .A1(n674), .A2(G478), .ZN(n672) );
  XOR2_X1 U727 ( .A(KEYINPUT118), .B(n670), .Z(n671) );
  XNOR2_X1 U728 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U729 ( .A1(n673), .A2(n680), .ZN(G63) );
  NAND2_X1 U730 ( .A1(n674), .A2(G469), .ZN(n679) );
  XOR2_X1 U731 ( .A(KEYINPUT116), .B(KEYINPUT57), .Z(n676) );
  XNOR2_X1 U732 ( .A(n676), .B(KEYINPUT58), .ZN(n677) );
  XNOR2_X1 U733 ( .A(n675), .B(n677), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n679), .B(n678), .ZN(n681) );
  NOR2_X1 U735 ( .A1(n681), .A2(n680), .ZN(G54) );
  NAND2_X1 U736 ( .A1(n682), .A2(G210), .ZN(n686) );
  XOR2_X1 U737 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n683) );
  XNOR2_X1 U738 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U739 ( .A(n686), .B(n685), .ZN(n688) );
  NAND2_X1 U740 ( .A1(n688), .A2(n687), .ZN(n690) );
  XNOR2_X1 U741 ( .A(KEYINPUT77), .B(KEYINPUT56), .ZN(n689) );
  XNOR2_X1 U742 ( .A(n690), .B(n689), .ZN(G51) );
  XOR2_X1 U743 ( .A(G101), .B(n691), .Z(G3) );
  NOR2_X1 U744 ( .A1(n694), .A2(n706), .ZN(n693) );
  XNOR2_X1 U745 ( .A(G104), .B(KEYINPUT105), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n693), .B(n692), .ZN(G6) );
  NOR2_X1 U747 ( .A1(n694), .A2(n709), .ZN(n699) );
  XOR2_X1 U748 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n696) );
  XNOR2_X1 U749 ( .A(G107), .B(KEYINPUT26), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U751 ( .A(KEYINPUT27), .B(n697), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(G9) );
  NOR2_X1 U753 ( .A1(n709), .A2(n703), .ZN(n701) );
  XNOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(G30) );
  XOR2_X1 U756 ( .A(n343), .B(n702), .Z(G45) );
  NOR2_X1 U757 ( .A1(n706), .A2(n703), .ZN(n704) );
  XOR2_X1 U758 ( .A(KEYINPUT108), .B(n704), .Z(n705) );
  XNOR2_X1 U759 ( .A(G146), .B(n705), .ZN(G48) );
  XNOR2_X1 U760 ( .A(G113), .B(KEYINPUT109), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(G15) );
  XOR2_X1 U762 ( .A(KEYINPUT110), .B(n710), .Z(n711) );
  XNOR2_X1 U763 ( .A(G116), .B(n711), .ZN(G18) );
  XNOR2_X1 U764 ( .A(G140), .B(n712), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n713), .B(KEYINPUT111), .ZN(G42) );
  BUF_X1 U766 ( .A(n714), .Z(n716) );
  NAND2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U768 ( .A1(G953), .A2(G224), .ZN(n717) );
  XNOR2_X1 U769 ( .A(KEYINPUT61), .B(n717), .ZN(n718) );
  NAND2_X1 U770 ( .A1(n718), .A2(G898), .ZN(n719) );
  NAND2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n728) );
  XNOR2_X1 U772 ( .A(n721), .B(KEYINPUT119), .ZN(n722) );
  XNOR2_X1 U773 ( .A(n722), .B(KEYINPUT120), .ZN(n723) );
  XNOR2_X1 U774 ( .A(G101), .B(n723), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n726), .B(KEYINPUT121), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(G69) );
  XNOR2_X1 U778 ( .A(n730), .B(KEYINPUT122), .ZN(n731) );
  XOR2_X1 U779 ( .A(n729), .B(n731), .Z(n735) );
  XNOR2_X1 U780 ( .A(n732), .B(n735), .ZN(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(n739) );
  XNOR2_X1 U782 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U783 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U784 ( .A1(G953), .A2(n737), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U786 ( .A(KEYINPUT123), .B(n740), .Z(G72) );
  XOR2_X1 U787 ( .A(G137), .B(KEYINPUT126), .Z(n741) );
  XNOR2_X1 U788 ( .A(n742), .B(n741), .ZN(G39) );
  XNOR2_X1 U789 ( .A(G119), .B(KEYINPUT125), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(n743), .ZN(G21) );
endmodule

