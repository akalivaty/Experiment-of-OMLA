//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  AND2_X1   g000(.A1(KEYINPUT71), .A2(G953), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT71), .A2(G953), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT76), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n196), .A2(new_n198), .A3(new_n203), .A4(new_n199), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(KEYINPUT66), .A3(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  AOI21_X1  g025(.A(G128), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT67), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(G128), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n215), .A2(new_n220), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT77), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G104), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n229), .B(G101), .C1(new_n224), .C2(new_n228), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G107), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G107), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(G104), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G107), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n225), .A3(new_n227), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n223), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n222), .A2(new_n209), .A3(new_n211), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(new_n217), .C1(G128), .C2(new_n219), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n230), .A3(new_n237), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n207), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n234), .A2(new_n225), .A3(new_n227), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G107), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n234), .B2(new_n224), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT0), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(new_n221), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n219), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n251), .A3(new_n221), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n210), .A2(G146), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n256), .B(new_n258), .C1(new_n259), .C2(new_n216), .ZN(new_n260));
  OAI211_X1 g074(.A(KEYINPUT65), .B(new_n252), .C1(new_n259), .C2(new_n216), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n255), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n236), .B1(new_n233), .B2(new_n235), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n250), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n238), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n215), .A2(new_n220), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n240), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT78), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n242), .A2(new_n272), .A3(new_n267), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n242), .B2(new_n267), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n266), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n207), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n193), .B1(new_n245), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n193), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n275), .B2(new_n276), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n280), .A2(KEYINPUT79), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n276), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n280), .B2(KEYINPUT79), .ZN(new_n283));
  OAI211_X1 g097(.A(G469), .B(new_n278), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n245), .A2(new_n280), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n265), .A2(new_n262), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n288), .A2(new_n250), .B1(new_n268), .B2(new_n270), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n289), .B(new_n207), .C1(new_n273), .C2(new_n274), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n279), .B1(new_n282), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n285), .A2(new_n286), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n284), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT9), .B(G234), .ZN(new_n296));
  OAI21_X1  g110(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n297), .B(KEYINPUT75), .Z(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G952), .ZN(new_n301));
  AOI211_X1 g115(.A(G953), .B(new_n301), .C1(G234), .C2(G237), .ZN(new_n302));
  INV_X1    g116(.A(new_n189), .ZN(new_n303));
  NAND2_X1  g117(.A1(G234), .A2(G237), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n303), .A2(G902), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT21), .B(G898), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G113), .B(G122), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(new_n224), .ZN(new_n310));
  INV_X1    g124(.A(G237), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n189), .A2(G214), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n210), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n189), .A2(G143), .A3(G214), .A4(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G131), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n203), .A3(new_n314), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT89), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT89), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n320), .A3(new_n317), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  OR3_X1    g138(.A1(new_n324), .A2(KEYINPUT16), .A3(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(G146), .A3(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n322), .B(KEYINPUT19), .Z(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G146), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n321), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n315), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n315), .A2(new_n331), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n322), .B(new_n208), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n310), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n310), .B(KEYINPUT90), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT17), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n316), .A2(new_n338), .A3(new_n317), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n323), .A2(new_n325), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n208), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n326), .C1(new_n316), .C2(new_n338), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n335), .B(new_n337), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n336), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(G475), .A2(G902), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n347), .C1(new_n336), .C2(new_n345), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n352));
  INV_X1    g166(.A(new_n343), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n339), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n344), .B1(new_n354), .B2(new_n310), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n286), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n349), .A2(new_n351), .B1(G475), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G478), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(KEYINPUT15), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n361));
  INV_X1    g175(.A(G122), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(G116), .ZN(new_n363));
  INV_X1    g177(.A(G116), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(KEYINPUT91), .A3(G122), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(G116), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G107), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(G107), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n360), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n210), .A2(G128), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n221), .A2(G143), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n195), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT13), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n210), .A3(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n374), .ZN(new_n378));
  OAI211_X1 g192(.A(G134), .B(new_n377), .C1(new_n378), .C2(new_n376), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT93), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n366), .A2(new_n367), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n228), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT92), .A3(new_n369), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n372), .A2(new_n375), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n366), .A2(KEYINPUT14), .B1(G116), .B2(new_n362), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n385), .A2(KEYINPUT95), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n385), .B2(KEYINPUT95), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n228), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n371), .A2(KEYINPUT94), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n371), .A2(KEYINPUT94), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n378), .A2(G134), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n375), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n384), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G217), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n296), .A2(new_n396), .A3(G953), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n384), .B(new_n397), .C1(new_n389), .C2(new_n394), .ZN(new_n400));
  AOI21_X1  g214(.A(G902), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n359), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n401), .A2(KEYINPUT96), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n405));
  AOI211_X1 g219(.A(new_n405), .B(G902), .C1(new_n399), .C2(new_n400), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n403), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n391), .A2(new_n393), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n386), .A2(new_n388), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n390), .B(new_n408), .C1(new_n409), .C2(new_n228), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n397), .B1(new_n410), .B2(new_n384), .ZN(new_n411));
  INV_X1    g225(.A(new_n400), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n286), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n359), .B1(new_n413), .B2(new_n402), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n300), .A2(new_n308), .A3(new_n357), .A4(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G122), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n364), .A2(G119), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT68), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n364), .B2(G119), .ZN(new_n422));
  INV_X1    g236(.A(G119), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n423), .A2(KEYINPUT68), .A3(G116), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT2), .B(G113), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT68), .B1(new_n423), .B2(G116), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n364), .A3(G119), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n419), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n426), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n427), .A2(new_n432), .B1(new_n263), .B2(new_n264), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n230), .A2(new_n237), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT5), .B(new_n420), .C1(new_n422), .C2(new_n424), .ZN(new_n435));
  INV_X1    g249(.A(G113), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n419), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n435), .A2(new_n438), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n433), .A2(new_n250), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n418), .B1(new_n440), .B2(KEYINPUT80), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n433), .A2(new_n250), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n434), .A2(new_n439), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT81), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n427), .A2(new_n432), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n265), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n440), .A2(KEYINPUT80), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n418), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n440), .A2(new_n417), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n458));
  NAND4_X1  g272(.A1(new_n451), .A2(new_n452), .A3(new_n458), .A4(new_n418), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n270), .A2(new_n324), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n262), .A2(G125), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G224), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G953), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n462), .B(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n457), .A2(new_n459), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(KEYINPUT7), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n460), .A2(new_n461), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n455), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n417), .B(KEYINPUT8), .Z(new_n471));
  XNOR2_X1  g285(.A(new_n438), .B(KEYINPUT83), .ZN(new_n472));
  INV_X1    g286(.A(new_n435), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n432), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n474), .B2(new_n434), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n439), .A2(new_n238), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(new_n465), .B2(KEYINPUT84), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(KEYINPUT84), .B2(new_n465), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n475), .A2(new_n476), .B1(new_n462), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT86), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n467), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n480), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n482), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G214), .B1(G237), .B2(G902), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n483), .B1(new_n487), .B2(KEYINPUT85), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n493), .B(new_n485), .C1(KEYINPUT85), .C2(new_n487), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT88), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n491), .A2(new_n497), .A3(new_n494), .A4(new_n492), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n416), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G472), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT72), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n205), .A2(new_n262), .A3(new_n206), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n205), .A2(new_n262), .A3(KEYINPUT69), .A4(new_n206), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n446), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n195), .A2(G137), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n197), .A2(G134), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n204), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n270), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n506), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n507), .B1(new_n506), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n501), .B(KEYINPUT28), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n506), .A2(new_n514), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n446), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n504), .A2(new_n505), .B1(new_n270), .B2(new_n513), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n507), .A3(new_n502), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n517), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n189), .A2(G210), .A3(new_n311), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT27), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n502), .B1(new_n223), .B2(new_n511), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n536), .A2(new_n446), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n515), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(new_n525), .A3(new_n531), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n502), .B(new_n540), .C1(new_n223), .C2(new_n511), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n521), .B2(new_n540), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n515), .B1(new_n542), .B2(new_n446), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n539), .B(new_n533), .C1(new_n531), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n500), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n531), .B1(new_n538), .B2(new_n525), .ZN(new_n546));
  INV_X1    g360(.A(new_n541), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n519), .B2(KEYINPUT30), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n522), .B(new_n531), .C1(new_n548), .C2(new_n507), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT31), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(KEYINPUT31), .A3(new_n531), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G472), .A2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT32), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n538), .A2(new_n525), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n532), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n542), .A2(new_n446), .ZN(new_n559));
  AND4_X1   g373(.A1(KEYINPUT31), .A2(new_n559), .A3(new_n522), .A4(new_n531), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT31), .B1(new_n543), .B2(new_n531), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n554), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n545), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n396), .B1(G234), .B2(new_n286), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n342), .A2(new_n326), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT73), .B1(new_n423), .B2(G128), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT73), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n221), .A3(G119), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n423), .A2(G128), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G110), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n423), .B2(G128), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n578), .A2(new_n579), .A3(new_n572), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n568), .B(new_n575), .C1(new_n576), .C2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n326), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT74), .B(G110), .Z(new_n583));
  AOI22_X1  g397(.A1(new_n580), .A2(new_n583), .B1(new_n573), .B2(new_n574), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n322), .A2(new_n208), .ZN(new_n585));
  OR3_X1    g399(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT22), .B(G137), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n586), .A3(new_n590), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n286), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT25), .A4(new_n286), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n567), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n592), .A2(new_n593), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n566), .A2(G902), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n599), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n565), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n499), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  AOI21_X1  g420(.A(new_n483), .B1(new_n467), .B2(new_n480), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n492), .B1(new_n484), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT98), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n413), .A2(new_n405), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n401), .A2(KEYINPUT96), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n358), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n398), .B2(KEYINPUT99), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n411), .B2(new_n412), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n399), .A2(new_n400), .A3(new_n614), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(G478), .A3(new_n286), .A4(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n357), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n621), .B(new_n492), .C1(new_n484), .C2(new_n607), .ZN(new_n622));
  AND4_X1   g436(.A1(new_n308), .A2(new_n609), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n603), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n300), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G472), .B1(new_n553), .B2(G902), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n553), .B2(new_n555), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND2_X1  g446(.A1(new_n487), .A2(new_n482), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n467), .A2(new_n480), .A3(new_n483), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n621), .B1(new_n635), .B2(new_n492), .ZN(new_n636));
  INV_X1    g450(.A(new_n622), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n356), .A2(G475), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n328), .B1(new_n318), .B2(KEYINPUT89), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n352), .B1(new_n640), .B2(new_n321), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n344), .B1(new_n641), .B2(new_n310), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n350), .B1(new_n642), .B2(new_n347), .ZN(new_n643));
  INV_X1    g457(.A(new_n351), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n415), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n628), .A2(new_n638), .A3(new_n308), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n587), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n601), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n598), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n627), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n499), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n302), .B1(new_n305), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n415), .A2(new_n645), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n609), .A2(new_n661), .A3(new_n622), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n654), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n300), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n565), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XOR2_X1   g482(.A(new_n660), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n300), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT103), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n670), .B(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n672), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n415), .A2(new_n357), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n492), .A3(new_n654), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n673), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n556), .A2(new_n564), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n520), .A2(new_n522), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n500), .B1(new_n682), .B2(new_n532), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n683), .A2(new_n549), .B1(G472), .B2(G902), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n681), .A2(KEYINPUT102), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT102), .B1(new_n681), .B2(new_n686), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n491), .A2(new_n494), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT38), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n680), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n210), .ZN(G45));
  INV_X1    g510(.A(new_n545), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n681), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n300), .A2(new_n664), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n612), .A2(new_n618), .ZN(new_n701));
  INV_X1    g515(.A(new_n660), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n701), .A2(new_n645), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n609), .A2(new_n703), .A3(new_n622), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n609), .A2(new_n703), .A3(KEYINPUT105), .A4(new_n622), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n208), .ZN(G48));
  OAI21_X1  g523(.A(new_n286), .B1(new_n287), .B2(new_n291), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  INV_X1    g525(.A(new_n292), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n299), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n565), .A2(new_n603), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n623), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR3_X1   g532(.A1(new_n711), .A2(new_n712), .A3(new_n298), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n415), .A2(new_n603), .A3(new_n645), .A4(new_n307), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n638), .A2(new_n698), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NAND2_X1  g536(.A1(new_n415), .A2(new_n357), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n307), .A3(new_n654), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n638), .A2(new_n698), .A3(new_n719), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT106), .B(G119), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G21));
  AND3_X1   g541(.A1(new_n609), .A2(new_n622), .A3(new_n678), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT107), .B(G472), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n562), .B2(new_n286), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n710), .A2(G469), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n299), .A3(new_n292), .A4(new_n308), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n551), .A2(new_n552), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n517), .B(new_n532), .C1(new_n523), .C2(new_n526), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n555), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n731), .A2(new_n733), .A3(new_n736), .A4(new_n603), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n728), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NAND4_X1  g553(.A1(new_n609), .A2(new_n703), .A3(new_n622), .A4(new_n719), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n731), .A2(new_n736), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n664), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n324), .ZN(G27));
  INV_X1    g558(.A(new_n492), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n491), .B2(new_n494), .ZN(new_n746));
  AND4_X1   g560(.A1(KEYINPUT42), .A2(new_n746), .A3(new_n300), .A4(new_n703), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n681), .A2(KEYINPUT108), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n556), .A2(new_n564), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n697), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n751), .A2(new_n752), .A3(new_n624), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n751), .B2(new_n624), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n747), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n746), .A2(new_n604), .A3(new_n300), .A4(new_n703), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  AND4_X1   g574(.A1(new_n604), .A2(new_n746), .A3(new_n300), .A4(new_n661), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n195), .ZN(G36));
  INV_X1    g576(.A(new_n746), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n619), .A2(new_n645), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT43), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n765), .A2(new_n627), .A3(new_n664), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n763), .B1(new_n766), .B2(KEYINPUT44), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(KEYINPUT44), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n278), .B1(new_n281), .B2(new_n283), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n285), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n772));
  OAI22_X1  g586(.A1(new_n771), .A2(new_n772), .B1(new_n770), .B2(new_n769), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n294), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n712), .B1(new_n775), .B2(new_n777), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n299), .A3(new_n669), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n768), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n299), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT47), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n746), .A2(new_n565), .A3(new_n603), .A4(new_n703), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  AND4_X1   g603(.A1(new_n624), .A2(new_n765), .A3(new_n302), .A4(new_n741), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n714), .A2(new_n492), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n693), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n763), .A2(new_n714), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n624), .A3(new_n690), .A4(new_n302), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT118), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT118), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n357), .A3(new_n619), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n302), .A3(new_n765), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n800), .A2(KEYINPUT117), .A3(new_n742), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT117), .B1(new_n800), .B2(new_n742), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n794), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n713), .A2(new_n298), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n786), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n746), .A3(new_n790), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n804), .A2(new_n807), .A3(KEYINPUT51), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n753), .A2(new_n754), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n302), .A3(new_n765), .A4(new_n795), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT48), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n797), .A2(new_n620), .A3(new_n798), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n636), .A2(new_n637), .A3(new_n714), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n301), .B(G953), .C1(new_n790), .C2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n810), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT119), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n810), .A2(new_n821), .A3(new_n811), .A4(new_n818), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n716), .A2(new_n721), .A3(new_n725), .A4(new_n738), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT112), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n816), .B(new_n698), .C1(new_n720), .C2(new_n724), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n716), .A4(new_n738), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n496), .A2(new_n498), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n620), .A2(new_n646), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n831), .A2(new_n625), .A3(new_n627), .A4(new_n307), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n605), .A2(new_n656), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n761), .B1(new_n755), .B2(new_n758), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n565), .A2(new_n723), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n620), .B2(new_n741), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n746), .A2(new_n300), .A3(new_n664), .A4(new_n702), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n829), .A2(new_n834), .A3(new_n835), .A4(new_n840), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n700), .A2(new_n662), .B1(new_n740), .B2(new_n742), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n708), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n598), .A2(new_n653), .A3(new_n660), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n295), .A2(new_n299), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n609), .A2(new_n622), .A3(new_n678), .A4(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n553), .A2(KEYINPUT32), .A3(new_n555), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n563), .B1(new_n562), .B2(new_n554), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n686), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT102), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n846), .B1(new_n851), .B2(new_n687), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n843), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n708), .A2(new_n842), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n841), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n854), .B2(new_n856), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n499), .A2(new_n604), .B1(new_n830), .B2(new_n832), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n656), .A2(new_n825), .A3(new_n862), .A4(new_n828), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n706), .A2(new_n707), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n666), .ZN(new_n865));
  INV_X1    g679(.A(new_n740), .ZN(new_n866));
  INV_X1    g680(.A(new_n742), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n866), .A2(new_n867), .B1(new_n663), .B2(new_n666), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n868), .A3(new_n853), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n855), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n853), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(KEYINPUT113), .A3(new_n871), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n761), .B(new_n839), .C1(new_n755), .C2(new_n758), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n861), .A2(new_n863), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT54), .B1(new_n859), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n824), .B(KEYINPUT116), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(KEYINPUT53), .A3(new_n834), .ZN(new_n879));
  INV_X1    g693(.A(new_n873), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n857), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n874), .A2(new_n883), .A3(new_n875), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n874), .B2(new_n875), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n877), .B1(new_n886), .B2(KEYINPUT54), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n823), .A2(new_n887), .B1(G952), .B2(G953), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n624), .A2(new_n764), .A3(new_n492), .A4(new_n299), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n713), .B(KEYINPUT49), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n693), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n691), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n189), .A2(G952), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT121), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n886), .A2(G902), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n896), .B2(new_n483), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n457), .A2(new_n459), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n466), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n894), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n897), .B2(new_n902), .ZN(G51));
  NOR2_X1   g718(.A1(new_n287), .A2(new_n291), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT122), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n861), .A2(new_n872), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n875), .B1(new_n907), .B2(new_n841), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT115), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n874), .A2(new_n883), .A3(new_n875), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n881), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT54), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n293), .B(KEYINPUT57), .Z(new_n913));
  OAI21_X1  g727(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n896), .A2(new_n774), .A3(new_n773), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n893), .B1(new_n914), .B2(new_n915), .ZN(G54));
  NAND4_X1  g730(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n346), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n346), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n893), .ZN(G60));
  AND2_X1   g734(.A1(new_n616), .A2(new_n617), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT59), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n894), .B1(new_n912), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n887), .B2(new_n923), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(G63));
  XNOR2_X1  g741(.A(new_n600), .B(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n911), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n930), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n886), .A2(new_n651), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n894), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n934), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT61), .B1(new_n934), .B2(KEYINPUT123), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  NOR2_X1   g751(.A1(new_n863), .A2(new_n303), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT125), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n306), .B2(new_n463), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n898), .B1(G898), .B2(new_n189), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n944));
  INV_X1    g758(.A(new_n843), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n695), .B2(new_n945), .ZN(new_n946));
  OR3_X1    g760(.A1(new_n695), .A2(new_n944), .A3(new_n945), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n671), .A2(new_n763), .A3(new_n831), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n946), .A2(new_n947), .B1(new_n604), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n788), .A2(new_n783), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n303), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n542), .B(new_n327), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(KEYINPUT126), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  INV_X1    g770(.A(new_n954), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n954), .B1(G900), .B2(new_n303), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n812), .A2(new_n728), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n843), .B1(new_n960), .B2(new_n782), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n950), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n835), .A2(KEYINPUT127), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n835), .A2(KEYINPUT127), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n959), .B1(new_n965), .B2(new_n303), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n955), .A2(new_n958), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n968), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n955), .A2(new_n958), .A3(new_n970), .A4(new_n966), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(G72));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  INV_X1    g788(.A(new_n863), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n965), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n532), .A3(new_n543), .ZN(new_n977));
  INV_X1    g791(.A(new_n549), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n543), .A2(new_n531), .ZN(new_n979));
  OAI221_X1 g793(.A(new_n974), .B1(new_n978), .B2(new_n979), .C1(new_n859), .C2(new_n876), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n949), .A2(new_n863), .A3(new_n951), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n974), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n543), .A2(new_n532), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n893), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n977), .A2(new_n980), .A3(new_n984), .ZN(G57));
endmodule


