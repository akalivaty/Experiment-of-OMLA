//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n651,
    new_n652, new_n655, new_n657, new_n658, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT65), .B(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  OAI22_X1  g050(.A1(new_n471), .A2(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n477), .B1(new_n468), .B2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(KEYINPUT65), .B(G2105), .Z(new_n480));
  AOI21_X1  g055(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n468), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n469), .A2(new_n480), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n486), .B2(KEYINPUT66), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(KEYINPUT66), .B2(new_n486), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT67), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND3_X1  g067(.A1(new_n469), .A2(G138), .A3(new_n470), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n468), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n475), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n497), .A2(G2105), .B1(G102), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n506), .A2(new_n511), .A3(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n511), .A2(G50), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n506), .A2(G62), .ZN(new_n520));
  INV_X1    g095(.A(G75), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n521), .B2(new_n504), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n519), .B1(new_n522), .B2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n516), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n508), .A2(new_n510), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n534), .A2(G51), .A3(G543), .A4(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n538), .B1(new_n503), .B2(new_n505), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n502), .A2(G543), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT69), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G63), .A2(G651), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n537), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AOI211_X1 g121(.A(KEYINPUT70), .B(new_n544), .C1(new_n539), .C2(new_n542), .ZN(new_n547));
  OAI211_X1 g122(.A(KEYINPUT72), .B(new_n536), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT69), .ZN(new_n550));
  AOI21_X1  g125(.A(KEYINPUT69), .B1(new_n540), .B2(new_n541), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT70), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n543), .A2(new_n537), .A3(new_n545), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT72), .B1(new_n555), .B2(new_n536), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n532), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(G168));
  NAND2_X1  g133(.A1(new_n543), .A2(G64), .ZN(new_n559));
  NAND2_X1  g134(.A1(G77), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n507), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n534), .A2(G52), .A3(G543), .A4(new_n535), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n514), .A2(G90), .A3(new_n515), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n564), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT73), .B1(new_n567), .B2(new_n561), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G171));
  INV_X1    g144(.A(G81), .ZN(new_n570));
  INV_X1    g145(.A(G43), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n534), .A2(G543), .A3(new_n535), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n516), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n543), .A2(G56), .ZN(new_n574));
  NAND2_X1  g149(.A1(G68), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n507), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G860), .ZN(G153));
  AND3_X1   g153(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G36), .ZN(G176));
  NAND2_X1  g155(.A1(G1), .A2(G3), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT8), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(G188));
  INV_X1    g158(.A(new_n515), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT68), .B1(new_n506), .B2(new_n511), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT74), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n514), .A2(new_n587), .A3(new_n515), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(G65), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(G65), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n506), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G78), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n504), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n589), .A2(G91), .B1(G651), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n535), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT9), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT76), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n584), .A2(KEYINPUT74), .A3(new_n585), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n587), .B1(new_n514), .B2(new_n515), .ZN(new_n601));
  OAI21_X1  g176(.A(G91), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(G651), .ZN(new_n603));
  AND4_X1   g178(.A1(KEYINPUT76), .A2(new_n602), .A3(new_n598), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G299));
  AND2_X1   g181(.A1(new_n566), .A2(new_n568), .ZN(G301));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n557), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n536), .B1(new_n546), .B2(new_n547), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT72), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n548), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n613), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(G286));
  NAND2_X1  g190(.A1(new_n589), .A2(G87), .ZN(new_n616));
  OAI21_X1  g191(.A(G651), .B1(new_n543), .B2(G74), .ZN(new_n617));
  INV_X1    g192(.A(new_n572), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G49), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(G288));
  NAND2_X1  g195(.A1(new_n506), .A2(G61), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(KEYINPUT78), .B2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G651), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT80), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n589), .B2(G86), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n626), .A2(new_n629), .ZN(G305));
  INV_X1    g205(.A(G85), .ZN(new_n631));
  INV_X1    g206(.A(G47), .ZN(new_n632));
  OAI22_X1  g207(.A1(new_n516), .A2(new_n631), .B1(new_n632), .B2(new_n572), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n543), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n634), .A2(new_n507), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G290));
  NAND2_X1  g212(.A1(G301), .A2(G868), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n639));
  OAI211_X1 g214(.A(G92), .B(new_n639), .C1(new_n600), .C2(new_n601), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n506), .A2(G66), .ZN(new_n641));
  NAND2_X1  g216(.A1(G79), .A2(G543), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT82), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n507), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n618), .B2(G54), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n639), .B1(new_n589), .B2(G92), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n638), .B1(G868), .B2(new_n648), .ZN(G284));
  OAI21_X1  g224(.A(new_n638), .B1(G868), .B2(new_n648), .ZN(G321));
  NAND2_X1  g225(.A1(G286), .A2(G868), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(G868), .B2(new_n605), .ZN(new_n652));
  MUX2_X1   g227(.A(new_n651), .B(new_n652), .S(KEYINPUT83), .Z(G297));
  MUX2_X1   g228(.A(new_n651), .B(new_n652), .S(KEYINPUT83), .Z(G280));
  INV_X1    g229(.A(G559), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n648), .B1(new_n655), .B2(G860), .ZN(G148));
  NAND2_X1  g231(.A1(new_n648), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G868), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(G868), .B2(new_n577), .ZN(G323));
  XNOR2_X1  g234(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g235(.A1(new_n482), .A2(G135), .ZN(new_n661));
  OAI221_X1 g236(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n662));
  INV_X1    g237(.A(G123), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n484), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(G2096), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n468), .A2(new_n475), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT13), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n670), .ZN(G156));
  INV_X1    g246(.A(G14), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT15), .B(G2435), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2438), .ZN(new_n674));
  XOR2_X1   g249(.A(G2427), .B(G2430), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2451), .B(G2454), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT16), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2443), .B(G2446), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1341), .B(G1348), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n672), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n691), .C1(new_n689), .C2(new_n688), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n685), .B(new_n686), .ZN(new_n693));
  INV_X1    g268(.A(new_n689), .ZN(new_n694));
  OAI21_X1  g269(.A(G14), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n688), .A2(new_n689), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT87), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g274(.A(G2084), .B(G2090), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G2067), .B(G2678), .Z(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G2072), .A2(G2078), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n444), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT18), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(KEYINPUT17), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n701), .A2(new_n702), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n708), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n711));
  INV_X1    g286(.A(new_n705), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n707), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2100), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT90), .B(G2096), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(G227));
  XNOR2_X1  g293(.A(G1971), .B(G1976), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT19), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(G1956), .B(G2474), .Z(new_n722));
  XOR2_X1   g297(.A(G1961), .B(G1966), .Z(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n724), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n719), .B(KEYINPUT19), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n722), .A2(new_n723), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT91), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n731), .A2(new_n721), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n725), .B(new_n729), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n734), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1991), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1996), .ZN(new_n738));
  XNOR2_X1  g313(.A(G1981), .B(G1986), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(G229));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n648), .B2(new_n744), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1348), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(G19), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n577), .B2(new_n744), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1341), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n751), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n750), .B1(new_n754), .B2(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n469), .A2(new_n480), .A3(G128), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT93), .Z(new_n759));
  OR2_X1    g334(.A1(new_n470), .A2(G116), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n762), .A2(new_n763), .A3(new_n464), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n760), .A2(new_n764), .B1(new_n482), .B2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n757), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G2067), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n755), .B(new_n772), .C1(G2090), .C2(new_n754), .ZN(new_n773));
  INV_X1    g348(.A(G1956), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n744), .A2(G20), .ZN(new_n775));
  NAND2_X1  g350(.A1(G299), .A2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(KEYINPUT23), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(KEYINPUT23), .B2(new_n775), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n747), .B(new_n773), .C1(new_n774), .C2(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n774), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(G29), .A2(G33), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT25), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G139), .B2(new_n482), .ZN(new_n785));
  NAND2_X1  g360(.A1(G115), .A2(G2104), .ZN(new_n786));
  INV_X1    g361(.A(G127), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n468), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT96), .B1(new_n788), .B2(new_n480), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n788), .A2(KEYINPUT96), .A3(new_n480), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n782), .B1(new_n791), .B2(new_n751), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(new_n442), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT97), .ZN(new_n794));
  OR2_X1    g369(.A1(G29), .A2(G32), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n482), .A2(G141), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT99), .Z(new_n797));
  NAND3_X1  g372(.A1(new_n469), .A2(new_n480), .A3(G129), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT100), .Z(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT26), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n802), .A2(new_n803), .B1(G105), .B2(new_n498), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n797), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n795), .B1(new_n805), .B2(new_n751), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G34), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(KEYINPUT24), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(KEYINPUT24), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n751), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G160), .B2(new_n751), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT98), .ZN(new_n814));
  INV_X1    g389(.A(G2084), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n808), .B1(new_n792), .B2(new_n442), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n794), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT101), .Z(new_n818));
  INV_X1    g393(.A(KEYINPUT102), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(new_n815), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n806), .A2(new_n807), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n751), .A2(G27), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G164), .B2(new_n751), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(G2078), .ZN(new_n824));
  INV_X1    g399(.A(G28), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT30), .ZN(new_n826));
  AOI21_X1  g401(.A(G29), .B1(new_n825), .B2(KEYINPUT30), .ZN(new_n827));
  OR2_X1    g402(.A1(KEYINPUT31), .A2(G11), .ZN(new_n828));
  NAND2_X1  g403(.A1(KEYINPUT31), .A2(G11), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n826), .A2(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n664), .B2(new_n751), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n823), .B2(G2078), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n820), .A2(new_n821), .A3(new_n824), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n744), .A2(G5), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G171), .B2(new_n744), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(G1961), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n744), .A2(G21), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G168), .B2(new_n744), .ZN(new_n839));
  INV_X1    g414(.A(G1966), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n837), .B(new_n841), .C1(G1961), .C2(new_n835), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n818), .A2(new_n819), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n819), .B1(new_n818), .B2(new_n842), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n781), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G288), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G16), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G16), .B2(G23), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT33), .B(G1976), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n744), .A2(G22), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(G166), .B2(new_n744), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(G1971), .Z(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n744), .A2(G6), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G305), .B2(G16), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT32), .B(G1981), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT34), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n482), .A2(G131), .ZN(new_n863));
  OAI221_X1 g438(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n864));
  INV_X1    g439(.A(G119), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n484), .ZN(new_n866));
  MUX2_X1   g441(.A(G25), .B(new_n866), .S(G29), .Z(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G1991), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n867), .B(new_n868), .Z(new_n869));
  INV_X1    g444(.A(KEYINPUT36), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(KEYINPUT92), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n744), .A2(G24), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n636), .B2(new_n744), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(G1986), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(G1986), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n862), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n870), .A2(KEYINPUT92), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n877), .B(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n845), .A2(new_n880), .ZN(G311));
  XNOR2_X1  g456(.A(new_n877), .B(new_n878), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n882), .A2(new_n781), .A3(new_n843), .A4(new_n844), .ZN(G150));
  INV_X1    g458(.A(new_n647), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n640), .A3(new_n645), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(new_n655), .ZN(new_n886));
  XOR2_X1   g461(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G93), .ZN(new_n889));
  INV_X1    g464(.A(G55), .ZN(new_n890));
  OAI22_X1  g465(.A1(new_n516), .A2(new_n889), .B1(new_n890), .B2(new_n572), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n543), .A2(G67), .ZN(new_n892));
  NAND2_X1  g467(.A1(G80), .A2(G543), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n507), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n577), .B(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G860), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n888), .A2(new_n897), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n895), .A2(new_n899), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(G145));
  XOR2_X1   g479(.A(new_n791), .B(KEYINPUT103), .Z(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n805), .A2(new_n766), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n805), .A2(new_n766), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n500), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n500), .A3(new_n908), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n905), .B1(new_n913), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n482), .A2(G142), .ZN(new_n916));
  OAI221_X1 g491(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n917));
  INV_X1    g492(.A(G130), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n484), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n866), .B(new_n919), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(new_n668), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT104), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n922), .A2(KEYINPUT104), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(KEYINPUT104), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n925), .A2(new_n912), .A3(new_n914), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n479), .A2(new_n480), .ZN(new_n929));
  OAI221_X1 g504(.A(new_n929), .B1(new_n473), .B2(new_n475), .C1(new_n472), .C2(new_n471), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(new_n664), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(new_n491), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT105), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n928), .B2(new_n933), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n924), .A2(new_n927), .A3(new_n936), .A4(new_n932), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT106), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g518(.A(new_n885), .B1(new_n599), .B2(new_n604), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n602), .A2(new_n598), .A3(new_n603), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT76), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n596), .A2(KEYINPUT76), .A3(new_n598), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n648), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n944), .A2(KEYINPUT41), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT41), .B1(new_n944), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n944), .A2(new_n949), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n657), .B(new_n896), .ZN(new_n955));
  MUX2_X1   g530(.A(new_n952), .B(new_n954), .S(new_n955), .Z(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(G305), .B(new_n846), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n636), .B(G303), .Z(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n957), .A2(new_n958), .A3(new_n962), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(G868), .B2(new_n895), .ZN(G295));
  OAI21_X1  g542(.A(new_n966), .B1(G868), .B2(new_n895), .ZN(G331));
  AOI21_X1  g543(.A(G301), .B1(new_n609), .B2(new_n614), .ZN(new_n969));
  NOR2_X1   g544(.A1(G171), .A2(new_n557), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n897), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT77), .B1(new_n613), .B2(new_n532), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n608), .B(new_n531), .C1(new_n612), .C2(new_n548), .ZN(new_n973));
  OAI21_X1  g548(.A(G171), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n970), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n896), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n952), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n971), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n974), .A2(KEYINPUT107), .A3(new_n975), .A4(new_n896), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n953), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n982), .B2(KEYINPUT108), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n953), .C1(new_n980), .C2(new_n981), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n986), .B2(new_n963), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n962), .B1(new_n983), .B2(new_n985), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT43), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n990));
  INV_X1    g565(.A(new_n985), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n963), .A4(new_n978), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n952), .A2(new_n981), .A3(new_n980), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n953), .B2(new_n977), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n994), .B2(new_n962), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n992), .A2(new_n995), .A3(KEYINPUT43), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n987), .B2(new_n988), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n992), .A2(new_n995), .A3(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(G1996), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n805), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G160), .A2(G40), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n494), .B2(new_n499), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1006), .A2(new_n1007), .A3(KEYINPUT45), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n766), .A2(G2067), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n759), .A2(new_n771), .A3(new_n765), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1008), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(KEYINPUT109), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(KEYINPUT109), .B2(new_n1014), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT110), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n866), .B(new_n868), .Z(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n636), .B(G1986), .Z(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1008), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n945), .B(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n500), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1006), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1007), .A2(new_n1028), .A3(KEYINPUT45), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT111), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G40), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n930), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1007), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT116), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1007), .A2(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1037), .C1(new_n1007), .C2(new_n1038), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT117), .B(G1956), .Z(new_n1045));
  AND3_X1   g620(.A1(new_n1044), .A2(KEYINPUT118), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT118), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1023), .B(new_n1035), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1007), .A2(new_n1037), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT120), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n771), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1054));
  INV_X1    g629(.A(G1348), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n885), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1035), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1023), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1049), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1044), .A2(KEYINPUT118), .A3(new_n1045), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1023), .B1(new_n1068), .B2(new_n1035), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT61), .B1(new_n1069), .B2(new_n1049), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1062), .A2(new_n1071), .A3(new_n1048), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1052), .A2(new_n885), .A3(new_n1056), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT60), .B1(new_n1074), .B2(new_n1057), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT58), .B(G1341), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1051), .A2(new_n1076), .B1(new_n1032), .B2(G1996), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n577), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n885), .A2(KEYINPUT60), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1052), .A2(new_n1056), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1063), .B1(new_n1073), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1032), .A2(KEYINPUT112), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1027), .A2(new_n1031), .A3(new_n1089), .A4(new_n1029), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n443), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1961), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1054), .A2(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1096));
  NAND2_X1  g671(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT53), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1032), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT125), .B1(new_n1093), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1101), .A2(new_n1102), .A3(G171), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(G171), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1107));
  AOI211_X1 g682(.A(KEYINPUT125), .B(new_n1100), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT126), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1027), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1030), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1095), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT123), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1095), .A2(new_n1114), .A3(new_n1111), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1110), .B1(new_n1118), .B2(G301), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1106), .A2(new_n1109), .A3(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1103), .A2(G301), .ZN(new_n1121));
  AOI21_X1  g696(.A(G301), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1110), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(G303), .A2(G8), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT55), .Z(new_n1125));
  AOI21_X1  g700(.A(G1971), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1054), .A2(G2090), .ZN(new_n1127));
  OAI211_X1 g702(.A(G8), .B(new_n1125), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT113), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1044), .A2(G2090), .ZN(new_n1130));
  OAI21_X1  g705(.A(G8), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1125), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1030), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1037), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n840), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1053), .A2(new_n815), .A3(new_n1037), .A4(new_n1041), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1134), .B(G8), .C1(new_n1139), .C2(new_n557), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n557), .A2(G8), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1134), .B(new_n1142), .C1(new_n1139), .C2(G8), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1133), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(G1976), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G288), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(KEYINPUT114), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1050), .A2(G8), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(KEYINPUT114), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT52), .B1(G288), .B2(new_n1148), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT52), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT115), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(G305), .B2(G1981), .ZN(new_n1160));
  INV_X1    g735(.A(G1981), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n626), .A2(KEYINPUT115), .A3(new_n1161), .A4(new_n629), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n628), .B1(G86), .B2(new_n517), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1164), .B2(new_n624), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT49), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT49), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1168), .B(new_n1165), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1151), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1158), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1123), .A2(new_n1129), .A3(new_n1147), .A4(new_n1172), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1087), .A2(new_n1120), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT62), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1139), .A2(G8), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1176), .A2(KEYINPUT51), .A3(new_n1141), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1175), .A2(new_n1122), .A3(new_n1179), .ZN(new_n1180));
  OR3_X1    g755(.A1(new_n1176), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1133), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1129), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1172), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1148), .B(new_n846), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1151), .B1(new_n1185), .B2(new_n1163), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1176), .A2(G286), .ZN(new_n1187));
  OAI21_X1  g762(.A(G8), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1132), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1172), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1186), .B1(new_n1190), .B2(KEYINPUT63), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1184), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1021), .B1(new_n1174), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1008), .A2(new_n1004), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT46), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1008), .B1(new_n1013), .B2(new_n805), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(KEYINPUT127), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1196), .A2(KEYINPUT127), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT47), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1009), .A2(G1986), .A3(G290), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT48), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1200), .B1(new_n1019), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n866), .A2(new_n868), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1017), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1009), .B1(new_n1205), .B2(new_n1012), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1193), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g783(.A1(G227), .A2(new_n462), .ZN(new_n1210));
  AND3_X1   g784(.A1(new_n698), .A2(new_n742), .A3(new_n1210), .ZN(new_n1211));
  OAI211_X1 g785(.A(new_n1211), .B(new_n942), .C1(new_n1000), .C2(new_n1001), .ZN(G225));
  INV_X1    g786(.A(G225), .ZN(G308));
endmodule


