//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  AOI22_X1  g031(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT64), .Z(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  AND2_X1   g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n459), .A2(G137), .ZN(new_n464));
  AND2_X1   g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(G160));
  OAI21_X1  g043(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n469));
  INV_X1    g044(.A(G100), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(new_n463), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT66), .Z(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT65), .B1(new_n475), .B2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n463), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n472), .B(new_n481), .C1(G124), .C2(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n463), .B2(G114), .ZN(new_n487));
  NOR2_X1   g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n488), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n490), .A2(KEYINPUT67), .A3(G2104), .A4(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n489), .A2(new_n493), .B1(new_n484), .B2(G126), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT68), .A2(G138), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n463), .B(new_n495), .C1(new_n473), .C2(new_n474), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n459), .A2(new_n498), .A3(new_n463), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(G543), .B1(new_n504), .B2(KEYINPUT69), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT70), .A2(G88), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT70), .A2(G88), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n515), .A2(new_n516), .A3(new_n505), .A4(new_n508), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(KEYINPUT71), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT71), .B1(new_n517), .B2(new_n518), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n516), .A2(G89), .A3(new_n505), .A4(new_n508), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  AND3_X1   g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(new_n529), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n525), .A2(new_n526), .A3(new_n530), .A4(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n505), .A2(new_n508), .A3(G63), .A4(G651), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n538), .A2(new_n540), .A3(G51), .A4(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n534), .A2(new_n530), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n526), .B1(new_n544), .B2(new_n525), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n524), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n525), .A2(new_n530), .A3(new_n534), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n548), .A2(KEYINPUT74), .A3(new_n535), .A4(new_n542), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G168));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n505), .A2(new_n508), .A3(new_n538), .A4(new_n540), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n516), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n505), .A2(new_n508), .A3(G64), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n537), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(G171));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n552), .B1(new_n553), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n505), .A2(new_n508), .A3(G56), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n537), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n538), .A2(new_n540), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n509), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n516), .A2(KEYINPUT76), .A3(new_n505), .A4(new_n508), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(G91), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n538), .A2(new_n540), .A3(G53), .A4(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n509), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n577), .A2(new_n579), .A3(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n509), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n574), .A2(new_n507), .ZN(new_n589));
  AOI22_X1  g164(.A1(G651), .A2(new_n588), .B1(new_n589), .B2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n575), .A2(G87), .A3(new_n576), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G288));
  NAND3_X1  g167(.A1(new_n505), .A2(new_n508), .A3(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(KEYINPUT77), .A3(G651), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n575), .A2(G86), .A3(new_n576), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n509), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT78), .B(G85), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n516), .A2(new_n607), .A3(new_n505), .A4(new_n508), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n516), .A2(G47), .A3(G543), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n575), .A2(G92), .A3(new_n576), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n575), .A2(new_n617), .A3(G92), .A4(new_n576), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n509), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(new_n589), .B2(G54), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n616), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n614), .B1(new_n623), .B2(G868), .ZN(G321));
  NOR2_X1   g200(.A1(G299), .A2(G868), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g202(.A(new_n626), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n476), .A2(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n484), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n480), .B2(G135), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT80), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n654), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT81), .Z(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT17), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n666), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT82), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n668), .A3(new_n666), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n668), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n667), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(G2096), .Z(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(G2100), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(G2100), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT84), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n689), .B(new_n690), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n693), .B(new_n694), .C1(new_n688), .C2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  INV_X1    g276(.A(G1981), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n700), .A2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n590), .A2(new_n591), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n707), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n712), .B1(G1971), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n707), .A2(G6), .ZN(new_n716));
  INV_X1    g291(.A(G305), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT32), .B(G1981), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n715), .B(new_n720), .C1(G1971), .C2(new_n714), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n707), .A2(G24), .ZN(new_n724));
  INV_X1    g299(.A(new_n607), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n610), .B1(new_n552), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT79), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n727), .A2(new_n728), .B1(G651), .B2(new_n605), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n724), .B1(new_n729), .B2(new_n707), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT86), .Z(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(new_n697), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n697), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n484), .A2(G119), .ZN(new_n736));
  NOR2_X1   g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT85), .Z(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G131), .B2(new_n480), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n734), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XOR2_X1   g318(.A(new_n742), .B(new_n743), .Z(new_n744));
  NOR3_X1   g319(.A1(new_n732), .A2(new_n733), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n722), .A2(new_n723), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT36), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n734), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n734), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n616), .A2(new_n618), .A3(new_n622), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n707), .A2(G4), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n707), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  INV_X1    g336(.A(G299), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n707), .ZN(new_n763));
  INV_X1    g338(.A(G1956), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n752), .A2(new_n758), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n734), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n484), .A2(G128), .ZN(new_n769));
  NOR2_X1   g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n480), .B2(G140), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(new_n734), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n707), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n566), .B2(new_n707), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  AND2_X1   g353(.A1(KEYINPUT24), .A2(G34), .ZN(new_n779));
  NOR2_X1   g354(.A1(KEYINPUT24), .A2(G34), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n734), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT87), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n467), .B2(new_n734), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G11), .ZN(new_n788));
  INV_X1    g363(.A(G28), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n789), .B2(KEYINPUT30), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT30), .B2(new_n789), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n645), .B2(G29), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n775), .A2(new_n778), .A3(new_n785), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n734), .A2(G33), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n463), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n480), .B2(G139), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n734), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G2072), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n707), .A2(G5), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G171), .B2(new_n707), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT91), .B(G1961), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n734), .A2(G27), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G164), .B2(new_n734), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n734), .A2(G32), .ZN(new_n814));
  NAND3_X1  g389(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT26), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n484), .A2(G129), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n480), .B2(G141), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n734), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT27), .B(G1996), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n805), .A2(new_n809), .A3(new_n813), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT89), .B(G1966), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT88), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n707), .A2(G21), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G168), .B2(new_n707), .ZN(new_n828));
  AOI211_X1 g403(.A(new_n796), .B(new_n824), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n826), .B2(new_n828), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n747), .A2(new_n766), .A3(new_n830), .ZN(G311));
  OR3_X1    g406(.A1(new_n747), .A2(new_n766), .A3(new_n830), .ZN(G150));
  INV_X1    g407(.A(new_n565), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n552), .A2(new_n560), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n589), .A2(G43), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n505), .A2(new_n508), .A3(G67), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G651), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT92), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n516), .A2(G55), .A3(G543), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n516), .A2(G93), .A3(new_n505), .A4(new_n508), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n842), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n537), .B1(new_n837), .B2(new_n838), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT92), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n836), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n566), .A2(new_n841), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n623), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  INV_X1    g430(.A(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n849), .A2(new_n856), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n773), .B(new_n501), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n820), .ZN(new_n863));
  INV_X1    g438(.A(new_n803), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n862), .A2(new_n820), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n820), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n803), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n484), .A2(G130), .ZN(new_n870));
  NOR2_X1   g445(.A1(G106), .A2(G2105), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n480), .B2(G142), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n636), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n741), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n865), .A2(new_n878), .A3(new_n868), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n645), .B(new_n467), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n877), .A2(KEYINPUT93), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT93), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n869), .A2(new_n885), .A3(new_n876), .ZN(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n884), .A2(new_n886), .A3(new_n879), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT94), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n883), .A2(new_n888), .A3(KEYINPUT94), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT40), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(G395));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n896));
  OAI211_X1 g471(.A(G288), .B(new_n512), .C1(new_n521), .C2(new_n520), .ZN(new_n897));
  NAND2_X1  g472(.A1(G305), .A2(new_n729), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n601), .A2(new_n600), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT77), .B1(new_n595), .B2(G651), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n597), .B(new_n537), .C1(new_n593), .C2(new_n594), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(G290), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G303), .A2(new_n709), .ZN(new_n904));
  AND4_X1   g479(.A1(new_n897), .A2(new_n898), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n898), .A2(new_n903), .B1(new_n904), .B2(new_n897), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n898), .A2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n897), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n898), .A2(new_n903), .A3(new_n904), .A4(new_n897), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT97), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n911), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT98), .B(KEYINPUT42), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n913), .A2(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(KEYINPUT99), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n851), .B(new_n631), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT96), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n577), .A2(new_n579), .A3(KEYINPUT95), .A4(new_n583), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n921), .A2(new_n618), .A3(new_n616), .A4(new_n622), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT95), .ZN(new_n923));
  AND2_X1   g498(.A1(G299), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n753), .A2(new_n923), .A3(G299), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT41), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G299), .A2(new_n923), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n623), .A2(new_n928), .A3(new_n921), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n753), .A2(new_n923), .A3(G299), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n920), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n920), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n919), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n925), .A2(new_n926), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n919), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n917), .A2(KEYINPUT99), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n918), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n918), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(G868), .B2(new_n849), .ZN(G295));
  OAI21_X1  g519(.A(new_n943), .B1(G868), .B2(new_n849), .ZN(G331));
  NAND2_X1  g520(.A1(new_n848), .A2(new_n850), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n546), .A2(new_n549), .A3(G301), .ZN(new_n947));
  AOI21_X1  g522(.A(G301), .B1(new_n546), .B2(new_n549), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G168), .A2(G171), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n546), .A2(new_n549), .A3(G301), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n851), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n933), .B2(new_n935), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n937), .A2(new_n949), .A3(new_n952), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n955), .A2(new_n907), .A3(new_n912), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n956), .A3(KEYINPUT101), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n955), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n913), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n851), .B1(new_n950), .B2(new_n951), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n947), .A2(new_n948), .A3(new_n946), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT96), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n972), .B2(new_n934), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n955), .A2(new_n907), .A3(new_n912), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n958), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n955), .A2(KEYINPUT102), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n968), .A2(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n937), .A2(new_n949), .A3(new_n952), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n913), .ZN(new_n981));
  INV_X1    g556(.A(G37), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n975), .A2(new_n981), .A3(new_n960), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n959), .A2(KEYINPUT103), .A3(new_n960), .A4(new_n981), .ZN(new_n986));
  AND4_X1   g561(.A1(KEYINPUT104), .A2(new_n985), .A3(new_n986), .A4(KEYINPUT43), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n983), .B2(new_n984), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT104), .B1(new_n989), .B2(new_n986), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n966), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n996), .ZN(G397));
  NAND3_X1  g572(.A1(new_n462), .A2(new_n466), .A3(G40), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n501), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT106), .Z(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT107), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(KEYINPUT107), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n773), .B(G2067), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n820), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1003), .B(KEYINPUT106), .ZN(new_n1010));
  INV_X1    g585(.A(G1996), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT46), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT125), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT126), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT126), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(KEYINPUT47), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1007), .B1(new_n1011), .B2(new_n820), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1005), .A2(new_n1006), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1013), .A2(new_n820), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n741), .B(new_n743), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G290), .A2(G1986), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1010), .A2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1033));
  XNOR2_X1  g608(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G2067), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n773), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n741), .A2(new_n743), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n1027), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1030), .A2(new_n1034), .B1(new_n1038), .B2(new_n1028), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1023), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT47), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1384), .B1(new_n494), .B2(new_n500), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT108), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n998), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n784), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1054));
  AOI211_X1 g629(.A(KEYINPUT108), .B(G1384), .C1(new_n494), .C2(new_n500), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1002), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n998), .B1(new_n1046), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n825), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1049), .A2(new_n1061), .A3(new_n784), .A4(new_n1050), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1052), .A2(new_n1060), .A3(G168), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1051), .A2(KEYINPUT113), .B1(new_n1059), .B2(new_n825), .ZN(new_n1068));
  AOI21_X1  g643(.A(G168), .B1(new_n1068), .B2(new_n1062), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT51), .B1(new_n1063), .B2(G8), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1043), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1052), .A2(new_n1062), .A3(new_n1060), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G286), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1063), .A2(G8), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1064), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1077), .A3(KEYINPUT62), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1046), .A2(KEYINPUT45), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1971), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1046), .A2(KEYINPUT112), .A3(new_n1045), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT50), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n999), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1083), .B1(new_n1089), .B2(G2090), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G8), .ZN(new_n1091));
  NOR3_X1   g666(.A1(G166), .A2(KEYINPUT55), .A3(new_n1065), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(G303), .B2(G8), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1065), .B1(new_n1098), .B2(new_n999), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n899), .A2(new_n702), .A3(new_n902), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT109), .B(G86), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n516), .A2(new_n1101), .A3(new_n505), .A4(new_n508), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT110), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n600), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1102), .B2(new_n600), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(new_n902), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT49), .B(new_n1100), .C1(new_n1107), .C2(new_n702), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT49), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G305), .A2(G1981), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n702), .B1(new_n1106), .B2(new_n902), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1099), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1099), .A2(new_n1108), .A3(new_n1112), .A4(KEYINPUT111), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1049), .A2(new_n751), .A3(new_n1050), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1065), .B1(new_n1118), .B2(new_n1083), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1095), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1044), .A2(new_n999), .A3(new_n1048), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n709), .A2(G1976), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(G8), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n709), .B2(G1976), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(KEYINPUT52), .B2(new_n1123), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1097), .A2(new_n1117), .A3(new_n1120), .A4(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT50), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n999), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1049), .A2(new_n1132), .A3(new_n1050), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1961), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1081), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n1135), .B2(new_n812), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1056), .A2(KEYINPUT53), .A3(new_n812), .A4(new_n1058), .ZN(new_n1138));
  AOI21_X1  g713(.A(G301), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1072), .A2(new_n1078), .A3(new_n1128), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(G1976), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1117), .A2(new_n1141), .A3(new_n709), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1100), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1120), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1117), .A2(new_n1127), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1143), .A2(new_n1099), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(G286), .A2(new_n1065), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1073), .A2(KEYINPUT114), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT114), .B1(new_n1073), .B2(new_n1147), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT63), .B(new_n1120), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1119), .A2(new_n1095), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1145), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1117), .A3(new_n1127), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT115), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1150), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1149), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1073), .A2(KEYINPUT114), .A3(new_n1147), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n1128), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1140), .B(new_n1146), .C1(new_n1156), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1089), .A2(new_n764), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(G2072), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1135), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT119), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n577), .A2(new_n583), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT57), .B1(new_n1167), .B2(KEYINPUT116), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(G299), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1162), .A2(KEYINPUT119), .A3(new_n1165), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1133), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1132), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n757), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1098), .A2(new_n1035), .A3(new_n999), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n753), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1162), .A2(new_n1169), .A3(new_n1165), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1170), .A2(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1162), .A2(new_n1169), .A3(new_n1165), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT120), .B1(new_n1081), .B2(G1996), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1079), .A2(new_n1186), .A3(new_n1011), .A4(new_n1080), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT58), .B(G1341), .Z(new_n1188));
  NAND2_X1  g763(.A1(new_n1121), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n566), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1169), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1180), .B1(new_n1195), .B2(new_n1179), .ZN(new_n1196));
  OR2_X1    g771(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1191), .A2(new_n1193), .A3(new_n1197), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1184), .A2(new_n1194), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(KEYINPUT60), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1175), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n623), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n753), .A4(new_n1175), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1200), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1178), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT54), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1080), .A2(KEYINPUT53), .A3(new_n812), .ZN(new_n1209));
  OR2_X1    g784(.A1(new_n1079), .A2(KEYINPUT124), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1079), .A2(KEYINPUT124), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR4_X1   g787(.A1(new_n1134), .A2(new_n1136), .A3(new_n1212), .A4(G171), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1208), .B1(new_n1139), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1134), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1136), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1216), .A2(new_n1138), .A3(G301), .A4(new_n1217), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1134), .A2(new_n1136), .A3(new_n1212), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1218), .B(KEYINPUT54), .C1(new_n1219), .C2(G301), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1214), .A2(new_n1215), .A3(new_n1220), .A4(new_n1128), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1221), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1161), .B1(new_n1207), .B2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n729), .A2(new_n697), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1010), .B1(new_n1031), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1030), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1042), .B1(new_n1223), .B2(new_n1226), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g802(.A1(new_n891), .A2(new_n892), .ZN(new_n1229));
  AND4_X1   g803(.A1(new_n457), .A2(new_n682), .A3(new_n664), .A4(new_n683), .ZN(new_n1230));
  OAI21_X1  g804(.A(new_n1230), .B1(new_n704), .B2(new_n705), .ZN(new_n1231));
  AND2_X1   g805(.A1(new_n992), .A2(new_n993), .ZN(new_n1232));
  NOR3_X1   g806(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .ZN(G308));
  INV_X1    g807(.A(G229), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n891), .A2(new_n892), .ZN(new_n1235));
  NAND4_X1  g809(.A1(new_n1234), .A2(new_n1235), .A3(new_n994), .A4(new_n1230), .ZN(G225));
endmodule


