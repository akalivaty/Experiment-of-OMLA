//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(new_n203), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT65), .B(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n214), .B1(new_n215), .B2(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT67), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT69), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n207), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G50), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G50), .B2(new_n250), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT8), .A2(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n202), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G58), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n265), .B2(KEYINPUT8), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n208), .A2(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n260), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n258), .B1(new_n254), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g0070(.A(new_n270), .B(KEYINPUT9), .Z(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G222), .A2(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G223), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n253), .B1(G33), .B2(G41), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n276), .B(new_n277), .C1(G77), .C2(new_n272), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n277), .A2(new_n283), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G226), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n278), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(G200), .B2(new_n287), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT10), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n271), .A2(new_n290), .B1(KEYINPUT71), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n287), .A2(G179), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n287), .ZN(new_n297));
  INV_X1    g0097(.A(new_n270), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n285), .A2(G232), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n284), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  OAI211_X1 g0104(.A(G1), .B(G13), .C1(new_n304), .C2(new_n281), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT72), .B1(new_n304), .B2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(G223), .A2(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G226), .B2(new_n274), .ZN(new_n313));
  INV_X1    g0113(.A(G87), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n311), .A2(new_n313), .B1(new_n304), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n305), .B1(new_n315), .B2(KEYINPUT74), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT74), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n317), .B1(new_n304), .B2(new_n314), .C1(new_n311), .C2(new_n313), .ZN(new_n318));
  AOI211_X1 g0118(.A(G179), .B(new_n303), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(new_n277), .A3(new_n318), .ZN(new_n321));
  INV_X1    g0121(.A(new_n303), .ZN(new_n322));
  AOI21_X1  g0122(.A(G169), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT75), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n321), .A2(new_n325), .A3(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT75), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n303), .B1(new_n316), .B2(new_n318), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n327), .C1(G169), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT70), .B(G58), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n216), .B1(new_n221), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G20), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n259), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n272), .B2(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n308), .A2(G33), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n310), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n221), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n331), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n333), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n311), .A2(new_n337), .A3(new_n208), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n337), .B1(new_n311), .B2(new_n208), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n344), .B(KEYINPUT16), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n348), .A3(new_n254), .ZN(new_n349));
  INV_X1    g0149(.A(new_n255), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n266), .A2(new_n256), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n266), .A2(new_n256), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT73), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n352), .A2(new_n355), .B1(new_n251), .B2(new_n267), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n330), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT18), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n288), .B(new_n303), .C1(new_n316), .C2(new_n318), .ZN(new_n360));
  INV_X1    g0160(.A(G200), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n321), .B2(new_n322), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n363), .A2(KEYINPUT17), .A3(new_n356), .A4(new_n349), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n321), .A2(G190), .A3(new_n322), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n361), .B2(new_n328), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n357), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n330), .A2(new_n370), .A3(new_n357), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n359), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n221), .A2(G20), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n373), .A2(KEYINPUT12), .A3(new_n207), .A4(G13), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n255), .A2(G68), .A3(new_n256), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n250), .A2(G68), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n375), .C1(KEYINPUT12), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n259), .A2(G50), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n219), .B2(new_n268), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n254), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT11), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n380), .A2(new_n381), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G97), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n274), .A2(G232), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G226), .B2(G1698), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n387), .B1(new_n389), .B2(new_n340), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n277), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n305), .A2(G274), .A3(new_n283), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(G238), .B2(new_n285), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n391), .B2(new_n393), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n386), .B(G169), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n325), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n386), .B1(new_n398), .B2(G169), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n385), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(G200), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n384), .C1(new_n288), .C2(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT8), .B(G58), .Z(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT15), .B(G87), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n268), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n254), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n255), .A2(G77), .A3(new_n256), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(G77), .C2(new_n250), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n277), .A2(new_n283), .A3(new_n220), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n272), .A2(G238), .A3(G1698), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n272), .A2(G232), .A3(new_n274), .ZN(new_n414));
  INV_X1    g0214(.A(G107), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n413), .B(new_n414), .C1(new_n415), .C2(new_n272), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n392), .B(new_n412), .C1(new_n416), .C2(new_n277), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(G169), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n325), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n411), .B1(G190), .B2(new_n417), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n361), .B2(new_n417), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n301), .A2(new_n372), .A3(new_n404), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n207), .A2(G45), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT5), .B(G41), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n277), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  NAND2_X1  g0230(.A1(KEYINPUT5), .A2(G41), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n429), .A2(G264), .B1(new_n280), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G294), .ZN(new_n434));
  INV_X1    g0234(.A(G257), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G1698), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G250), .B2(G1698), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n434), .B1(new_n311), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n277), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G179), .ZN(new_n441));
  AOI21_X1  g0241(.A(G169), .B1(new_n433), .B2(new_n439), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n254), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT78), .B(G116), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n445), .A2(G20), .A3(new_n304), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n415), .A2(G20), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT23), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT22), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n208), .A2(new_n306), .A3(new_n309), .A4(new_n310), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G87), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n208), .A3(G87), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT83), .B1(new_n340), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n453), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT83), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n272), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n449), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT24), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n306), .A2(new_n309), .A3(new_n208), .A4(new_n310), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT22), .B1(new_n461), .B2(new_n314), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n454), .A3(new_n457), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n449), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n444), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  XOR2_X1   g0266(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n467));
  NOR2_X1   g0267(.A1(new_n250), .A2(G107), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n207), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n250), .A2(new_n470), .A3(new_n253), .A4(new_n252), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n415), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n443), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n463), .A2(new_n464), .A3(new_n449), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n464), .B1(new_n463), .B2(new_n449), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n254), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n473), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT85), .A3(new_n443), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n440), .A2(G200), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n288), .B2(new_n440), .ZN(new_n484));
  OR3_X1    g0284(.A1(new_n466), .A2(new_n484), .A3(new_n474), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n477), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  AOI21_X1  g0287(.A(G20), .B1(G33), .B2(G283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n304), .A2(G97), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n488), .A2(new_n489), .B1(new_n252), .B2(new_n253), .ZN(new_n490));
  INV_X1    g0290(.A(G116), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT78), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT78), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G116), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n494), .A3(G20), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT20), .B1(new_n490), .B2(new_n495), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n492), .A2(new_n494), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n471), .A2(new_n491), .B1(new_n499), .B2(new_n250), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n487), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n488), .A2(new_n489), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n495), .A2(new_n254), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n495), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n500), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(KEYINPUT82), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n325), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n429), .A2(G270), .B1(new_n280), .B2(new_n432), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n340), .A2(G303), .ZN(new_n512));
  AND2_X1   g0312(.A1(G264), .A2(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n306), .A2(new_n309), .A3(new_n310), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n309), .A2(new_n310), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n435), .A2(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(KEYINPUT81), .A3(new_n306), .A4(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT81), .ZN(new_n519));
  INV_X1    g0319(.A(new_n517), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n311), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n515), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n511), .B1(new_n522), .B2(new_n305), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n487), .B(new_n500), .C1(new_n505), .C2(new_n506), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT82), .B1(new_n507), .B2(new_n508), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(G200), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n288), .C2(new_n523), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n501), .A2(new_n509), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT21), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(G169), .A4(new_n523), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n296), .B1(new_n501), .B2(new_n509), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n535), .B2(new_n523), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n525), .B(new_n530), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n207), .A3(G45), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT77), .B1(new_n282), .B2(G1), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n305), .A2(G250), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n305), .A2(G274), .A3(new_n427), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n220), .A2(G1698), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G238), .B2(G1698), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n311), .A2(new_n545), .B1(new_n304), .B2(new_n445), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n543), .B1(new_n277), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G190), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  INV_X1    g0350(.A(G97), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n314), .A2(new_n551), .A3(new_n415), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n387), .A2(new_n208), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n268), .A2(KEYINPUT19), .A3(new_n551), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n203), .A2(new_n461), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n254), .B1(new_n251), .B2(new_n407), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n471), .A2(new_n314), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n547), .C2(new_n361), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT80), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n549), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n546), .A2(new_n277), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(new_n542), .A3(new_n541), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(KEYINPUT80), .A3(new_n557), .A4(new_n558), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n557), .B1(new_n471), .B2(new_n407), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n296), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n547), .A2(new_n325), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT79), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT79), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n547), .A2(new_n572), .A3(new_n325), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n220), .A2(G1698), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT4), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G283), .ZN(new_n580));
  AND2_X1   g0380(.A1(KEYINPUT4), .A2(G244), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n339), .A2(new_n310), .A3(new_n581), .A4(new_n274), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n277), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n429), .A2(G257), .B1(new_n280), .B2(new_n432), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n296), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n432), .A2(G274), .A3(new_n305), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n428), .A2(new_n427), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n305), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(new_n435), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  INV_X1    g0392(.A(new_n577), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n311), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(new_n580), .A3(new_n579), .A4(new_n582), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n591), .B1(new_n595), .B2(new_n277), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n325), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n259), .A2(G77), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT76), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n600), .A2(new_n551), .A3(G107), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n599), .B1(new_n208), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n415), .B1(new_n338), .B2(new_n341), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n254), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n251), .A2(new_n551), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n471), .B2(new_n551), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n587), .A2(new_n597), .A3(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n272), .A2(new_n337), .A3(G20), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT7), .B1(new_n340), .B2(new_n208), .ZN(new_n613));
  OAI21_X1  g0413(.A(G107), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(new_n599), .C1(new_n208), .C2(new_n603), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n608), .B1(new_n615), .B2(new_n254), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n586), .A2(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n596), .A2(G190), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n566), .A2(new_n575), .A3(new_n611), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n537), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n425), .A2(new_n486), .A3(new_n621), .ZN(G372));
  NOR2_X1   g0422(.A1(new_n481), .A2(new_n484), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n564), .A2(new_n557), .A3(new_n558), .A4(new_n548), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n619), .A2(new_n611), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n523), .B(G169), .C1(new_n526), .C2(new_n527), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT21), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n533), .B1(new_n524), .B2(new_n510), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n475), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n611), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n566), .A2(new_n575), .A3(new_n633), .A4(KEYINPUT26), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n625), .A2(new_n624), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n611), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n637), .A3(KEYINPUT86), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n561), .A2(new_n565), .B1(new_n569), .B2(new_n574), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n633), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n632), .A2(new_n624), .A3(new_n638), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n425), .A2(new_n642), .ZN(new_n643));
  AOI221_X4 g0443(.A(KEYINPUT18), .B1(new_n356), .B2(new_n349), .C1(new_n324), .C2(new_n329), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n370), .B1(new_n330), .B2(new_n357), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n403), .A2(new_n420), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n647), .A2(new_n401), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n364), .A2(new_n368), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n299), .B1(new_n650), .B2(new_n294), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n643), .A2(new_n651), .ZN(G369));
  INV_X1    g0452(.A(G13), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n653), .A2(G1), .A3(G20), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT87), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT27), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G213), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n481), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n486), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n475), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n662), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  INV_X1    g0468(.A(new_n662), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n630), .B(new_n530), .C1(new_n528), .C2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n525), .B1(new_n534), .B2(new_n536), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n531), .A3(new_n662), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n630), .A2(new_n662), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n486), .A2(new_n675), .B1(new_n665), .B2(new_n669), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n211), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G1), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n552), .A2(G116), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n681), .A2(new_n683), .B1(new_n217), .B2(new_n680), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n621), .A2(new_n486), .A3(new_n669), .ZN(new_n686));
  AOI21_X1  g0486(.A(G179), .B1(new_n433), .B2(new_n439), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n523), .A2(new_n586), .A3(new_n563), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n689));
  NOR2_X1   g0489(.A1(G250), .A2(G1698), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n435), .B2(G1698), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n306), .A3(new_n309), .A4(new_n310), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n305), .B1(new_n692), .B2(new_n434), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n589), .A2(G264), .A3(new_n305), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n588), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n325), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n547), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT89), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n523), .A4(new_n586), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n584), .B(new_n585), .C1(new_n305), .C2(new_n522), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n325), .B1(new_n429), .B2(G270), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n547), .A2(new_n439), .A3(new_n433), .A4(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n700), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n433), .A2(new_n702), .A3(new_n439), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n563), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n522), .A2(new_n305), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n707), .A4(new_n596), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n689), .A2(new_n699), .A3(new_n704), .A4(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT31), .B1(new_n709), .B2(new_n662), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n704), .A3(new_n688), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n669), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n710), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n668), .B1(new_n686), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n669), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT90), .B1(new_n642), .B2(new_n669), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT29), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n566), .A2(new_n575), .A3(new_n633), .A4(new_n635), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT26), .B1(new_n636), .B2(new_n611), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(new_n624), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n630), .A2(new_n477), .A3(new_n482), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n627), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n669), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT91), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT91), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n730), .A3(new_n669), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n720), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n716), .B1(new_n719), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n685), .B1(new_n734), .B2(G1), .ZN(G364));
  INV_X1    g0535(.A(new_n673), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n653), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n207), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n679), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n670), .A2(new_n672), .A3(new_n668), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n736), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n670), .A2(new_n672), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n208), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n272), .B1(new_n750), .B2(G303), .ZN(new_n751));
  NAND2_X1  g0551(.A1(G20), .A2(G179), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT95), .B1(new_n752), .B2(new_n361), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT95), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(G20), .A3(G179), .A4(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G190), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n751), .A2(KEYINPUT97), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(KEYINPUT97), .B2(new_n751), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n288), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n208), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n748), .A2(new_n288), .A3(new_n361), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n763), .A2(G294), .B1(new_n765), .B2(G329), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n748), .A2(new_n288), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n753), .A2(G190), .A3(new_n755), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n766), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT93), .ZN(new_n773));
  AOI21_X1  g0573(.A(G200), .B1(new_n752), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(KEYINPUT93), .A2(G20), .A3(G179), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n288), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n774), .A2(G190), .A3(new_n775), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n772), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n760), .A2(new_n771), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n765), .A2(G159), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(KEYINPUT32), .B1(G97), .B2(new_n763), .ZN(new_n782));
  INV_X1    g0582(.A(new_n757), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n782), .B1(KEYINPUT32), .B2(new_n781), .C1(new_n203), .C2(new_n783), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n272), .B1(new_n749), .B2(new_n314), .C1(new_n415), .C2(new_n768), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n201), .A2(new_n770), .B1(new_n777), .B2(new_n332), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n776), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT94), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT94), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G77), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n780), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n253), .B1(G20), .B2(new_n296), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n740), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n746), .A2(new_n795), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n678), .A2(new_n340), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n491), .B2(new_n678), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n248), .A2(G45), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT92), .Z(new_n802));
  NOR2_X1   g0602(.A1(new_n678), .A2(new_n576), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n217), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n797), .B1(new_n798), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n747), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n743), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  INV_X1    g0609(.A(new_n718), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n669), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n421), .A2(new_n662), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n662), .A2(new_n411), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n423), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n421), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n810), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n817), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n642), .A2(new_n819), .A3(new_n669), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n740), .B1(new_n821), .B2(new_n716), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n716), .B2(new_n821), .ZN(new_n823));
  INV_X1    g0623(.A(new_n770), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G150), .A2(new_n757), .B1(new_n824), .B2(G137), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  INV_X1    g0627(.A(G159), .ZN(new_n828));
  INV_X1    g0628(.A(new_n792), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n826), .B1(new_n827), .B2(new_n777), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT34), .Z(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n576), .B1(new_n832), .B2(new_n764), .ZN(new_n833));
  INV_X1    g0633(.A(new_n768), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n763), .A2(new_n265), .B1(new_n834), .B2(G68), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n201), .B2(new_n749), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n831), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G303), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n838), .A2(new_n770), .B1(new_n777), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n750), .A2(G107), .B1(new_n834), .B2(G87), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n757), .A2(G283), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n763), .A2(G97), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n272), .B1(new_n765), .B2(G311), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n840), .B(new_n845), .C1(new_n499), .C2(new_n792), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n795), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n795), .A2(new_n744), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n741), .B1(new_n219), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n745), .C2(new_n819), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n823), .A2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(KEYINPUT103), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n649), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n364), .A2(new_n368), .A3(KEYINPUT103), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(new_n359), .A3(new_n371), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n660), .B1(new_n349), .B2(new_n356), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n357), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n858), .B2(new_n363), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n358), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n358), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n348), .A2(new_n254), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT7), .B1(new_n576), .B2(G20), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(G68), .A3(new_n345), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT16), .B1(new_n869), .B2(new_n344), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n356), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n660), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n357), .B2(new_n367), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n869), .A2(new_n344), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n331), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n254), .A3(new_n348), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n324), .A2(new_n329), .B1(new_n877), .B2(new_n356), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n873), .ZN(new_n880));
  AOI221_X4 g0680(.A(new_n866), .B1(new_n879), .B2(new_n863), .C1(new_n372), .C2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT40), .B1(new_n865), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n669), .A2(new_n384), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n401), .A2(new_n403), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n404), .A2(new_n883), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n817), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n619), .A2(new_n611), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n630), .A2(new_n639), .A3(new_n530), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n477), .A2(new_n482), .A3(new_n485), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n889), .A2(new_n890), .A3(new_n662), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n709), .A2(new_n662), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n712), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  INV_X1    g0697(.A(new_n894), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n710), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n686), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n887), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n882), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n886), .A2(new_n885), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n819), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n686), .A2(new_n899), .A3(new_n897), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT105), .B1(new_n891), .B2(new_n895), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n873), .B1(new_n646), .B2(new_n369), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n879), .A2(new_n863), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n866), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n372), .A2(new_n880), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n879), .A2(new_n863), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n910), .A2(KEYINPUT101), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT101), .B1(new_n910), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n907), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n425), .B1(new_n896), .B2(new_n900), .ZN(new_n920));
  OAI21_X1  g0720(.A(G330), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  INV_X1    g0722(.A(new_n903), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n820), .A2(new_n813), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT100), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT100), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n820), .A2(new_n926), .A3(new_n813), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT101), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n911), .B2(new_n912), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n881), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n910), .A2(KEYINPUT101), .A3(new_n913), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n646), .A2(new_n872), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT39), .B1(new_n881), .B2(new_n930), .ZN(new_n936));
  XNOR2_X1  g0736(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n855), .A2(new_n856), .B1(new_n861), .B2(new_n863), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n913), .B(new_n937), .C1(new_n938), .C2(KEYINPUT38), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n401), .A2(new_n662), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT102), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n935), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n810), .A2(new_n720), .A3(new_n811), .ZN(new_n946));
  INV_X1    g0746(.A(new_n731), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n730), .B1(new_n727), .B2(new_n669), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT29), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n949), .A3(new_n425), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n651), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n945), .B(new_n951), .Z(new_n952));
  OR2_X1    g0752(.A1(new_n922), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n922), .A2(new_n952), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(new_n207), .C2(new_n737), .ZN(new_n955));
  INV_X1    g0755(.A(new_n603), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n491), .B(new_n215), .C1(new_n956), .C2(KEYINPUT35), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(KEYINPUT35), .B2(new_n956), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT36), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n221), .A2(new_n332), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n960), .A2(new_n219), .A3(new_n217), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n203), .A2(G50), .ZN(new_n962));
  OAI211_X1 g0762(.A(G1), .B(new_n653), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT99), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n955), .A2(new_n965), .ZN(G367));
  INV_X1    g0766(.A(new_n803), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n798), .B1(new_n211), .B2(new_n407), .C1(new_n967), .C2(new_n239), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n740), .ZN(new_n969));
  INV_X1    g0769(.A(G150), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n827), .A2(new_n770), .B1(new_n777), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n340), .B1(new_n765), .B2(G137), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n332), .B2(new_n749), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n762), .A2(new_n203), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n768), .A2(new_n219), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n828), .B2(new_n783), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n971), .B(new_n977), .C1(G50), .C2(new_n792), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n792), .A2(G283), .ZN(new_n979));
  INV_X1    g0779(.A(new_n777), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G311), .A2(new_n824), .B1(new_n980), .B2(G303), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n839), .B2(new_n783), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n750), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n834), .A2(G97), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n415), .C2(new_n762), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n749), .A2(new_n445), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n311), .B1(new_n986), .B2(new_n764), .C1(new_n987), .C2(KEYINPUT46), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n982), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n978), .B1(new_n979), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT47), .Z(new_n991));
  AOI21_X1  g0791(.A(new_n969), .B1(new_n991), .B2(new_n795), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n557), .A2(new_n558), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n662), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n624), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT106), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n625), .A2(new_n994), .A3(new_n624), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT107), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n746), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n992), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n679), .B(new_n1006), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n671), .A2(new_n669), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n664), .A2(new_n666), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n486), .A2(new_n675), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n673), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n736), .A3(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n716), .B(new_n1014), .C1(new_n719), .C2(new_n732), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT111), .B1(new_n667), .B2(new_n673), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n888), .B1(new_n616), .B2(new_n669), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n633), .A2(new_n662), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1008), .A2(new_n890), .B1(new_n475), .B2(new_n662), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1019), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n667), .A2(KEYINPUT111), .A3(new_n673), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT44), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1016), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT44), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1028), .B(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1016), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n1026), .A4(new_n1025), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1015), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(KEYINPUT112), .B(new_n1007), .C1(new_n1035), .C2(new_n733), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT112), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n733), .B1(new_n1038), .B2(new_n1014), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1007), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1036), .A2(new_n1041), .A3(new_n738), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1010), .A2(new_n1023), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT42), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1017), .B1(new_n477), .B2(new_n482), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n669), .B1(new_n1045), .B2(new_n633), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1001), .B(KEYINPUT43), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT109), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1047), .A2(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(KEYINPUT109), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n674), .A2(new_n1023), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT108), .Z(new_n1055));
  AND3_X1   g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1005), .B1(new_n1042), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1061), .B(new_n1005), .C1(new_n1042), .C2(new_n1058), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1060), .A2(new_n1062), .ZN(G387));
  AOI22_X1  g0863(.A1(G311), .A2(new_n757), .B1(new_n980), .B2(G317), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n778), .B2(new_n770), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G303), .B2(new_n792), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT115), .Z(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT48), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1066), .B(KEYINPUT115), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n763), .A2(G283), .B1(new_n750), .B2(G294), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT116), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1068), .A2(new_n1071), .A3(KEYINPUT49), .A4(new_n1072), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n311), .B1(new_n764), .B2(new_n769), .C1(new_n445), .C2(new_n768), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G77), .A2(new_n750), .B1(new_n765), .B2(G150), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT114), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n407), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n763), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1083), .A2(new_n576), .A3(new_n984), .A4(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G159), .A2(new_n824), .B1(new_n789), .B2(G68), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n201), .B2(new_n777), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1082), .A2(KEYINPUT114), .B1(new_n783), .B2(new_n267), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n795), .B1(new_n1081), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT117), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n664), .A2(new_n666), .A3(new_n746), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n236), .A2(new_n282), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1094), .A2(new_n803), .B1(new_n683), .B2(new_n799), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n405), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(G50), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT50), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n282), .B1(new_n203), .B2(new_n219), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n683), .B(new_n1099), .C1(new_n1098), .C2(new_n1097), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1095), .A2(new_n1100), .B1(G107), .B2(new_n211), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n741), .B1(new_n1101), .B2(new_n798), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1080), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1090), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n796), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1093), .A2(new_n1102), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT117), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1103), .A2(new_n1112), .B1(new_n739), .B2(new_n1014), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n733), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n679), .A3(new_n1015), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(G393));
  AOI21_X1  g0916(.A(new_n1038), .B1(new_n734), .B2(new_n1014), .ZN(new_n1117));
  OR3_X1    g0917(.A1(new_n1117), .A2(new_n1035), .A3(new_n680), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1038), .A2(new_n739), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n244), .A2(new_n967), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n798), .B1(new_n551), .B2(new_n211), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n740), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n762), .A2(new_n445), .B1(new_n749), .B2(new_n767), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n340), .B1(new_n764), .B2(new_n778), .C1(new_n415), .C2(new_n768), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G303), .C2(new_n757), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n986), .A2(new_n770), .B1(new_n777), .B2(new_n772), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT52), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(new_n839), .C2(new_n776), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT119), .Z(new_n1129));
  AOI22_X1  g0929(.A1(new_n757), .A2(G50), .B1(new_n763), .B2(G77), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n829), .B2(new_n1096), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT118), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n970), .A2(new_n770), .B1(new_n777), .B2(new_n828), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT51), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n314), .A2(new_n768), .B1(new_n749), .B2(new_n221), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n311), .B(new_n1135), .C1(G143), .C2(new_n765), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1129), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1122), .B1(new_n1138), .B2(new_n795), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1002), .B2(new_n1019), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1118), .A2(new_n1119), .A3(new_n1140), .ZN(G390));
  AOI21_X1  g0941(.A(new_n668), .B1(new_n906), .B2(new_n905), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n887), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n927), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n926), .B1(new_n820), .B2(new_n813), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n903), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n940), .B1(new_n1147), .B2(new_n942), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n729), .A2(new_n731), .A3(new_n813), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n816), .A3(new_n903), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n913), .B1(new_n938), .B2(KEYINPUT38), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1151), .A2(new_n942), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1144), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n716), .A2(new_n817), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n903), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n928), .A2(new_n943), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1153), .B(new_n1157), .C1(new_n1158), .C2(new_n940), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n425), .A2(new_n1142), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n950), .A2(new_n651), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1143), .B1(new_n903), .B2(new_n1156), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1149), .A2(new_n816), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1142), .A2(new_n819), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n1157), .C1(new_n1166), .C2(new_n903), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1162), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1160), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1155), .A2(new_n1168), .A3(new_n1159), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n679), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1155), .A2(new_n1159), .A3(new_n739), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n848), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n740), .B1(new_n1174), .B2(new_n266), .ZN(new_n1175));
  INV_X1    g0975(.A(G125), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n272), .B1(new_n764), .B2(new_n1176), .C1(new_n762), .C2(new_n828), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n750), .A2(G150), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT53), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(G50), .C2(new_n834), .ZN(new_n1180));
  INV_X1    g0980(.A(G128), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1181), .A2(new_n770), .B1(new_n777), .B2(new_n832), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G137), .B2(new_n757), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT54), .B(G143), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1180), .B(new_n1183), .C1(new_n829), .C2(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n762), .A2(new_n219), .B1(new_n768), .B2(new_n203), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n340), .B1(new_n764), .B2(new_n839), .C1(new_n314), .C2(new_n749), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(G107), .C2(new_n757), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G283), .A2(new_n824), .B1(new_n980), .B2(G116), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n551), .C2(new_n829), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT120), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n796), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1185), .A2(KEYINPUT120), .A3(new_n1190), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1175), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n940), .B2(new_n745), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1172), .A2(new_n1173), .A3(new_n1195), .ZN(G378));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n301), .A2(new_n298), .A3(new_n872), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n294), .B(new_n300), .C1(new_n270), .C2(new_n660), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT122), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1197), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n918), .B2(G330), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n907), .A2(KEYINPUT40), .A3(new_n1151), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n901), .B1(new_n931), .B2(new_n932), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G330), .B(new_n1206), .C1(new_n1207), .C2(KEYINPUT40), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1203), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1209), .A2(KEYINPUT122), .A3(new_n1200), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n945), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n918), .A2(G330), .A3(new_n1204), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n945), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1212), .A2(new_n1213), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1162), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1171), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(KEYINPUT123), .B(new_n945), .C1(new_n1205), .C2(new_n1211), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n680), .B1(new_n1225), .B2(new_n1220), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1218), .A2(new_n739), .A3(new_n1221), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1201), .A2(new_n744), .A3(new_n1203), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n749), .A2(new_n219), .B1(new_n764), .B2(new_n767), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n311), .A2(new_n281), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n768), .A2(new_n332), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT121), .Z(new_n1234));
  AOI21_X1  g1034(.A(new_n974), .B1(G97), .B2(new_n757), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n824), .A2(G116), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G107), .A2(new_n980), .B1(new_n789), .B2(new_n1084), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT58), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1231), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n762), .A2(new_n970), .B1(new_n749), .B2(new_n1184), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G128), .A2(new_n980), .B1(new_n789), .B2(G137), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1176), .B2(new_n770), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(G132), .C2(new_n757), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n834), .A2(G159), .ZN(new_n1249));
  AOI211_X1 g1049(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1242), .B1(new_n1239), .B2(new_n1238), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n795), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n741), .B1(new_n201), .B2(new_n848), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1229), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1228), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1227), .A2(new_n1259), .ZN(G375));
  OAI21_X1  g1060(.A(new_n740), .B1(new_n1174), .B2(G68), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n749), .A2(new_n828), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1232), .B(new_n1262), .C1(G50), .C2(new_n763), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n311), .B1(new_n765), .B2(G128), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1184), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n757), .A2(new_n1265), .B1(new_n789), .B2(G150), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G132), .A2(new_n824), .B1(new_n980), .B2(G137), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n829), .A2(new_n415), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n272), .B(new_n975), .C1(G303), .C2(new_n765), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n980), .A2(G283), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n763), .A2(new_n1084), .B1(new_n750), .B2(G97), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n499), .A2(new_n757), .B1(new_n824), .B2(G294), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1268), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1261), .B1(new_n1275), .B2(new_n795), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n903), .B2(new_n745), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n738), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1168), .A2(new_n1040), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1162), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(G381));
  INV_X1    g1083(.A(G378), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(G390), .A2(G384), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1284), .A2(new_n1282), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  OR3_X1    g1087(.A1(G375), .A2(new_n1287), .A3(G387), .ZN(G407));
  AOI21_X1  g1088(.A(new_n1258), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n661), .A3(new_n1284), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G407), .A2(G213), .A3(new_n1290), .ZN(G409));
  NAND4_X1  g1091(.A1(new_n1218), .A2(new_n1220), .A3(new_n1007), .A4(new_n1221), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1256), .B1(new_n1293), .B2(new_n739), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G378), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1289), .B2(G378), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n658), .A2(G343), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G384), .B(KEYINPUT124), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1278), .A2(KEYINPUT60), .A3(new_n1162), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n679), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1169), .A2(KEYINPUT60), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1300), .B1(new_n1301), .B2(new_n1281), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1298), .B1(new_n1302), .B2(new_n1279), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1299), .A2(new_n679), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1281), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1279), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  OR2_X1    g1106(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1303), .A2(new_n1308), .ZN(new_n1309));
  NOR4_X1   g1109(.A1(new_n1296), .A2(KEYINPUT62), .A3(new_n1297), .A4(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1227), .A2(G378), .A3(new_n1259), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1284), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1297), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1297), .A2(G2897), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1303), .A2(new_n1308), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1303), .B2(new_n1308), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1311), .B1(new_n1315), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1309), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1315), .B2(new_n1323), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1310), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1059), .B(G390), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n808), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1285), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1042), .A2(new_n1058), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1004), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1061), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1333));
  INV_X1    g1133(.A(G390), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1328), .B1(new_n1059), .B2(G390), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1335), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1336), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1329), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT125), .ZN(new_n1341));
  AOI211_X1 g1141(.A(new_n1297), .B(new_n1309), .C1(new_n1312), .C2(new_n1314), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1341), .B1(new_n1342), .B2(KEYINPUT63), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1297), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(new_n1345), .A3(new_n1323), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1346), .A2(KEYINPUT125), .A3(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1343), .A2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1323), .ZN(new_n1350));
  OAI22_X1  g1150(.A1(new_n1296), .A2(new_n1297), .B1(new_n1319), .B2(new_n1318), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT61), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1350), .A2(new_n1340), .A3(new_n1351), .A4(new_n1352), .ZN(new_n1353));
  OAI22_X1  g1153(.A1(new_n1325), .A2(new_n1340), .B1(new_n1349), .B2(new_n1353), .ZN(G405));
  NAND2_X1  g1154(.A1(G375), .A2(new_n1284), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1312), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1340), .A2(new_n1357), .ZN(new_n1358));
  OAI211_X1 g1158(.A(new_n1356), .B(new_n1329), .C1(new_n1339), .C2(new_n1338), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1358), .A2(new_n1359), .A3(new_n1323), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1323), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1360), .A2(new_n1361), .ZN(G402));
endmodule


