//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT98), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n202), .B(KEYINPUT98), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT100), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n210), .A2(KEYINPUT99), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(KEYINPUT99), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(new_n206), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G8gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT97), .B(G29gat), .Z(new_n224));
  OAI221_X1 g023(.A(new_n221), .B1(KEYINPUT15), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n213), .A2(new_n230), .A3(new_n217), .A4(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT101), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT102), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n213), .A2(new_n217), .A3(new_n227), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n229), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n234), .B(KEYINPUT13), .Z(new_n241));
  NAND3_X1  g040(.A1(new_n218), .A2(KEYINPUT102), .A3(new_n228), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n229), .A2(new_n234), .A3(new_n232), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT101), .A3(new_n235), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  INV_X1    g046(.A(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT11), .B(G169gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT12), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n237), .A2(new_n243), .A3(new_n245), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT89), .B(KEYINPUT0), .Z(new_n258));
  XNOR2_X1  g057(.A(G1gat), .B(G29gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G57gat), .B(G85gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT80), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(G155gat), .A3(G162gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G141gat), .B(G148gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n264), .B(new_n269), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT82), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(new_n265), .A3(new_n270), .ZN(new_n279));
  INV_X1    g078(.A(G148gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G141gat), .ZN(new_n281));
  INV_X1    g080(.A(G141gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G148gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n263), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT82), .A3(new_n269), .ZN(new_n286));
  OR2_X1    g085(.A1(KEYINPUT84), .A2(G155gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT84), .A2(G155gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(G162gat), .A3(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n289), .A2(KEYINPUT2), .B1(new_n264), .B2(new_n265), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n284), .B(KEYINPUT83), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n277), .A2(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G113gat), .B(G120gat), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT69), .ZN(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G127gat), .B(G134gat), .Z(new_n299));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n293), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT1), .B1(new_n295), .B2(KEYINPUT70), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n298), .A2(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT4), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n286), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n290), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT87), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n292), .A2(KEYINPUT87), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n303), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT4), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n275), .A2(new_n276), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT82), .B1(new_n285), .B2(new_n269), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n308), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT85), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n307), .A2(new_n321), .A3(new_n316), .A4(new_n308), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n303), .B1(new_n309), .B2(KEYINPUT3), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n323), .A2(KEYINPUT86), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT86), .B1(new_n323), .B2(new_n324), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n306), .B(new_n315), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n327), .A2(KEYINPUT5), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n292), .A2(new_n303), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n305), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT88), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT88), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n334), .B(new_n329), .C1(new_n305), .C2(new_n331), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(KEYINPUT5), .A3(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT4), .B(new_n303), .C1(new_n311), .C2(new_n312), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n304), .A2(new_n314), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n328), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n324), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n323), .A2(KEYINPUT86), .A3(new_n324), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n336), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n262), .B1(new_n330), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT6), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n343), .A2(new_n344), .B1(new_n314), .B2(new_n313), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT5), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n328), .A4(new_n306), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n333), .A2(KEYINPUT5), .A3(new_n335), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n325), .A2(new_n326), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n339), .ZN(new_n354));
  INV_X1    g153(.A(new_n262), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n347), .A2(new_n348), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(KEYINPUT6), .B(new_n262), .C1(new_n330), .C2(new_n346), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT66), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT66), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n364));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT24), .ZN(new_n370));
  INV_X1    g169(.A(G183gat), .ZN(new_n371));
  INV_X1    g170(.A(G190gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n372), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G176gat), .ZN(new_n377));
  AND2_X1   g176(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n379));
  OAI211_X1 g178(.A(KEYINPUT23), .B(new_n377), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT67), .B(G190gat), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n373), .B(new_n374), .C1(new_n384), .C2(G183gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n367), .A2(KEYINPUT23), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(KEYINPUT25), .A3(new_n386), .A4(new_n369), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n368), .A2(new_n389), .A3(new_n365), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n367), .A2(KEYINPUT26), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(new_n391), .C1(new_n371), .C2(new_n372), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT67), .B(G190gat), .Z(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT27), .B(G183gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n394), .A2(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n394), .A2(new_n396), .A3(new_n397), .A4(new_n395), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n388), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n402), .A2(new_n403), .B1(G226gat), .B2(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n394), .A2(new_n395), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n398), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n387), .A2(new_n383), .B1(new_n407), .B2(new_n393), .ZN(new_n408));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G211gat), .ZN(new_n411));
  INV_X1    g210(.A(G218gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414));
  NAND2_X1  g213(.A1(G211gat), .A2(G218gat), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT77), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT76), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G197gat), .B(G204gat), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT22), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n418), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n427), .B(KEYINPUT77), .C1(new_n416), .C2(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n404), .A2(new_n410), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n409), .B1(new_n408), .B2(KEYINPUT29), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT78), .ZN(new_n435));
  INV_X1    g234(.A(new_n410), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT78), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(new_n409), .C1(new_n408), .C2(KEYINPUT29), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n439), .B2(new_n432), .ZN(new_n440));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n360), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OR3_X1    g245(.A1(new_n440), .A2(new_n360), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n443), .ZN(new_n448));
  OAI211_X1 g247(.A(KEYINPUT79), .B(new_n360), .C1(new_n440), .C2(new_n443), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n359), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n323), .A2(new_n403), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n431), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n309), .A2(new_n310), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n292), .A2(KEYINPUT87), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n429), .A2(new_n403), .A3(new_n430), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n429), .A2(KEYINPUT90), .A3(new_n403), .A4(new_n430), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n316), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n457), .B(new_n458), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n454), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n316), .B1(new_n459), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n309), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT29), .B1(new_n320), .B2(new_n322), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n469), .B(new_n454), .C1(new_n470), .C2(new_n432), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT93), .B(G22gat), .C1(new_n465), .C2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G78gat), .B(G106gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G50gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n464), .B1(new_n470), .B2(new_n432), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n453), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT92), .B(G22gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n471), .ZN(new_n481));
  INV_X1    g280(.A(G22gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n479), .B2(new_n471), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(KEYINPUT93), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT94), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n476), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n483), .B2(KEYINPUT93), .ZN(new_n487));
  OAI21_X1  g286(.A(G22gat), .B1(new_n465), .B2(new_n472), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n487), .A2(new_n490), .A3(new_n491), .A4(new_n481), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n465), .A2(new_n472), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(new_n480), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n485), .A2(new_n492), .B1(new_n494), .B2(new_n486), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n452), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n303), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n402), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n408), .A2(new_n303), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(G227gat), .A2(G233gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G43gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n388), .A2(new_n303), .A3(new_n401), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n303), .B1(new_n388), .B2(new_n401), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n501), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT71), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n516), .B(new_n501), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT72), .B1(new_n518), .B2(KEYINPUT32), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n523));
  AOI211_X1 g322(.A(new_n522), .B(new_n523), .C1(new_n515), .C2(new_n517), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n520), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT73), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(new_n520), .C1(new_n521), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n516), .B1(new_n500), .B2(new_n501), .ZN(new_n530));
  INV_X1    g329(.A(new_n517), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT32), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n511), .A2(new_n519), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n507), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g335(.A(new_n534), .B(new_n506), .C1(new_n526), .C2(new_n528), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT75), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(KEYINPUT36), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n532), .A2(new_n522), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n518), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n527), .B1(new_n544), .B2(new_n520), .ZN(new_n545));
  INV_X1    g344(.A(new_n528), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n535), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n506), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n529), .A2(new_n535), .A3(new_n507), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n496), .B1(new_n539), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT95), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n485), .A2(new_n492), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n494), .A2(new_n486), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT38), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n443), .B1(new_n440), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n435), .A2(new_n431), .A3(new_n438), .A4(new_n436), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n432), .B1(new_n404), .B2(new_n410), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(KEYINPUT37), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n443), .B(new_n560), .C1(new_n440), .C2(KEYINPUT37), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n556), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n439), .A2(new_n432), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n433), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n556), .B1(new_n440), .B2(KEYINPUT37), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n557), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n357), .A2(new_n568), .A3(new_n358), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n327), .A2(new_n329), .ZN(new_n570));
  OR3_X1    g369(.A1(new_n305), .A2(new_n329), .A3(new_n331), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT39), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT39), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n327), .A2(new_n573), .A3(new_n329), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n355), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n572), .A2(KEYINPUT40), .A3(new_n355), .A4(new_n574), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n347), .A4(new_n450), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n555), .A2(new_n569), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n541), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(new_n536), .B2(new_n537), .ZN(new_n582));
  INV_X1    g381(.A(new_n538), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n548), .A2(new_n549), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n586), .A3(new_n496), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n552), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n548), .A2(new_n549), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n555), .ZN(new_n590));
  AOI211_X1 g389(.A(KEYINPUT96), .B(new_n450), .C1(new_n357), .C2(new_n358), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT35), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n548), .A2(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n257), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT104), .B(KEYINPUT7), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n602), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G99gat), .B(G106gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n230), .A2(new_n231), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n611), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n228), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT105), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n618), .A3(new_n615), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n600), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n619), .A3(new_n600), .ZN(new_n622));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  AND3_X1   g424(.A1(new_n621), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n621), .B2(new_n622), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g429(.A1(G71gat), .A2(G78gat), .ZN(new_n631));
  OR2_X1    g430(.A1(G71gat), .A2(G78gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT9), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G57gat), .B(G64gat), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT103), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(KEYINPUT9), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n631), .A3(new_n632), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n213), .B(new_n217), .C1(new_n630), .C2(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(G183gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(G183gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n640), .A2(new_n630), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(new_n411), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G127gat), .B(G155gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(G231gat), .A2(G233gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n651), .B1(new_n647), .B2(new_n648), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n653), .B2(new_n658), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n629), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n611), .B(new_n640), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(KEYINPUT10), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n614), .A2(KEYINPUT10), .A3(new_n637), .A4(new_n639), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G230gat), .A2(G233gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n669), .B2(KEYINPUT106), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n667), .B(new_n675), .C1(KEYINPUT106), .C2(new_n669), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT107), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n661), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n598), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n359), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n209), .ZN(G1324gat));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n451), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n207), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n689), .B2(new_n691), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n687), .A2(KEYINPUT108), .A3(KEYINPUT42), .A4(new_n688), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(G1325gat));
  INV_X1    g495(.A(G15gat), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n582), .A2(new_n584), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n582), .B2(new_n584), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n684), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n684), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n589), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n697), .B2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n684), .A2(new_n555), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NAND2_X1  g507(.A1(new_n659), .A2(new_n660), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n677), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n598), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n629), .ZN(new_n712));
  INV_X1    g511(.A(new_n359), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n224), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(KEYINPUT45), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n585), .A2(KEYINPUT109), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n357), .A2(new_n358), .A3(new_n568), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n495), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n719), .A2(new_n579), .B1(new_n495), .B2(new_n452), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n582), .A2(new_n584), .A3(new_n698), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n717), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n597), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT44), .B1(new_n723), .B2(new_n629), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n628), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n588), .B2(new_n597), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n256), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT110), .B1(new_n253), .B2(new_n255), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(new_n734), .A3(new_n710), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n359), .ZN(new_n736));
  OAI22_X1  g535(.A1(new_n715), .A2(new_n716), .B1(new_n224), .B2(new_n736), .ZN(G1328gat));
  NAND3_X1  g536(.A1(new_n712), .A2(new_n223), .A3(new_n450), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n735), .B2(new_n451), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(G1329gat));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n712), .A2(new_n743), .A3(new_n589), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  OAI21_X1  g544(.A(G43gat), .B1(new_n735), .B2(new_n701), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1330gat));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n711), .A2(new_n495), .A3(new_n629), .ZN(new_n751));
  INV_X1    g550(.A(G50gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n735), .A2(new_n752), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n750), .B(new_n753), .C1(new_n754), .C2(new_n555), .ZN(new_n755));
  INV_X1    g554(.A(new_n753), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n735), .A2(new_n752), .A3(new_n555), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT48), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(G1331gat));
  AND2_X1   g558(.A1(new_n723), .A2(new_n661), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n734), .A2(new_n678), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n713), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g564(.A1(new_n762), .A2(new_n451), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n762), .B2(new_n701), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(new_n589), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G71gat), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g573(.A1(new_n763), .A2(new_n495), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g575(.A1(new_n734), .A2(new_n709), .A3(new_n678), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n729), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n778), .A2(new_n605), .A3(new_n359), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n734), .A2(new_n709), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n580), .A2(new_n496), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n699), .A2(new_n700), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n594), .A2(new_n595), .A3(new_n591), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n595), .B1(new_n594), .B2(new_n591), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n629), .B(new_n780), .C1(new_n782), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n723), .A2(new_n788), .A3(new_n629), .A4(new_n780), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n677), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(new_n359), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n779), .B1(new_n605), .B2(new_n791), .ZN(G1336gat));
  OAI21_X1  g591(.A(G92gat), .B1(new_n778), .B2(new_n451), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n790), .A2(new_n451), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(G92gat), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n796), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n793), .B(new_n798), .C1(new_n794), .C2(G92gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1337gat));
  XNOR2_X1  g599(.A(KEYINPUT112), .B(G99gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n778), .B2(new_n701), .ZN(new_n802));
  INV_X1    g601(.A(new_n589), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n803), .A2(new_n801), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n790), .B2(new_n804), .ZN(G1338gat));
  OAI21_X1  g604(.A(new_n629), .B1(new_n782), .B2(new_n785), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n725), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n585), .A2(new_n586), .A3(new_n496), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n586), .B1(new_n585), .B2(new_n496), .ZN(new_n809));
  INV_X1    g608(.A(new_n580), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n726), .B1(new_n811), .B2(new_n785), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n807), .A2(new_n812), .A3(new_n495), .A4(new_n777), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n790), .A2(G106gat), .A3(new_n555), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT53), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND4_X1   g615(.A1(new_n495), .A2(new_n787), .A3(new_n677), .A4(new_n789), .ZN(new_n817));
  INV_X1    g616(.A(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT53), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n729), .A2(new_n821), .A3(new_n495), .A4(new_n777), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n822), .A3(G106gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n819), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n819), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n816), .B1(new_n825), .B2(new_n826), .ZN(G1339gat));
  INV_X1    g626(.A(new_n709), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n663), .A2(new_n664), .A3(new_n668), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n667), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n665), .A2(new_n666), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n673), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n673), .A4(new_n832), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n676), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n731), .B2(new_n732), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n240), .A2(new_n242), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n840), .A2(new_n241), .B1(new_n234), .B2(new_n233), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n251), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n255), .A3(new_n677), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n629), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n255), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n837), .A2(new_n628), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n828), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n661), .A2(new_n678), .A3(new_n733), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n495), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n359), .A2(new_n450), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n589), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n257), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n733), .A2(G113gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(G1340gat));
  INV_X1    g653(.A(new_n851), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n677), .ZN(new_n856));
  INV_X1    g655(.A(G120gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(KEYINPUT116), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(KEYINPUT116), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n856), .B2(new_n858), .ZN(G1341gat));
  NAND2_X1  g660(.A1(new_n855), .A2(new_n709), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g662(.A1(new_n855), .A2(new_n629), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(G134gat), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT56), .B1(new_n864), .B2(G134gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n843), .B1(new_n837), .B2(new_n257), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n846), .B1(new_n628), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n848), .B1(new_n871), .B2(new_n709), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(new_n495), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n555), .B1(new_n847), .B2(new_n848), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n869), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n701), .A2(new_n850), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n734), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(KEYINPUT117), .A3(G141gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n876), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n256), .A2(new_n282), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n881), .B2(new_n880), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT117), .B1(new_n877), .B2(G141gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n878), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n884), .A2(KEYINPUT58), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n875), .A2(new_n876), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n282), .B1(new_n890), .B2(new_n256), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n886), .A2(new_n887), .B1(new_n888), .B2(new_n891), .ZN(G1344gat));
  NOR3_X1   g691(.A1(new_n879), .A2(G148gat), .A3(new_n678), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT119), .Z(new_n894));
  AND3_X1   g693(.A1(new_n680), .A2(new_n257), .A3(new_n682), .ZN(new_n895));
  OR3_X1    g694(.A1(new_n837), .A2(new_n628), .A3(KEYINPUT120), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT120), .B1(new_n837), .B2(new_n628), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n255), .A3(new_n842), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n870), .A2(new_n628), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n709), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n869), .B(new_n495), .C1(new_n895), .C2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n901), .B(new_n677), .C1(new_n869), .C2(new_n874), .ZN(new_n902));
  INV_X1    g701(.A(new_n876), .ZN(new_n903));
  OAI21_X1  g702(.A(G148gat), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(KEYINPUT59), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n280), .C1(new_n890), .C2(new_n677), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(G1345gat));
  AND2_X1   g706(.A1(new_n287), .A2(new_n288), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n889), .B2(new_n828), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n874), .A2(new_n709), .A3(new_n876), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(G1346gat));
  NOR2_X1   g712(.A1(new_n879), .A2(new_n628), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(G162gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n889), .A2(new_n628), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n713), .A2(new_n451), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n589), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n849), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n734), .C1(new_n379), .C2(new_n378), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(KEYINPUT122), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n920), .A2(KEYINPUT122), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n849), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n257), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n922), .A2(new_n926), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n377), .A3(new_n677), .ZN(new_n928));
  OAI21_X1  g727(.A(G176gat), .B1(new_n925), .B2(new_n678), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT123), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n921), .A2(new_n395), .A3(new_n709), .ZN(new_n932));
  OAI21_X1  g731(.A(G183gat), .B1(new_n925), .B2(new_n828), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n921), .A2(new_n394), .A3(new_n629), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n925), .A2(new_n628), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(G190gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n937), .B2(G190gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n701), .A2(new_n918), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n874), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  XOR2_X1   g744(.A(KEYINPUT124), .B(G197gat), .Z(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n734), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n901), .B1(new_n869), .B2(new_n874), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(new_n257), .A3(new_n942), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n950), .B2(new_n947), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT125), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n944), .A2(G204gat), .A3(new_n678), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n902), .B2(new_n942), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n945), .A2(new_n411), .A3(new_n709), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n949), .A2(new_n942), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n709), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  NOR2_X1   g761(.A1(new_n628), .A2(new_n412), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n629), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT126), .B1(new_n965), .B2(new_n412), .ZN(new_n966));
  OAI211_X1 g765(.A(KEYINPUT126), .B(new_n412), .C1(new_n944), .C2(new_n628), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n964), .B(KEYINPUT127), .C1(new_n966), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1355gat));
endmodule


