//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  AND4_X1   g008(.A1(new_n202), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n204), .B2(new_n206), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n202), .B1(new_n211), .B2(new_n208), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n208), .ZN(new_n214));
  XNOR2_X1  g013(.A(G113gat), .B(G120gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n209), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n207), .A2(KEYINPUT69), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT27), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n225), .B2(KEYINPUT27), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n221), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n233), .B(new_n221), .C1(new_n227), .C2(new_n230), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT28), .A3(new_n229), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT68), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239));
  INV_X1    g038(.A(new_n237), .ZN(new_n240));
  AOI211_X1 g039(.A(new_n239), .B(new_n240), .C1(new_n232), .C2(new_n234), .ZN(new_n241));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT26), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n242), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n238), .A2(new_n241), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n225), .A2(new_n229), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT24), .A3(new_n242), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n242), .A2(KEYINPUT24), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n244), .A2(KEYINPUT23), .ZN(new_n255));
  OR3_X1    g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n243), .B1(new_n244), .B2(KEYINPUT23), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n255), .B(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n260), .B(new_n262), .C1(new_n259), .C2(new_n253), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n263), .B2(new_n254), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n220), .B1(new_n249), .B2(new_n264), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n229), .B(new_n228), .C1(new_n236), .C2(new_n222), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n233), .B1(new_n266), .B2(new_n221), .ZN(new_n267));
  INV_X1    g066(.A(new_n234), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n237), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n239), .ZN(new_n270));
  INV_X1    g069(.A(new_n248), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n235), .A2(KEYINPUT68), .A3(new_n237), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n220), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n254), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n257), .B2(new_n256), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n265), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G227gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n278), .A2(new_n280), .B1(new_n281), .B2(KEYINPUT33), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G99gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT71), .B(G71gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n274), .B1(new_n273), .B2(new_n276), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT33), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n290), .A2(new_n279), .B1(KEYINPUT32), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  INV_X1    g092(.A(new_n286), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI221_X1 g094(.A(KEYINPUT32), .B1(new_n291), .B2(new_n286), .C1(new_n290), .C2(new_n279), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n287), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n287), .A2(new_n295), .A3(new_n296), .A4(KEYINPUT73), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n278), .A2(new_n280), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n302), .A2(KEYINPUT34), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(KEYINPUT34), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(KEYINPUT74), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n305), .A2(new_n296), .A3(new_n287), .A4(new_n295), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n301), .A2(KEYINPUT75), .A3(new_n309), .ZN(new_n314));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(G211gat), .ZN(new_n316));
  INV_X1    g115(.A(G218gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(KEYINPUT22), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G141gat), .B(G148gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n324), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n324), .B(new_n328), .C1(new_n322), .C2(KEYINPUT2), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n321), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT86), .ZN(new_n335));
  INV_X1    g134(.A(new_n332), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT85), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT3), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT85), .B1(new_n321), .B2(KEYINPUT29), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G228gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n335), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n344), .B(KEYINPUT87), .Z(new_n345));
  AOI211_X1 g144(.A(new_n342), .B(new_n343), .C1(new_n337), .C2(new_n332), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n334), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G22gat), .B(G50gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n349), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G85gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n211), .A2(new_n202), .A3(new_n208), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT1), .B1(new_n207), .B2(KEYINPUT69), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n215), .A2(new_n216), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n208), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n213), .A2(KEYINPUT80), .A3(new_n219), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n336), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n336), .A2(new_n219), .A3(new_n213), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n363), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n333), .B1(new_n372), .B2(new_n373), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n379), .A2(new_n347), .B1(KEYINPUT4), .B2(new_n376), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n363), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n333), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n368), .A2(new_n371), .A3(new_n364), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT80), .B1(new_n213), .B2(new_n219), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n347), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n376), .A2(KEYINPUT4), .ZN(new_n389));
  AND4_X1   g188(.A1(new_n378), .A2(new_n388), .A3(new_n389), .A4(new_n383), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT5), .B(new_n377), .C1(new_n384), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n381), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n388), .B(new_n392), .C1(KEYINPUT4), .C2(new_n376), .ZN(new_n393));
  OR3_X1    g192(.A1(new_n393), .A2(KEYINPUT5), .A3(new_n363), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n361), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n391), .A2(new_n361), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G226gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(new_n343), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n273), .B2(new_n276), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n273), .A2(new_n276), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n408), .B2(new_n404), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n321), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n405), .A2(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n403), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n273), .B2(new_n276), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n412), .B1(new_n403), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n411), .B1(new_n414), .B2(KEYINPUT78), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n410), .B1(new_n415), .B2(new_n321), .ZN(new_n416));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417));
  INV_X1    g216(.A(G92gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT79), .B(G64gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT30), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n411), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n409), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n321), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n421), .B1(new_n428), .B2(new_n410), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n431), .A3(new_n422), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n401), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT83), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n414), .A2(new_n427), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n436), .B1(new_n426), .B2(new_n427), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n421), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n416), .A2(new_n422), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT30), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n432), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n401), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT35), .B1(new_n357), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n391), .A2(new_n361), .A3(new_n394), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(new_n395), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n448), .B2(new_n397), .ZN(new_n449));
  NOR4_X1   g248(.A1(new_n447), .A2(new_n395), .A3(KEYINPUT90), .A4(KEYINPUT6), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n400), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n441), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT35), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n297), .A2(new_n303), .A3(new_n304), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n313), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n355), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(new_n441), .A3(KEYINPUT92), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n455), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n421), .B1(new_n437), .B2(KEYINPUT37), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n414), .A2(new_n427), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT37), .B(new_n463), .C1(new_n426), .C2(new_n427), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT38), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n439), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT91), .B1(new_n451), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n466), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n422), .B1(new_n416), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n429), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n399), .A2(KEYINPUT90), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n446), .A3(new_n397), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n472), .A2(new_n473), .A3(new_n400), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n416), .A2(new_n470), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT38), .B1(new_n462), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n374), .A2(new_n376), .A3(new_n363), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  OR3_X1    g281(.A1(new_n481), .A2(KEYINPUT88), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n393), .A2(new_n363), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT88), .B1(new_n481), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n393), .A2(new_n482), .A3(new_n363), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n361), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n489), .A2(KEYINPUT89), .A3(KEYINPUT40), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n490), .A2(new_n493), .A3(new_n395), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(KEYINPUT40), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n432), .A3(new_n440), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(new_n356), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n312), .A2(KEYINPUT36), .A3(new_n313), .A4(new_n314), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n457), .A2(KEYINPUT77), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT77), .B1(new_n457), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n444), .A2(new_n355), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n498), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n461), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G43gat), .B(G50gat), .Z(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n510), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n519), .A2(new_n512), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G1gat), .B2(new_n527), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(G8gat), .Z(new_n531));
  XOR2_X1   g330(.A(new_n526), .B(new_n531), .Z(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT13), .Z(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n531), .B1(new_n525), .B2(new_n522), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n526), .B(KEYINPUT17), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n531), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT97), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT18), .B1(new_n540), .B2(KEYINPUT98), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT98), .A2(KEYINPUT18), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n539), .B1(KEYINPUT97), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n535), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G169gat), .B(G197gat), .Z(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT93), .B(KEYINPUT11), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT94), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT12), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n535), .B(new_n553), .C1(new_n541), .C2(new_n543), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n552), .A2(KEYINPUT99), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT99), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT100), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(G71gat), .B2(G78gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT101), .ZN(new_n561));
  INV_X1    g360(.A(G64gat), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n562), .A2(G57gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(G57gat), .ZN(new_n564));
  AND2_X1   g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n563), .A2(new_n564), .B1(KEYINPUT9), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n565), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OR3_X1    g368(.A1(new_n566), .A2(G71gat), .A3(G78gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n531), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n225), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n572), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G211gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n578), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(new_n418), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT102), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT102), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT7), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n591), .A2(KEYINPUT103), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(KEYINPUT103), .C1(new_n587), .C2(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n585), .B2(new_n418), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n537), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n526), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G134gat), .B(G162gat), .Z(new_n606));
  AOI21_X1  g405(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n605), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n598), .B(new_n571), .Z(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n598), .A2(new_n571), .A3(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G230gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n343), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n620), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n617), .B1(new_n613), .B2(new_n614), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND4_X1   g429(.A1(new_n583), .A2(new_n584), .A3(new_n610), .A4(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n507), .A2(new_n558), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n401), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G1gat), .ZN(G1324gat));
  INV_X1    g434(.A(new_n441), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n637), .A2(KEYINPUT105), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(KEYINPUT105), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G8gat), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  NAND3_X1  g441(.A1(new_n637), .A2(KEYINPUT42), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n641), .B(new_n643), .C1(new_n646), .C2(new_n647), .ZN(G1325gat));
  INV_X1    g447(.A(new_n457), .ZN(new_n649));
  AOI21_X1  g448(.A(G15gat), .B1(new_n632), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n504), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n651), .A2(G15gat), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n632), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT106), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n632), .A2(new_n355), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G22gat), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  AOI21_X1  g457(.A(new_n610), .B1(new_n461), .B2(new_n506), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n584), .A2(new_n583), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n630), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n659), .A2(new_n558), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n513), .A3(new_n633), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n609), .B(KEYINPUT108), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n461), .B2(new_n506), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n668), .B2(new_n659), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n552), .A2(new_n554), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n662), .ZN(new_n674));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674), .B2(new_n401), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n665), .A2(new_n675), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n663), .A2(new_n514), .A3(new_n636), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT46), .Z(new_n678));
  OAI21_X1  g477(.A(G36gat), .B1(new_n674), .B2(new_n441), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1329gat));
  OAI21_X1  g479(.A(G43gat), .B1(new_n674), .B2(new_n504), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT47), .B1(new_n681), .B2(KEYINPUT109), .ZN(new_n682));
  INV_X1    g481(.A(G43gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n663), .A2(new_n683), .A3(new_n649), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n682), .B(new_n685), .ZN(G1330gat));
  INV_X1    g485(.A(KEYINPUT48), .ZN(new_n687));
  INV_X1    g486(.A(G50gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n663), .A2(new_n688), .A3(new_n355), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT110), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n672), .A2(new_n673), .A3(new_n355), .A4(new_n662), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n691), .A2(G50gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n687), .B1(new_n691), .B2(G50gat), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n694), .A2(KEYINPUT111), .A3(new_n689), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT111), .B1(new_n694), .B2(new_n689), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(G1331gat));
  AND2_X1   g496(.A1(new_n584), .A2(new_n583), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n673), .A2(new_n630), .ZN(new_n699));
  AND4_X1   g498(.A1(new_n507), .A2(new_n698), .A3(new_n610), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n633), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n636), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT49), .B(G64gat), .Z(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(G1333gat));
  AOI21_X1  g505(.A(G71gat), .B1(new_n700), .B2(new_n649), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n651), .A2(G71gat), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n700), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1334gat));
  NAND2_X1  g510(.A1(new_n700), .A2(new_n355), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT113), .B(G78gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1335gat));
  NOR3_X1   g513(.A1(new_n698), .A2(new_n673), .A3(new_n630), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n672), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n585), .A3(new_n401), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n698), .A2(new_n673), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT114), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n507), .A2(new_n718), .A3(new_n609), .A4(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n719), .A2(KEYINPUT114), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n722), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n659), .A2(new_n724), .A3(new_n718), .A4(new_n720), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(new_n629), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(new_n401), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n717), .B1(new_n727), .B2(new_n585), .ZN(G1336gat));
  NAND3_X1  g527(.A1(new_n672), .A2(new_n636), .A3(new_n715), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(G92gat), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n726), .A2(G92gat), .A3(new_n441), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT52), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT115), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n733), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n734), .A2(G92gat), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n731), .A2(KEYINPUT52), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(G1337gat));
  OAI21_X1  g537(.A(G99gat), .B1(new_n716), .B2(new_n504), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n457), .A2(G99gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n726), .B2(new_n740), .ZN(G1338gat));
  AOI21_X1  g540(.A(new_n668), .B1(new_n507), .B2(new_n609), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n355), .B(new_n715), .C1(new_n742), .C2(new_n670), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G106gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n356), .A2(G106gat), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n723), .A2(new_n629), .A3(new_n725), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT53), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n672), .A2(KEYINPUT116), .A3(new_n355), .A4(new_n715), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(G106gat), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n748), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT117), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n748), .B(new_n757), .C1(new_n752), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1339gat));
  NAND3_X1  g558(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n619), .A2(KEYINPUT54), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n624), .B1(new_n627), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n763), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n766), .A2(new_n625), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n673), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n538), .A2(new_n533), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n532), .A2(new_n534), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n550), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n554), .A2(new_n629), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT118), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n554), .A2(new_n629), .A3(new_n775), .A4(new_n772), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n769), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT119), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n769), .A2(new_n779), .A3(new_n774), .A4(new_n776), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n666), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n554), .A2(new_n772), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n667), .A2(new_n768), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n698), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR4_X1   g583(.A1(new_n660), .A2(new_n673), .A3(new_n609), .A4(new_n629), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n357), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n633), .A3(new_n787), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n788), .A2(KEYINPUT120), .A3(new_n636), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT120), .B1(new_n788), .B2(new_n636), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n789), .A2(new_n205), .A3(new_n673), .A4(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n786), .A2(new_n458), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n636), .A2(new_n401), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G113gat), .B1(new_n794), .B2(new_n557), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(G1340gat));
  NAND4_X1  g595(.A1(new_n789), .A2(new_n203), .A3(new_n629), .A4(new_n790), .ZN(new_n797));
  OAI21_X1  g596(.A(G120gat), .B1(new_n794), .B2(new_n630), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1341gat));
  INV_X1    g598(.A(G127gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n794), .A2(new_n800), .A3(new_n660), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n788), .A2(new_n636), .A3(new_n660), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n800), .ZN(G1342gat));
  NAND3_X1  g602(.A1(new_n792), .A2(new_n609), .A3(new_n793), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n805), .A3(G134gat), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n805), .B1(new_n804), .B2(G134gat), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n788), .A2(G134gat), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n636), .A2(new_n610), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n809), .A2(KEYINPUT56), .A3(new_n810), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n807), .A2(new_n808), .B1(new_n811), .B2(new_n812), .ZN(G1343gat));
  NAND3_X1  g612(.A1(new_n786), .A2(new_n633), .A3(new_n355), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n814), .A2(new_n636), .A3(new_n651), .ZN(new_n815));
  INV_X1    g614(.A(G141gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n558), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n355), .B1(new_n784), .B2(new_n785), .ZN(new_n819));
  XNOR2_X1  g618(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n673), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n631), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n783), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n768), .B1(new_n555), .B2(new_n556), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n609), .B1(new_n825), .B2(new_n773), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n660), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n356), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n819), .A2(new_n821), .B1(new_n828), .B2(KEYINPUT57), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n504), .A2(new_n793), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n829), .A2(new_n557), .A3(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n817), .B(new_n818), .C1(new_n816), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n673), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n814), .A2(G141gat), .A3(new_n636), .A4(new_n651), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n834), .A2(G141gat), .B1(new_n835), .B2(new_n558), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n818), .ZN(G1344gat));
  INV_X1    g636(.A(G148gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n815), .A2(new_n838), .A3(new_n629), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840));
  INV_X1    g639(.A(new_n830), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n355), .B(new_n820), .C1(new_n784), .C2(new_n785), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n631), .A2(new_n557), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n768), .A2(new_n609), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT123), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n768), .A2(new_n847), .A3(new_n609), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n846), .A2(new_n782), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n660), .B1(new_n849), .B2(new_n826), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n851), .B2(new_n355), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n629), .B(new_n841), .C1(new_n843), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n838), .B1(new_n853), .B2(KEYINPUT124), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n843), .A2(new_n852), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n629), .A4(new_n841), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n840), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g657(.A(KEYINPUT59), .B(new_n838), .C1(new_n833), .C2(new_n629), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n839), .B1(new_n858), .B2(new_n859), .ZN(G1345gat));
  AOI21_X1  g659(.A(G155gat), .B1(new_n815), .B2(new_n698), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n660), .A2(new_n326), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n833), .B2(new_n862), .ZN(G1346gat));
  INV_X1    g662(.A(new_n814), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(new_n327), .A3(new_n504), .A4(new_n810), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n829), .A2(new_n666), .A3(new_n830), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n327), .ZN(G1347gat));
  NOR2_X1   g666(.A1(new_n441), .A2(new_n633), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n786), .A2(new_n458), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869), .B2(new_n557), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n786), .A2(new_n787), .A3(new_n868), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n822), .A2(G169gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1348gat));
  INV_X1    g672(.A(G176gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n871), .B2(new_n630), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT125), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n869), .A2(new_n874), .A3(new_n630), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1349gat));
  OAI21_X1  g677(.A(G183gat), .B1(new_n869), .B2(new_n660), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n698), .A2(new_n236), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n871), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g681(.A(G190gat), .B1(new_n869), .B2(new_n610), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT126), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n886), .B(G190gat), .C1(new_n869), .C2(new_n610), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n885), .B1(new_n884), .B2(new_n887), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n667), .A2(new_n229), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n888), .A2(new_n889), .B1(new_n871), .B2(new_n890), .ZN(G1351gat));
  AND2_X1   g690(.A1(new_n504), .A2(new_n868), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n855), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G197gat), .B1(new_n893), .B2(new_n557), .ZN(new_n894));
  INV_X1    g693(.A(new_n819), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n892), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n822), .A2(G197gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1352gat));
  OR3_X1    g697(.A1(new_n896), .A2(G204gat), .A3(new_n630), .ZN(new_n899));
  XOR2_X1   g698(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n855), .A2(new_n629), .A3(new_n892), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G204gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n901), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(G1353gat));
  INV_X1    g705(.A(new_n896), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n316), .A3(new_n698), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n855), .A2(new_n698), .A3(new_n892), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT63), .B1(new_n909), .B2(G211gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1354gat));
  OAI21_X1  g711(.A(G218gat), .B1(new_n893), .B2(new_n610), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n907), .A2(new_n317), .A3(new_n667), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1355gat));
endmodule


