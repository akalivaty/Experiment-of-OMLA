

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  NOR2_X2 U322 ( .A1(n579), .A2(n485), .ZN(n486) );
  XNOR2_X1 U323 ( .A(n412), .B(n411), .ZN(n525) );
  XNOR2_X1 U324 ( .A(n302), .B(n301), .ZN(n306) );
  XNOR2_X1 U325 ( .A(n324), .B(n422), .ZN(n529) );
  XOR2_X1 U326 ( .A(G36GAT), .B(n397), .Z(n290) );
  XOR2_X1 U327 ( .A(KEYINPUT62), .B(n581), .Z(n291) );
  NOR2_X1 U328 ( .A1(n558), .A2(n403), .ZN(n404) );
  INV_X1 U329 ( .A(KEYINPUT48), .ZN(n411) );
  XNOR2_X1 U330 ( .A(n294), .B(KEYINPUT33), .ZN(n295) );
  XNOR2_X1 U331 ( .A(n374), .B(G50GAT), .ZN(n375) );
  INV_X1 U332 ( .A(n413), .ZN(n299) );
  XNOR2_X1 U333 ( .A(n334), .B(n295), .ZN(n297) );
  XNOR2_X1 U334 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U335 ( .A(n300), .B(n299), .ZN(n301) );
  AND2_X1 U336 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U337 ( .A(KEYINPUT124), .B(n566), .ZN(n578) );
  NOR2_X1 U338 ( .A1(n529), .A2(n448), .ZN(n557) );
  XNOR2_X1 U339 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U340 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  XOR2_X1 U341 ( .A(G78GAT), .B(G204GAT), .Z(n293) );
  XNOR2_X1 U342 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n334) );
  AND2_X1 U344 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  INV_X1 U345 ( .A(KEYINPUT32), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .Z(n345) );
  XNOR2_X1 U348 ( .A(n345), .B(KEYINPUT31), .ZN(n300) );
  XNOR2_X1 U349 ( .A(G176GAT), .B(G92GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n298), .B(G64GAT), .ZN(n413) );
  XNOR2_X1 U351 ( .A(G120GAT), .B(G148GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n303), .B(G57GAT), .ZN(n425) );
  XNOR2_X1 U353 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n304), .B(KEYINPUT74), .ZN(n396) );
  XNOR2_X1 U355 ( .A(n425), .B(n396), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n572) );
  XOR2_X1 U357 ( .A(n572), .B(KEYINPUT41), .Z(n544) );
  XOR2_X1 U358 ( .A(n544), .B(KEYINPUT109), .Z(n531) );
  XOR2_X1 U359 ( .A(G176GAT), .B(G71GAT), .Z(n308) );
  XNOR2_X1 U360 ( .A(KEYINPUT20), .B(KEYINPUT65), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n319) );
  XOR2_X1 U362 ( .A(G134GAT), .B(G190GAT), .Z(n311) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n309), .B(KEYINPUT85), .ZN(n426) );
  XNOR2_X1 U365 ( .A(G99GAT), .B(n426), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G127GAT), .Z(n313) );
  NAND2_X1 U368 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U370 ( .A(n315), .B(n314), .Z(n317) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(G15GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U374 ( .A(KEYINPUT17), .B(G183GAT), .Z(n321) );
  XNOR2_X1 U375 ( .A(G169GAT), .B(KEYINPUT86), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U377 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n422) );
  XOR2_X1 U379 ( .A(KEYINPUT3), .B(G162GAT), .Z(n326) );
  XNOR2_X1 U380 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U382 ( .A(G141GAT), .B(n327), .Z(n433) );
  XOR2_X1 U383 ( .A(G148GAT), .B(KEYINPUT88), .Z(n329) );
  XNOR2_X1 U384 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U386 ( .A(G22GAT), .B(n330), .Z(n332) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U389 ( .A(n333), .B(KEYINPUT91), .Z(n339) );
  XOR2_X1 U390 ( .A(n334), .B(KEYINPUT22), .Z(n336) );
  XOR2_X1 U391 ( .A(G50GAT), .B(KEYINPUT77), .Z(n356) );
  XNOR2_X1 U392 ( .A(n356), .B(KEYINPUT23), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n337), .B(KEYINPUT87), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n433), .B(n340), .ZN(n344) );
  XOR2_X1 U397 ( .A(KEYINPUT21), .B(G218GAT), .Z(n342) );
  XNOR2_X1 U398 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(G197GAT), .B(n343), .Z(n417) );
  XOR2_X1 U401 ( .A(n344), .B(n417), .Z(n463) );
  XOR2_X1 U402 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n347) );
  XOR2_X1 U403 ( .A(G29GAT), .B(G134GAT), .Z(n441) );
  XNOR2_X1 U404 ( .A(n441), .B(n345), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U406 ( .A(n348), .B(KEYINPUT79), .Z(n353) );
  XOR2_X1 U407 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n350) );
  XNOR2_X1 U408 ( .A(KEYINPUT80), .B(KEYINPUT78), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U410 ( .A(G218GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U412 ( .A(G36GAT), .B(G190GAT), .Z(n416) );
  XOR2_X1 U413 ( .A(n354), .B(n416), .Z(n358) );
  XNOR2_X1 U414 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n355), .B(KEYINPUT7), .ZN(n378) );
  XNOR2_X1 U416 ( .A(n378), .B(n356), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U418 ( .A(G92GAT), .B(G106GAT), .Z(n360) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U421 ( .A(G162GAT), .B(n361), .Z(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n558) );
  XOR2_X1 U423 ( .A(KEYINPUT72), .B(KEYINPUT69), .Z(n365) );
  XNOR2_X1 U424 ( .A(KEYINPUT70), .B(KEYINPUT30), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n382) );
  XNOR2_X1 U426 ( .A(G15GAT), .B(G22GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n366), .B(G8GAT), .ZN(n397) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n290), .B(n367), .ZN(n376) );
  XOR2_X1 U430 ( .A(G141GAT), .B(G113GAT), .Z(n369) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(G29GAT), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U433 ( .A(KEYINPUT68), .B(KEYINPUT73), .Z(n371) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(G1GAT), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U436 ( .A(n373), .B(n372), .Z(n374) );
  XOR2_X1 U437 ( .A(n377), .B(KEYINPUT29), .Z(n380) );
  XNOR2_X1 U438 ( .A(n378), .B(KEYINPUT71), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n567) );
  NAND2_X1 U441 ( .A1(n567), .A2(n544), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n383), .B(KEYINPUT46), .ZN(n402) );
  XOR2_X1 U443 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n385) );
  XNOR2_X1 U444 ( .A(KEYINPUT84), .B(KEYINPUT14), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n392) );
  XOR2_X1 U446 ( .A(G64GAT), .B(G57GAT), .Z(n387) );
  XNOR2_X1 U447 ( .A(G155GAT), .B(G211GAT), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U449 ( .A(G1GAT), .B(G127GAT), .Z(n440) );
  XOR2_X1 U450 ( .A(n388), .B(n440), .Z(n390) );
  XNOR2_X1 U451 ( .A(G183GAT), .B(G78GAT), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n401) );
  XOR2_X1 U454 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n394) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(n395), .B(KEYINPUT81), .Z(n399) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n484) );
  NAND2_X1 U461 ( .A1(n402), .A2(n484), .ZN(n403) );
  XNOR2_X1 U462 ( .A(KEYINPUT47), .B(n404), .ZN(n410) );
  INV_X1 U463 ( .A(n558), .ZN(n469) );
  XNOR2_X1 U464 ( .A(n469), .B(KEYINPUT36), .ZN(n579) );
  NOR2_X1 U465 ( .A1(n484), .A2(n579), .ZN(n406) );
  XNOR2_X1 U466 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n408) );
  NOR2_X1 U468 ( .A1(n567), .A2(n572), .ZN(n407) );
  NAND2_X1 U469 ( .A1(n408), .A2(n407), .ZN(n409) );
  NAND2_X1 U470 ( .A1(n410), .A2(n409), .ZN(n412) );
  XOR2_X1 U471 ( .A(n413), .B(KEYINPUT99), .Z(n415) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U474 ( .A(n416), .B(G204GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(G8GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n514) );
  NOR2_X1 U479 ( .A1(n525), .A2(n514), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n424), .B(KEYINPUT54), .ZN(n565) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n445) );
  XOR2_X1 U482 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(KEYINPUT97), .B(n429), .Z(n431) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U488 ( .A(n432), .B(KEYINPUT94), .Z(n435) );
  XNOR2_X1 U489 ( .A(n433), .B(KEYINPUT6), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U491 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n437) );
  XNOR2_X1 U492 ( .A(G85GAT), .B(KEYINPUT92), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n461) );
  XNOR2_X1 U498 ( .A(KEYINPUT98), .B(n461), .ZN(n563) );
  NAND2_X1 U499 ( .A1(n565), .A2(n563), .ZN(n446) );
  NOR2_X1 U500 ( .A1(n463), .A2(n446), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  NAND2_X1 U502 ( .A1(n531), .A2(n557), .ZN(n452) );
  XOR2_X1 U503 ( .A(G176GAT), .B(KEYINPUT56), .Z(n450) );
  XNOR2_X1 U504 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n449) );
  XOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n454) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n474) );
  NOR2_X1 U508 ( .A1(n529), .A2(n514), .ZN(n455) );
  NOR2_X1 U509 ( .A1(n463), .A2(n455), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(KEYINPUT25), .ZN(n459) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(n514), .ZN(n462) );
  NAND2_X1 U512 ( .A1(n463), .A2(n529), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT26), .ZN(n561) );
  OR2_X1 U514 ( .A1(n462), .A2(n561), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n461), .A2(n460), .ZN(n468) );
  NOR2_X1 U517 ( .A1(n462), .A2(n563), .ZN(n523) );
  XNOR2_X1 U518 ( .A(KEYINPUT67), .B(KEYINPUT28), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n527) );
  NAND2_X1 U520 ( .A1(n523), .A2(n527), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT100), .B(n465), .Z(n466) );
  NAND2_X1 U522 ( .A1(n466), .A2(n529), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n483) );
  INV_X1 U524 ( .A(n484), .ZN(n575) );
  NAND2_X1 U525 ( .A1(n469), .A2(n575), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  AND2_X1 U527 ( .A1(n483), .A2(n471), .ZN(n500) );
  INV_X1 U528 ( .A(n567), .ZN(n499) );
  NOR2_X1 U529 ( .A1(n572), .A2(n499), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT76), .ZN(n487) );
  NAND2_X1 U531 ( .A1(n500), .A2(n487), .ZN(n480) );
  NOR2_X1 U532 ( .A1(n563), .A2(n480), .ZN(n473) );
  XOR2_X1 U533 ( .A(n474), .B(n473), .Z(G1324GAT) );
  NOR2_X1 U534 ( .A1(n514), .A2(n480), .ZN(n476) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n529), .A2(n480), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n479), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n527), .A2(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(G1327GAT) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT37), .B(n486), .Z(n511) );
  NAND2_X1 U546 ( .A1(n511), .A2(n487), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(n488), .ZN(n497) );
  NOR2_X1 U548 ( .A1(n497), .A2(n563), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n497), .A2(n514), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1329GAT) );
  NOR2_X1 U555 ( .A1(n497), .A2(n529), .ZN(n495) );
  XNOR2_X1 U556 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U558 ( .A(G43GAT), .B(n496), .Z(G1330GAT) );
  NOR2_X1 U559 ( .A1(n497), .A2(n527), .ZN(n498) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n498), .Z(G1331GAT) );
  AND2_X1 U561 ( .A1(n499), .A2(n531), .ZN(n510) );
  NAND2_X1 U562 ( .A1(n510), .A2(n500), .ZN(n506) );
  NOR2_X1 U563 ( .A1(n563), .A2(n506), .ZN(n501) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n501), .Z(n502) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n506), .ZN(n503) );
  XOR2_X1 U567 ( .A(KEYINPUT110), .B(n503), .Z(n504) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U569 ( .A1(n529), .A2(n506), .ZN(n505) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n527), .A2(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  NAND2_X1 U575 ( .A1(n511), .A2(n510), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n563), .A2(n519), .ZN(n512) );
  XOR2_X1 U577 ( .A(KEYINPUT112), .B(n512), .Z(n513) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n519), .ZN(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U583 ( .A1(n529), .A2(n519), .ZN(n518) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U585 ( .A1(n527), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT115), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  INV_X1 U589 ( .A(n523), .ZN(n524) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(KEYINPUT116), .B(n526), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n527), .A2(n541), .ZN(n528) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n538), .A2(n567), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n533) );
  NAND2_X1 U597 ( .A1(n538), .A2(n531), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n536) );
  NAND2_X1 U601 ( .A1(n538), .A2(n575), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n537), .Z(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n558), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  INV_X1 U607 ( .A(n541), .ZN(n542) );
  NOR2_X1 U608 ( .A1(n561), .A2(n542), .ZN(n550) );
  AND2_X1 U609 ( .A1(n567), .A2(n550), .ZN(n543) );
  XOR2_X1 U610 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  XOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .Z(n546) );
  NAND2_X1 U612 ( .A1(n550), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n575), .A2(n550), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n552) );
  NAND2_X1 U619 ( .A1(n550), .A2(n558), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n567), .ZN(n554) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT123), .Z(n556) );
  NAND2_X1 U625 ( .A1(n557), .A2(n575), .ZN(n555) );
  XNOR2_X1 U626 ( .A(n556), .B(n555), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .Z(n569) );
  INV_X1 U631 ( .A(n561), .ZN(n562) );
  AND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n578), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n578), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n291), .ZN(G1355GAT) );
endmodule

