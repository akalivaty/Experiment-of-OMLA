

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  INV_X1 U321 ( .A(KEYINPUT102), .ZN(n413) );
  XNOR2_X1 U322 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U323 ( .A(n462), .B(KEYINPUT111), .ZN(n463) );
  INV_X1 U324 ( .A(KEYINPUT93), .ZN(n332) );
  XNOR2_X1 U325 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n469) );
  XNOR2_X1 U326 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U327 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U328 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U329 ( .A(n335), .B(n334), .ZN(n338) );
  XNOR2_X1 U330 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U331 ( .A(n416), .B(KEYINPUT103), .ZN(n417) );
  XNOR2_X1 U332 ( .A(n418), .B(n417), .ZN(n516) );
  XNOR2_X1 U333 ( .A(n348), .B(n370), .ZN(n520) );
  XNOR2_X1 U334 ( .A(n478), .B(G176GAT), .ZN(n479) );
  XNOR2_X1 U335 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n451) );
  XNOR2_X1 U336 ( .A(n480), .B(n479), .ZN(G1349GAT) );
  XNOR2_X1 U337 ( .A(n452), .B(n451), .ZN(G1329GAT) );
  XOR2_X1 U338 ( .A(G134GAT), .B(KEYINPUT72), .Z(n312) );
  XOR2_X1 U339 ( .A(G36GAT), .B(G190GAT), .Z(n335) );
  XOR2_X1 U340 ( .A(n312), .B(n335), .Z(n290) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U342 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U343 ( .A(G92GAT), .B(KEYINPUT10), .Z(n292) );
  XNOR2_X1 U344 ( .A(KEYINPUT9), .B(KEYINPUT71), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U346 ( .A(n294), .B(n293), .Z(n299) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n379) );
  XOR2_X1 U348 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U349 ( .A(G218GAT), .B(KEYINPUT64), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n379), .B(n297), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U353 ( .A(G29GAT), .B(G43GAT), .Z(n301) );
  XNOR2_X1 U354 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n432) );
  XOR2_X1 U356 ( .A(G85GAT), .B(KEYINPUT69), .Z(n303) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(G106GAT), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n439) );
  XOR2_X1 U359 ( .A(n432), .B(n439), .Z(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n555) );
  XNOR2_X1 U361 ( .A(KEYINPUT36), .B(n555), .ZN(n583) );
  XOR2_X1 U362 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U365 ( .A(KEYINPUT90), .B(n308), .Z(n310) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U368 ( .A(n311), .B(KEYINPUT87), .Z(n319) );
  XOR2_X1 U369 ( .A(n312), .B(G85GAT), .Z(n316) );
  XOR2_X1 U370 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n314) );
  XNOR2_X1 U371 ( .A(G141GAT), .B(KEYINPUT85), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n369) );
  XNOR2_X1 U373 ( .A(n369), .B(G162GAT), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n317), .B(KEYINPUT6), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U377 ( .A(G155GAT), .B(G148GAT), .Z(n321) );
  XNOR2_X1 U378 ( .A(G29GAT), .B(G1GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U381 ( .A(KEYINPUT77), .B(G127GAT), .Z(n325) );
  XNOR2_X1 U382 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U384 ( .A(G113GAT), .B(n326), .Z(n358) );
  XOR2_X1 U385 ( .A(KEYINPUT91), .B(KEYINPUT88), .Z(n328) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(KEYINPUT89), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n358), .B(n329), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n527) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XOR2_X1 U391 ( .A(G64GAT), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U392 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n438) );
  XOR2_X1 U394 ( .A(n338), .B(n438), .Z(n343) );
  XOR2_X1 U395 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n340) );
  XNOR2_X1 U396 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n351) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n341), .B(KEYINPUT74), .ZN(n399) );
  XNOR2_X1 U400 ( .A(n351), .B(n399), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n348) );
  XNOR2_X1 U402 ( .A(G211GAT), .B(KEYINPUT83), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n344), .B(KEYINPUT21), .ZN(n345) );
  XOR2_X1 U404 ( .A(n345), .B(KEYINPUT84), .Z(n347) );
  XNOR2_X1 U405 ( .A(G197GAT), .B(G218GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n370) );
  INV_X1 U407 ( .A(KEYINPUT27), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n520), .B(n349), .ZN(n350) );
  XOR2_X1 U409 ( .A(n350), .B(KEYINPUT94), .Z(n390) );
  XOR2_X1 U410 ( .A(n351), .B(G99GAT), .Z(n353) );
  NAND2_X1 U411 ( .A1(G227GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U413 ( .A(n354), .B(G134GAT), .Z(n360) );
  XOR2_X1 U414 ( .A(G176GAT), .B(G183GAT), .Z(n356) );
  XNOR2_X1 U415 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n368) );
  XOR2_X1 U419 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n362) );
  XNOR2_X1 U420 ( .A(KEYINPUT78), .B(KEYINPUT20), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U422 ( .A(KEYINPUT79), .B(G71GAT), .Z(n364) );
  XNOR2_X1 U423 ( .A(G43GAT), .B(G190GAT), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U425 ( .A(n366), .B(n365), .Z(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n391) );
  INV_X1 U427 ( .A(n391), .ZN(n530) );
  XOR2_X1 U428 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n372) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U431 ( .A(G148GAT), .B(G78GAT), .Z(n442) );
  XOR2_X1 U432 ( .A(G22GAT), .B(G155GAT), .Z(n398) );
  XOR2_X1 U433 ( .A(n442), .B(n398), .Z(n374) );
  NAND2_X1 U434 ( .A1(G228GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U436 ( .A(n376), .B(n375), .Z(n382) );
  XOR2_X1 U437 ( .A(G204GAT), .B(KEYINPUT24), .Z(n378) );
  XNOR2_X1 U438 ( .A(G106GAT), .B(KEYINPUT86), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n472) );
  NOR2_X1 U442 ( .A1(n530), .A2(n472), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n383), .B(KEYINPUT26), .ZN(n567) );
  AND2_X1 U444 ( .A1(n390), .A2(n567), .ZN(n546) );
  XNOR2_X1 U445 ( .A(KEYINPUT96), .B(n546), .ZN(n387) );
  NAND2_X1 U446 ( .A1(n530), .A2(n520), .ZN(n384) );
  NAND2_X1 U447 ( .A1(n472), .A2(n384), .ZN(n385) );
  XNOR2_X1 U448 ( .A(KEYINPUT25), .B(n385), .ZN(n386) );
  NOR2_X1 U449 ( .A1(n387), .A2(n386), .ZN(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT97), .B(n388), .Z(n389) );
  NOR2_X1 U451 ( .A1(n527), .A2(n389), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n472), .B(KEYINPUT28), .ZN(n494) );
  NAND2_X1 U453 ( .A1(n390), .A2(n494), .ZN(n532) );
  NAND2_X1 U454 ( .A1(n527), .A2(n391), .ZN(n392) );
  NOR2_X1 U455 ( .A1(n532), .A2(n392), .ZN(n393) );
  XOR2_X1 U456 ( .A(KEYINPUT95), .B(n393), .Z(n394) );
  NOR2_X1 U457 ( .A1(n395), .A2(n394), .ZN(n482) );
  XNOR2_X1 U458 ( .A(G15GAT), .B(G1GAT), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n396), .B(KEYINPUT66), .ZN(n419) );
  XOR2_X1 U460 ( .A(G71GAT), .B(G57GAT), .Z(n397) );
  XOR2_X1 U461 ( .A(KEYINPUT13), .B(n397), .Z(n448) );
  XNOR2_X1 U462 ( .A(n419), .B(n448), .ZN(n412) );
  XOR2_X1 U463 ( .A(n399), .B(n398), .Z(n401) );
  XNOR2_X1 U464 ( .A(G127GAT), .B(G78GAT), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U466 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n403) );
  NAND2_X1 U467 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U469 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U470 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n407) );
  XNOR2_X1 U471 ( .A(G211GAT), .B(G64GAT), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n408), .B(KEYINPUT76), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n552) );
  INV_X1 U476 ( .A(n552), .ZN(n579) );
  NOR2_X1 U477 ( .A1(n482), .A2(n579), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U479 ( .A1(n583), .A2(n415), .ZN(n418) );
  INV_X1 U480 ( .A(KEYINPUT37), .ZN(n416) );
  XOR2_X1 U481 ( .A(G50GAT), .B(n419), .Z(n421) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U484 ( .A(n422), .B(G36GAT), .Z(n430) );
  XOR2_X1 U485 ( .A(G197GAT), .B(G22GAT), .Z(n424) );
  XNOR2_X1 U486 ( .A(G169GAT), .B(G113GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U488 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n426) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(G8GAT), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n431), .B(KEYINPUT29), .ZN(n434) );
  XOR2_X1 U494 ( .A(n432), .B(KEYINPUT30), .Z(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n570) );
  XNOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT32), .ZN(n436) );
  AND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U499 ( .A(n437), .B(KEYINPUT31), .Z(n441) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n446) );
  XNOR2_X1 U502 ( .A(G120GAT), .B(n442), .ZN(n444) );
  INV_X1 U503 ( .A(KEYINPUT33), .ZN(n443) );
  XOR2_X1 U504 ( .A(n448), .B(n447), .Z(n575) );
  NOR2_X1 U505 ( .A1(n570), .A2(n575), .ZN(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT70), .B(n449), .Z(n485) );
  NOR2_X1 U507 ( .A1(n516), .A2(n485), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n450), .B(KEYINPUT38), .ZN(n502) );
  NAND2_X1 U509 ( .A1(n502), .A2(n520), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n474) );
  NOR2_X1 U511 ( .A1(n583), .A2(n552), .ZN(n454) );
  XNOR2_X1 U512 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n570), .A2(n455), .ZN(n456) );
  NOR2_X1 U515 ( .A1(n575), .A2(n456), .ZN(n457) );
  XOR2_X1 U516 ( .A(KEYINPUT113), .B(n457), .Z(n466) );
  XNOR2_X1 U517 ( .A(KEYINPUT41), .B(n575), .ZN(n477) );
  NOR2_X1 U518 ( .A1(n570), .A2(n477), .ZN(n459) );
  INV_X1 U519 ( .A(KEYINPUT46), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT110), .B(n579), .ZN(n559) );
  INV_X1 U522 ( .A(n555), .ZN(n562) );
  NOR2_X1 U523 ( .A1(n559), .A2(n562), .ZN(n460) );
  NAND2_X1 U524 ( .A1(n461), .A2(n460), .ZN(n464) );
  INV_X1 U525 ( .A(KEYINPUT47), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT48), .ZN(n529) );
  XOR2_X1 U528 ( .A(n520), .B(KEYINPUT118), .Z(n468) );
  NOR2_X1 U529 ( .A1(n529), .A2(n468), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n527), .A2(n471), .ZN(n568) );
  NAND2_X1 U531 ( .A1(n568), .A2(n472), .ZN(n473) );
  XOR2_X1 U532 ( .A(n474), .B(n473), .Z(n475) );
  AND2_X1 U533 ( .A1(n475), .A2(n530), .ZN(n476) );
  XOR2_X1 U534 ( .A(n476), .B(KEYINPUT121), .Z(n563) );
  INV_X1 U535 ( .A(n477), .ZN(n535) );
  NAND2_X1 U536 ( .A1(n563), .A2(n535), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n478) );
  NOR2_X1 U538 ( .A1(n562), .A2(n552), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n481), .B(KEYINPUT16), .ZN(n484) );
  INV_X1 U540 ( .A(n482), .ZN(n483) );
  NAND2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n505) );
  NOR2_X1 U542 ( .A1(n485), .A2(n505), .ZN(n495) );
  NAND2_X1 U543 ( .A1(n495), .A2(n527), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n486), .B(KEYINPUT34), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n489) );
  NAND2_X1 U547 ( .A1(n495), .A2(n520), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U551 ( .A1(n495), .A2(n530), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  XOR2_X1 U554 ( .A(G22GAT), .B(KEYINPUT101), .Z(n497) );
  INV_X1 U555 ( .A(n494), .ZN(n523) );
  NAND2_X1 U556 ( .A1(n495), .A2(n523), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  NAND2_X1 U559 ( .A1(n527), .A2(n502), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n502), .A2(n530), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT40), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n502), .A2(n523), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n507) );
  NAND2_X1 U567 ( .A1(n535), .A2(n570), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(KEYINPUT106), .ZN(n517) );
  NOR2_X1 U569 ( .A1(n517), .A2(n505), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n512), .A2(n527), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n520), .A2(n512), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT107), .Z(n511) );
  NAND2_X1 U576 ( .A1(n512), .A2(n530), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n523), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  XOR2_X1 U582 ( .A(G85GAT), .B(KEYINPUT109), .Z(n519) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n524), .A2(n527), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n524), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n530), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  INV_X1 U593 ( .A(n570), .ZN(n557) );
  INV_X1 U594 ( .A(n527), .ZN(n528) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n530), .A2(n545), .ZN(n531) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n557), .A2(n542), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT114), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U602 ( .A1(n542), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U606 ( .A1(n542), .A2(n559), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U610 ( .A1(n542), .A2(n562), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n554) );
  NOR2_X1 U613 ( .A1(n570), .A2(n554), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n477), .A2(n554), .ZN(n550) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n552), .A2(n554), .ZN(n553) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n563), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(n561), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(KEYINPUT124), .B(n569), .ZN(n582) );
  NOR2_X1 U635 ( .A1(n582), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U641 ( .A(n582), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n575), .A2(n580), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

