//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  AND2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT69), .Z(G261));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT70), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(KEYINPUT70), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n457), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n465), .B2(new_n466), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n494), .B(new_n497), .C1(new_n466), .C2(new_n465), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(G164));
  AND2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(new_n503), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n501), .A2(new_n500), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n507), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n515), .A2(new_n516), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n525), .A2(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n513), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT72), .B(G52), .Z(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n523), .A2(new_n533), .B1(new_n517), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  INV_X1    g112(.A(G68), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n526), .A2(new_n537), .B1(new_n538), .B2(new_n503), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI221_X1 g116(.A(KEYINPUT73), .B1(new_n538), .B2(new_n503), .C1(new_n526), .C2(new_n537), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(G651), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n517), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT74), .B(G43), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n544), .A2(G81), .B1(new_n504), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n509), .B2(new_n510), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT76), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n559), .B(new_n556), .C1(new_n526), .C2(new_n554), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(G651), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n517), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n511), .A2(new_n522), .A3(new_n564), .A4(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n561), .A2(new_n566), .A3(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  INV_X1    g147(.A(G49), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n523), .A2(KEYINPUT77), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT77), .B1(new_n523), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n511), .A2(G74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n544), .B2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G288));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n523), .A2(new_n580), .B1(new_n517), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n511), .A2(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n513), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n526), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(G72), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n544), .A2(G85), .B1(new_n504), .B2(G47), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n591), .A2(new_n592), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n526), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n603), .B(new_n599), .C1(new_n526), .C2(new_n600), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(G651), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n517), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n504), .A2(G54), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n598), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n598), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n547), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n612), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n477), .A2(new_n478), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n472), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n479), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n481), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n464), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n633), .A2(new_n634), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XOR2_X1   g220(.A(G2427), .B(G2430), .Z(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n632), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n640), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n675), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n679), .C1(new_n672), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(G229));
  NAND2_X1  g264(.A1(new_n613), .A2(G16), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G4), .B2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G1348), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G35), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G162), .B2(new_n694), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT29), .Z(new_n697));
  INV_X1    g272(.A(G2090), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n692), .B2(new_n691), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(G27), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G164), .B2(new_n694), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT93), .Z(new_n703));
  AOI211_X1 g278(.A(new_n693), .B(new_n700), .C1(G2078), .C2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n694), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n481), .A2(G129), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n472), .A2(G105), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G141), .B2(new_n479), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT26), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n705), .B1(new_n714), .B2(new_n694), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT27), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1996), .ZN(new_n717));
  OAI22_X1  g292(.A1(new_n697), .A2(new_n698), .B1(new_n703), .B2(G2078), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G19), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n548), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT87), .B(G1341), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n704), .A2(new_n717), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n694), .A2(G33), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT88), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n479), .A2(G139), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n728), .B(new_n729), .C1(new_n464), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n694), .A2(G26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n479), .A2(G140), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n481), .A2(G128), .ZN(new_n738));
  OR2_X1    g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(new_n694), .ZN(new_n743));
  INV_X1    g318(.A(G2067), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT31), .B(G11), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n748), .A2(G28), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n694), .B1(new_n748), .B2(G28), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n747), .B1(new_n749), .B2(new_n750), .C1(new_n639), .C2(new_n694), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(G160), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n694), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n751), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n734), .A2(new_n745), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n760), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n760), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n765), .A2(G1961), .B1(new_n752), .B2(new_n757), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n763), .B(new_n766), .C1(G1961), .C2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n762), .A2(G1966), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT91), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n732), .A2(new_n733), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT89), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n760), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n617), .B2(new_n760), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n724), .A2(new_n759), .A3(new_n770), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G6), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n586), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  INV_X1    g357(.A(G1981), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n760), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n760), .ZN(new_n786));
  INV_X1    g361(.A(G1971), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n760), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(G288), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n760), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT33), .B(G1976), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n784), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n796));
  NOR2_X1   g371(.A1(G25), .A2(G29), .ZN(new_n797));
  AOI22_X1  g372(.A1(G119), .A2(new_n481), .B1(new_n479), .B2(G131), .ZN(new_n798));
  OR2_X1    g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(KEYINPUT83), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(KEYINPUT83), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT84), .Z(new_n804));
  AOI21_X1  g379(.A(new_n797), .B1(new_n804), .B2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT85), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n760), .A2(G24), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n595), .A2(new_n596), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n760), .ZN(new_n811));
  AOI21_X1  g386(.A(KEYINPUT86), .B1(new_n811), .B2(G1986), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G1986), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n795), .A2(new_n796), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n779), .A2(new_n817), .A3(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  NOR2_X1   g395(.A1(new_n612), .A2(new_n620), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n523), .A2(new_n824), .B1(new_n517), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n511), .A2(G67), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n513), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n830), .A2(new_n543), .A3(new_n546), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n543), .B2(new_n546), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n823), .B(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n830), .A2(new_n836), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT95), .B(KEYINPUT37), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(G145));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n479), .A2(G142), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n481), .A2(G130), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n464), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT97), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n630), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n804), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n804), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n713), .A2(new_n741), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n713), .A2(new_n741), .ZN(new_n857));
  OAI21_X1  g432(.A(G164), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n496), .A2(new_n498), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n487), .A2(new_n491), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n862), .A3(new_n855), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n858), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n858), .A2(new_n863), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n731), .B(KEYINPUT96), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n854), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT99), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n868), .A2(new_n865), .B1(new_n851), .B2(new_n852), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n756), .B(new_n639), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n485), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT100), .Z(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n854), .A2(new_n876), .A3(new_n865), .A4(new_n868), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n873), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n871), .B1(new_n869), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n854), .A2(KEYINPUT98), .A3(new_n865), .A4(new_n868), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n843), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n869), .A2(new_n882), .ZN(new_n887));
  INV_X1    g462(.A(new_n871), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n873), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n890), .A2(KEYINPUT40), .A3(new_n879), .A4(new_n878), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n886), .A2(new_n891), .ZN(G395));
  NOR2_X1   g467(.A1(new_n830), .A2(G868), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT101), .B1(new_n831), .B2(new_n832), .ZN(new_n895));
  INV_X1    g470(.A(new_n830), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n547), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n830), .A2(new_n543), .A3(new_n546), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n895), .A2(new_n624), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n624), .B1(new_n895), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G299), .A2(KEYINPUT102), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n561), .A2(new_n566), .A3(new_n568), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n613), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n612), .A2(KEYINPUT102), .A3(G299), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n910), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n901), .B2(new_n902), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n918));
  NAND2_X1  g493(.A1(G290), .A2(G288), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n810), .A2(new_n790), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G166), .B(G305), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n918), .A3(new_n920), .ZN(new_n924));
  XNOR2_X1  g499(.A(G166), .B(new_n586), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n923), .B(KEYINPUT42), .C1(new_n926), .C2(new_n921), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n916), .A2(new_n917), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n916), .A2(new_n917), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n913), .A2(KEYINPUT104), .A3(new_n915), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n919), .A2(new_n920), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT103), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n924), .A3(new_n925), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT42), .B1(new_n938), .B2(new_n923), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n931), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n894), .B1(new_n941), .B2(new_n622), .ZN(G295));
  AND3_X1   g517(.A1(new_n913), .A2(KEYINPUT104), .A3(new_n915), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT104), .B1(new_n913), .B2(new_n915), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n929), .A2(new_n930), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n932), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n622), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT105), .B1(new_n948), .B2(new_n893), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(new_n894), .C1(new_n941), .C2(new_n622), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(G331));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n953));
  NAND2_X1  g528(.A1(G171), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n831), .B2(new_n832), .ZN(new_n956));
  AOI21_X1  g531(.A(G168), .B1(G301), .B2(KEYINPUT106), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n897), .A2(new_n954), .A3(new_n899), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n909), .B(new_n912), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n958), .ZN(new_n962));
  INV_X1    g537(.A(new_n957), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n956), .A2(new_n958), .A3(new_n957), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n914), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(KEYINPUT107), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n971), .B2(new_n927), .ZN(new_n972));
  INV_X1    g547(.A(new_n927), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT43), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n974), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n967), .A2(new_n927), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n879), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT44), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n972), .B2(new_n974), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n976), .A2(KEYINPUT43), .A3(new_n979), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(G8), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(G166), .B2(new_n987), .ZN(new_n990));
  OAI211_X1 g565(.A(G8), .B(new_n988), .C1(new_n507), .C2(new_n518), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n862), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n470), .A2(new_n473), .ZN(new_n997));
  INV_X1    g572(.A(G125), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n477), .B2(new_n478), .ZN(new_n999));
  INV_X1    g574(.A(new_n468), .ZN(new_n1000));
  OAI21_X1  g575(.A(G2105), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1001), .A3(G40), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n994), .A2(new_n996), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n1009));
  AND4_X1   g584(.A1(KEYINPUT109), .A2(new_n997), .A3(new_n1001), .A4(G40), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n994), .A4(new_n996), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1008), .A2(new_n1012), .A3(new_n787), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n862), .B2(new_n995), .ZN(new_n1015));
  AOI211_X1 g590(.A(KEYINPUT50), .B(G1384), .C1(new_n860), .C2(new_n861), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(new_n698), .A3(new_n1011), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n987), .B(new_n992), .C1(new_n1013), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n992), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G164), .A2(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(new_n987), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n582), .A2(new_n585), .A3(G1981), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT49), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G61), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n526), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n584), .ZN(new_n1032));
  OAI21_X1  g607(.A(G651), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n544), .A2(G86), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n504), .A2(G48), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n783), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT116), .A3(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1029), .B(new_n1038), .C1(new_n783), .C2(new_n586), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n586), .A2(new_n783), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1036), .A2(KEYINPUT116), .A3(new_n1037), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1037), .B1(new_n1036), .B2(KEYINPUT116), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1026), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n790), .A2(G1976), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1045), .A2(new_n1047), .A3(G8), .A4(new_n1024), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1024), .B(G8), .C1(new_n1046), .C2(G288), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1019), .A2(new_n1022), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n862), .A2(new_n995), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1053), .A2(KEYINPUT108), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n1053), .B2(KEYINPUT108), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2078), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1057), .A2(KEYINPUT53), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1002), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(G160), .A2(KEYINPUT125), .A3(G40), .ZN(new_n1061));
  AND4_X1   g636(.A1(new_n996), .A2(new_n1058), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1063));
  INV_X1    g638(.A(new_n498), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n497), .B1(new_n628), .B2(new_n494), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1014), .B(new_n995), .C1(new_n1066), .C2(new_n492), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1063), .A2(new_n1067), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT124), .B(G1961), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1056), .A2(new_n1062), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(G2078), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(KEYINPUT53), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G171), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1006), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT123), .A3(new_n1057), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1006), .B2(G2078), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(KEYINPUT53), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1078), .B(new_n1079), .C1(KEYINPUT53), .C2(new_n1071), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1073), .B(KEYINPUT54), .C1(new_n1080), .C2(G171), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1052), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  AND3_X1   g658(.A1(G299), .A2(new_n1083), .A3(KEYINPUT57), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(G299), .B2(new_n1083), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1068), .A2(new_n776), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1011), .A2(new_n994), .A3(new_n996), .A4(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1086), .A2(KEYINPUT120), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1025), .A2(new_n744), .B1(new_n1068), .B2(new_n692), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(new_n612), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1097), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1090), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1068), .A2(new_n692), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1011), .A2(new_n744), .A3(new_n1023), .ZN(new_n1102));
  AND4_X1   g677(.A1(KEYINPUT60), .A2(new_n1101), .A3(new_n612), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n612), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1095), .A2(KEYINPUT60), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1103), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1097), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1100), .B(new_n1108), .C1(new_n1109), .C2(KEYINPUT61), .ZN(new_n1110));
  INV_X1    g685(.A(G1996), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1024), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1006), .B2(G1996), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n548), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1117), .B2(new_n548), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1098), .B1(new_n1110), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT118), .B1(new_n1068), .B2(G2084), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1017), .A2(new_n1124), .A3(new_n752), .A4(new_n1011), .ZN(new_n1125));
  INV_X1    g700(.A(G1966), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1006), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(G8), .A3(G286), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(G8), .C1(new_n1128), .C2(G286), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1129), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1080), .A2(G171), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1072), .A2(G171), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1082), .A2(new_n1122), .A3(new_n1135), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(KEYINPUT62), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1143), .B(new_n1129), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1144));
  NOR4_X1   g719(.A1(new_n1136), .A2(new_n1022), .A3(new_n1019), .A4(new_n1051), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1051), .A2(KEYINPUT117), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1044), .A2(new_n1148), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1019), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1044), .A2(new_n1046), .A3(new_n790), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1026), .B1(new_n1152), .B2(new_n1027), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1022), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1021), .A2(new_n1020), .A3(G8), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1051), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1128), .A2(G8), .A3(G168), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1162), .A2(new_n1150), .A3(KEYINPUT63), .A4(new_n1158), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1154), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1141), .A2(new_n1146), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1055), .A2(new_n1011), .A3(new_n1054), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT110), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT110), .A4(new_n1011), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT112), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n741), .B(new_n744), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n714), .B2(new_n1111), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT112), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1168), .A2(new_n1174), .A3(new_n1169), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1171), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1168), .A2(new_n1111), .A3(new_n1169), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1177), .A2(new_n713), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT113), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(KEYINPUT113), .A3(new_n1178), .ZN(new_n1182));
  INV_X1    g757(.A(new_n807), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n804), .A2(new_n1183), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n804), .A2(new_n1183), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1171), .B(new_n1175), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1181), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1170), .ZN(new_n1188));
  NOR2_X1   g763(.A1(G290), .A2(G1986), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1189), .A2(KEYINPUT111), .ZN(new_n1190));
  NAND2_X1  g765(.A1(G290), .A2(G1986), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1190), .B(new_n1191), .Z(new_n1192));
  AOI21_X1  g767(.A(new_n1187), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1165), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1181), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n742), .A2(new_n744), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1177), .B(KEYINPUT46), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n714), .A2(new_n1172), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1199), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(KEYINPUT47), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT47), .ZN(new_n1204));
  OAI211_X1 g779(.A(new_n1199), .B(new_n1204), .C1(new_n1195), .C2(new_n1201), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1207));
  XOR2_X1   g782(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1208));
  XNOR2_X1  g783(.A(new_n1207), .B(new_n1208), .ZN(new_n1209));
  AND4_X1   g784(.A1(new_n1181), .A2(new_n1209), .A3(new_n1182), .A4(new_n1186), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1198), .A2(new_n1206), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1194), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g787(.A1(new_n983), .A2(new_n984), .ZN(new_n1214));
  OR3_X1    g788(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1215), .B1(new_n687), .B2(new_n688), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1216), .B1(new_n880), .B2(new_n885), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1214), .A2(new_n1217), .ZN(G308));
  OAI221_X1 g792(.A(new_n1216), .B1(new_n880), .B2(new_n885), .C1(new_n983), .C2(new_n984), .ZN(G225));
endmodule


