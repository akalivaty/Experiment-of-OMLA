//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G50), .A3(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n206), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n211), .A2(new_n222), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n229), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n206), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G50), .A2(G58), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n206), .B1(new_n259), .B2(new_n213), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n252), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n252), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(G50), .B1(new_n206), .B2(G1), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n261), .B1(G50), .B2(new_n262), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G226), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n268), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n283), .A2(G223), .B1(G77), .B2(new_n281), .ZN(new_n284));
  INV_X1    g0084(.A(G222), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AOI211_X1 g0088(.A(new_n274), .B(new_n276), .C1(new_n288), .C2(new_n268), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n267), .B1(new_n289), .B2(G169), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n289), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT67), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n267), .B(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(G190), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n300), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n292), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n268), .A2(new_n273), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n274), .B1(G238), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n306), .B(new_n307), .C1(new_n287), .C2(new_n275), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n268), .ZN(new_n309));
  XOR2_X1   g0109(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n305), .B2(new_n309), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  OR3_X1    g0115(.A1(new_n314), .A2(KEYINPUT14), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n305), .A2(new_n309), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT69), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT69), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n320), .A3(KEYINPUT13), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n319), .A2(G179), .A3(new_n321), .A4(new_n311), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT14), .B1(new_n314), .B2(new_n315), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n325));
  INV_X1    g0125(.A(G77), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n254), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(new_n252), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n263), .A2(new_n213), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n264), .B(G68), .C1(G1), .C2(new_n206), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  AND4_X1   g0135(.A1(G190), .A2(new_n319), .A3(new_n321), .A4(new_n311), .ZN(new_n336));
  INV_X1    g0136(.A(new_n334), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n314), .B2(new_n294), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n253), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT15), .B(G87), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n254), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n252), .ZN(new_n345));
  OAI21_X1  g0145(.A(G77), .B1(new_n206), .B2(G1), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n345), .B1(G77), .B2(new_n262), .C1(new_n265), .C2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n274), .B1(G244), .B2(new_n304), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n286), .A2(G232), .A3(new_n282), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n286), .A2(G1698), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n349), .B1(new_n350), .B2(new_n286), .C1(new_n351), .C2(new_n214), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n268), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n347), .B1(new_n354), .B2(G169), .ZN(new_n355));
  INV_X1    g0155(.A(new_n354), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(G179), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(G200), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n347), .B1(G190), .B2(new_n354), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n303), .A2(new_n335), .A3(new_n340), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n281), .A2(new_n206), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n366), .A2(G68), .ZN(new_n367));
  INV_X1    g0167(.A(G58), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n213), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n223), .ZN(new_n370));
  INV_X1    g0170(.A(G159), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n257), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n363), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT70), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(KEYINPUT70), .B(new_n363), .C1(new_n367), .C2(new_n372), .ZN(new_n376));
  INV_X1    g0176(.A(new_n252), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n372), .B1(new_n366), .B2(G68), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(KEYINPUT16), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n375), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n253), .B1(new_n205), .B2(G20), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n264), .B1(new_n263), .B2(new_n253), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n283), .A2(G226), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT71), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n286), .A2(G223), .A3(new_n282), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(KEYINPUT72), .B1(G33), .B2(G87), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(KEYINPUT72), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n268), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n274), .B1(G232), .B2(new_n304), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G169), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n291), .B2(new_n391), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(G200), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n389), .A2(G190), .A3(new_n390), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n382), .A4(new_n380), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n380), .A2(new_n397), .A3(new_n382), .A4(new_n396), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n383), .A2(new_n403), .A3(new_n393), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n395), .A2(new_n399), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n362), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n366), .A2(G107), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n350), .A2(KEYINPUT6), .A3(G97), .ZN(new_n409));
  XOR2_X1   g0209(.A(G97), .B(G107), .Z(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(KEYINPUT6), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n252), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n262), .A2(G97), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n205), .A2(G33), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n377), .A2(new_n262), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n418), .B2(G97), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n281), .A2(G1698), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT4), .A3(G244), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G283), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(new_n216), .C2(new_n351), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT4), .B1(new_n421), .B2(G244), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n268), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n205), .B(G45), .C1(new_n271), .C2(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT74), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n271), .A2(KEYINPUT5), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n272), .A2(G1), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT74), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT5), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G41), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n268), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(G257), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n270), .A2(new_n434), .A3(new_n428), .A4(new_n429), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n426), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G169), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n291), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n420), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n420), .A2(KEYINPUT73), .ZN(new_n445));
  INV_X1    g0245(.A(new_n440), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G190), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT73), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n414), .A2(new_n448), .A3(new_n419), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n440), .A2(G200), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n445), .A2(new_n447), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G116), .ZN(new_n452));
  INV_X1    g0252(.A(G244), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n452), .B1(new_n351), .B2(new_n453), .C1(new_n214), .C2(new_n287), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n268), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n430), .A2(new_n269), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n216), .B1(new_n272), .B2(G1), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n436), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT75), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n458), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n454), .B2(new_n268), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT75), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n291), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n286), .A2(new_n206), .A3(G68), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n206), .B1(new_n307), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G87), .B2(new_n203), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n467), .B1(new_n254), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n252), .B1(new_n263), .B2(new_n343), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n343), .B2(new_n417), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n463), .B(new_n460), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n465), .B(new_n474), .C1(new_n475), .C2(G169), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n461), .A2(G190), .A3(new_n464), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n418), .A2(G87), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(new_n480), .C1(new_n475), .C2(new_n294), .ZN(new_n481));
  AND4_X1   g0281(.A1(new_n444), .A2(new_n451), .A3(new_n476), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n279), .A2(G33), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n484));
  OAI21_X1  g0284(.A(G303), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n278), .A2(new_n280), .A3(G257), .A4(new_n282), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n278), .A2(new_n280), .A3(G264), .A4(G1698), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n268), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n429), .B1(new_n427), .B2(KEYINPUT74), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n431), .B1(new_n430), .B2(new_n433), .ZN(new_n491));
  OAI211_X1 g0291(.A(G270), .B(new_n436), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n492), .A3(new_n438), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT21), .A3(G169), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n490), .A2(new_n491), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(new_n270), .B1(new_n488), .B2(new_n268), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G179), .A3(new_n492), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n423), .B(new_n206), .C1(G33), .C2(new_n470), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  AOI221_X4 g0300(.A(KEYINPUT76), .B1(new_n500), .B2(G20), .C1(new_n251), .C2(new_n229), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT76), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(G20), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n252), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n499), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(KEYINPUT20), .B(new_n499), .C1(new_n501), .C2(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n263), .A2(G116), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n417), .B2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n498), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT77), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n507), .B2(new_n508), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n494), .B2(new_n497), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT77), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n315), .B1(new_n496), .B2(new_n492), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(new_n521), .A3(KEYINPUT78), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT78), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n493), .A2(G169), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n516), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT79), .A4(new_n526), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n493), .A2(G200), .ZN(new_n532));
  INV_X1    g0332(.A(G190), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n516), .C1(new_n533), .C2(new_n493), .ZN(new_n534));
  OAI211_X1 g0334(.A(G264), .B(new_n436), .C1(new_n490), .C2(new_n491), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n435), .A2(KEYINPUT82), .A3(G264), .A4(new_n436), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n278), .A2(new_n280), .A3(G257), .A4(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n278), .A2(new_n280), .A3(G250), .A4(new_n282), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT81), .A4(new_n542), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n268), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n539), .A2(G190), .A3(new_n438), .A4(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n537), .A3(new_n538), .A4(new_n438), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n278), .A2(new_n280), .A3(new_n206), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT22), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n286), .A2(new_n553), .A3(new_n206), .A4(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n452), .A2(G20), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n206), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n350), .A2(KEYINPUT23), .A3(G20), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n555), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n556), .B1(new_n555), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n252), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n262), .A2(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(KEYINPUT80), .B(KEYINPUT25), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n565), .B(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(G107), .B2(new_n418), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n548), .A2(new_n550), .A3(new_n564), .A4(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n539), .A2(new_n291), .A3(new_n438), .A4(new_n547), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n568), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n549), .A2(new_n315), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n482), .A2(new_n531), .A3(new_n534), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n407), .A2(new_n575), .ZN(G372));
  INV_X1    g0376(.A(new_n358), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n335), .B1(new_n339), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n402), .A2(new_n399), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g0380(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n383), .A2(KEYINPUT84), .A3(new_n393), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT84), .B1(new_n383), .B2(new_n393), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT84), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n394), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n383), .A2(KEYINPUT84), .A3(new_n393), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n581), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n580), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n301), .A2(new_n302), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n292), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT83), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n463), .A2(new_n294), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(new_n479), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n480), .B(KEYINPUT83), .C1(new_n294), .C2(new_n463), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n477), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n459), .A2(new_n315), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n465), .A2(new_n474), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n569), .A2(new_n601), .A3(new_n444), .A4(new_n451), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n517), .B1(new_n529), .B2(new_n530), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n573), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT26), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n446), .A2(G179), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n441), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n445), .A2(new_n449), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n601), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n607), .A2(new_n441), .B1(new_n414), .B2(new_n419), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n611), .A2(new_n476), .A3(new_n481), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n600), .C1(new_n606), .C2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n406), .B1(new_n605), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n593), .A2(new_n614), .ZN(G369));
  NAND3_X1  g0415(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n616), .A2(KEYINPUT27), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(KEYINPUT27), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(G213), .A3(new_n618), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT86), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(KEYINPUT86), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OR3_X1    g0425(.A1(new_n603), .A2(new_n516), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n531), .B(new_n534), .C1(new_n516), .C2(new_n625), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G330), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n629), .A2(KEYINPUT87), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT87), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n628), .B2(G330), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n571), .A2(new_n624), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n569), .A2(new_n573), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT88), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n573), .A2(new_n625), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n569), .A2(new_n573), .A3(new_n639), .A4(new_n635), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT89), .B1(new_n531), .B2(new_n624), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n517), .B(KEYINPUT77), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n524), .A2(new_n516), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT21), .B1(new_n647), .B2(KEYINPUT78), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT79), .B1(new_n648), .B2(new_n525), .ZN(new_n649));
  INV_X1    g0449(.A(new_n530), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n625), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n641), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n573), .A2(new_n624), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n644), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n529), .A2(new_n530), .ZN(new_n658));
  AOI211_X1 g0458(.A(KEYINPUT89), .B(new_n624), .C1(new_n658), .C2(new_n646), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n651), .B2(new_n625), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n655), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(KEYINPUT90), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n643), .A2(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n209), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G1), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n227), .B2(new_n668), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n609), .A2(new_n608), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n598), .A2(new_n600), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n611), .A2(new_n476), .A3(new_n481), .A4(new_n606), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT92), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n600), .B(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n531), .A2(new_n573), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n602), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT29), .B1(new_n681), .B2(new_n624), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n683), .B(new_n625), .C1(new_n605), .C2(new_n613), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT31), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n492), .A2(new_n539), .A3(new_n496), .A4(new_n547), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n443), .A2(new_n475), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT30), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n443), .A2(new_n475), .A3(new_n686), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n440), .A2(new_n291), .A3(new_n493), .A4(new_n459), .ZN(new_n692));
  INV_X1    g0492(.A(new_n549), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT91), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  AOI211_X1 g0497(.A(new_n697), .B(new_n694), .C1(new_n688), .C2(new_n690), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n685), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n699), .A2(new_n624), .B1(new_n575), .B2(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n624), .A2(KEYINPUT31), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n691), .B2(new_n695), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n682), .B(new_n684), .C1(new_n703), .C2(new_n630), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n672), .B1(new_n705), .B2(G1), .ZN(G364));
  AND2_X1   g0506(.A1(new_n206), .A2(G13), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n205), .B1(new_n707), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n667), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n634), .B(new_n711), .C1(G330), .C2(new_n628), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n666), .A2(new_n281), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G355), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G116), .B2(new_n209), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n246), .A2(G45), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n666), .A2(new_n286), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n228), .B2(new_n272), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n229), .B1(G20), .B2(new_n315), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n710), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n206), .A2(new_n291), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n729), .A2(new_n533), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G322), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n281), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n733), .B1(G311), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n728), .A2(G190), .A3(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT94), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n738), .A2(KEYINPUT94), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G326), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n206), .A2(G179), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n533), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n533), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n206), .ZN(new_n750));
  INV_X1    g0550(.A(G294), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n752));
  INV_X1    g0552(.A(G303), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n729), .A2(G190), .A3(new_n294), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT33), .B(G317), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n748), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n745), .A2(new_n734), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT95), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT95), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G329), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n737), .A2(new_n744), .A3(new_n757), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(G159), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n752), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n755), .A2(G68), .B1(G87), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n470), .B2(new_n750), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G50), .B2(new_n743), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n746), .A2(new_n350), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n731), .A2(new_n368), .B1(new_n735), .B2(new_n326), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT93), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n281), .B(new_n773), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n772), .B(new_n776), .C1(new_n775), .C2(new_n774), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n764), .B1(new_n768), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n727), .B1(new_n778), .B2(new_n724), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n723), .B(KEYINPUT98), .Z(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n628), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n712), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  OAI21_X1  g0583(.A(new_n625), .B1(new_n605), .B2(new_n613), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n360), .A2(new_n359), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n347), .A2(new_n624), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n358), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n358), .A2(new_n625), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n784), .B(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n699), .A2(new_n624), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n575), .A2(KEYINPUT31), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n702), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n630), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n710), .B1(new_n792), .B2(new_n798), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n721), .B1(new_n787), .B2(new_n789), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n724), .A2(new_n721), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n750), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G97), .B1(new_n769), .B2(G107), .ZN(new_n806));
  INV_X1    g0606(.A(new_n755), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n215), .B2(new_n746), .C1(new_n747), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n286), .B1(new_n736), .B2(G116), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n751), .B2(new_n731), .C1(new_n761), .C2(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n808), .B(new_n811), .C1(G303), .C2(new_n743), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n286), .B1(new_n750), .B2(new_n368), .ZN(new_n813));
  INV_X1    g0613(.A(G50), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n814), .A2(new_n752), .B1(new_n746), .B2(new_n213), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(new_n762), .C2(G132), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT99), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n730), .A2(G143), .B1(G159), .B2(new_n736), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n255), .B2(new_n807), .C1(new_n742), .C2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n812), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n724), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n710), .B1(G77), .B2(new_n804), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT100), .Z(new_n825));
  AOI22_X1  g0625(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  OR2_X1    g0627(.A1(new_n411), .A2(KEYINPUT35), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n411), .A2(KEYINPUT35), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n828), .A2(G116), .A3(new_n230), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT36), .Z(new_n831));
  OR3_X1    g0631(.A1(new_n227), .A2(new_n326), .A3(new_n369), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n814), .A2(G68), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n205), .B(G13), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n622), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n590), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n373), .A2(new_n379), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n382), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n836), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n405), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n383), .A2(new_n836), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n394), .A2(new_n843), .A3(new_n844), .A4(new_n400), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n393), .A2(new_n839), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n846), .A2(new_n400), .A3(new_n840), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(new_n847), .B2(new_n844), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n625), .B(new_n790), .C1(new_n605), .C2(new_n613), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n788), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n324), .A2(KEYINPUT101), .A3(new_n334), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT101), .B1(new_n324), .B2(new_n334), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n336), .A2(new_n338), .B1(new_n337), .B2(new_n625), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n337), .A2(new_n625), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n324), .B2(new_n339), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n852), .A2(new_n854), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n851), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n865), .A2(new_n849), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n843), .B1(new_n590), .B2(new_n579), .ZN(new_n869));
  INV_X1    g0669(.A(new_n845), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n400), .B(new_n843), .C1(new_n583), .C2(new_n584), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n868), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n851), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n842), .A2(KEYINPUT102), .A3(KEYINPUT38), .A4(new_n848), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n867), .B1(new_n877), .B2(new_n866), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n625), .B1(new_n855), .B2(new_n856), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n837), .B(new_n864), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n682), .A2(new_n684), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n406), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n883), .A2(new_n593), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n881), .B(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n790), .B1(new_n858), .B2(new_n861), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n696), .A2(new_n698), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n701), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n890), .B2(new_n795), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n877), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n886), .B1(new_n865), .B2(new_n849), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n700), .A2(new_n889), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n893), .A2(new_n894), .A3(new_n887), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n407), .B1(new_n795), .B2(new_n890), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n630), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n205), .B2(new_n707), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n885), .A2(new_n900), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n835), .B1(new_n902), .B2(new_n903), .ZN(G367));
  INV_X1    g0704(.A(new_n746), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n805), .A2(G107), .B1(new_n905), .B2(G97), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n751), .B2(new_n807), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n281), .B1(new_n747), .B2(new_n735), .C1(new_n731), .C2(new_n753), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT46), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n769), .A2(G116), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(G317), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n911), .B1(new_n909), .B2(new_n910), .C1(new_n912), .C2(new_n761), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n907), .B(new_n913), .C1(G311), .C2(new_n743), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT104), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n286), .B1(new_n731), .B2(new_n255), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n750), .A2(new_n213), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n368), .A2(new_n752), .B1(new_n746), .B2(new_n326), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n819), .B2(new_n761), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n755), .A2(G159), .B1(G50), .B2(new_n736), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n743), .A2(G143), .B1(KEYINPUT105), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(KEYINPUT105), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n915), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT47), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n724), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n717), .A2(new_n241), .ZN(new_n927));
  INV_X1    g0727(.A(new_n343), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n726), .B1(new_n666), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n711), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n625), .A2(new_n480), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n674), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(new_n465), .A3(new_n474), .A4(new_n599), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n926), .B(new_n930), .C1(new_n780), .C2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n609), .A2(new_n624), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n444), .A3(new_n451), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n609), .A2(new_n608), .A3(new_n624), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n656), .B2(new_n663), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(KEYINPUT45), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n944), .B(new_n941), .C1(new_n656), .C2(new_n663), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n656), .A2(new_n663), .A3(new_n941), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n656), .A2(new_n663), .A3(KEYINPUT44), .A4(new_n941), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n642), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n942), .B(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n643), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n645), .A2(new_n641), .A3(new_n653), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n634), .A2(new_n661), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n661), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n631), .B2(new_n633), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n704), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(new_n705), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n667), .B(KEYINPUT41), .Z(new_n963));
  OAI21_X1  g0763(.A(new_n708), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n941), .B1(KEYINPUT42), .B2(new_n662), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n654), .B2(new_n655), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT42), .B1(new_n661), .B2(new_n941), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n444), .C2(new_n624), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n968), .A2(KEYINPUT103), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT103), .B1(new_n968), .B2(new_n969), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n643), .A2(new_n941), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n936), .B1(new_n964), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(G387));
  NOR2_X1   g0778(.A1(new_n960), .A2(new_n668), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n957), .A2(new_n959), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n705), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n657), .A2(new_n780), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n669), .B(new_n272), .C1(new_n213), .C2(new_n326), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT107), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n253), .A2(G50), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT108), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(KEYINPUT50), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(KEYINPUT50), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n718), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n238), .A2(G45), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT106), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n669), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n713), .A2(new_n995), .B1(new_n350), .B2(new_n666), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n726), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n730), .A2(G317), .B1(G303), .B2(new_n736), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n810), .B2(new_n807), .C1(new_n742), .C2(new_n732), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT48), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n805), .A2(G283), .B1(new_n769), .B2(G294), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n762), .A2(G326), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n286), .B1(new_n905), .B2(G116), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n286), .B1(new_n735), .B2(new_n213), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n807), .A2(new_n253), .B1(new_n326), .B2(new_n752), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G97), .C2(new_n905), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G50), .A2(new_n730), .B1(new_n805), .B2(new_n928), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n743), .A2(G159), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n762), .A2(G150), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n823), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n997), .A2(new_n711), .A3(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n980), .A2(new_n709), .B1(new_n982), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n981), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(G393));
  NAND2_X1  g0825(.A1(new_n961), .A2(new_n667), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n960), .B1(new_n952), .B2(new_n955), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT113), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n952), .A2(new_n955), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n960), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT113), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n667), .A4(new_n961), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n952), .A2(new_n955), .A3(new_n709), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n725), .B1(new_n470), .B2(new_n209), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n717), .B2(new_n249), .ZN(new_n1037));
  INV_X1    g0837(.A(G143), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n761), .A2(new_n1038), .B1(new_n213), .B2(new_n752), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(KEYINPUT112), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n286), .B1(new_n735), .B2(new_n253), .C1(new_n215), .C2(new_n746), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n807), .A2(new_n814), .B1(new_n326), .B2(new_n750), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(KEYINPUT112), .B2(new_n1039), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n742), .A2(new_n255), .B1(new_n371), .B2(new_n731), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT51), .Z(new_n1046));
  OAI22_X1  g0846(.A1(new_n742), .A2(new_n912), .B1(new_n810), .B2(new_n731), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT52), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n807), .A2(new_n753), .B1(new_n752), .B2(new_n747), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G116), .B2(new_n805), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n286), .B(new_n773), .C1(G294), .C2(new_n736), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n732), .C2(new_n761), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1044), .A2(new_n1046), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n711), .B(new_n1037), .C1(new_n1053), .C2(new_n724), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n723), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n940), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1035), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT114), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT114), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1034), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(G390));
  NOR3_X1   g0863(.A1(new_n894), .A2(new_n630), .A3(new_n887), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n590), .A2(new_n579), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n843), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n872), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT38), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n875), .A2(new_n876), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n879), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n602), .A2(new_n680), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n624), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n787), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n789), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT115), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1071), .B1(new_n1078), .B2(new_n863), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n880), .B1(new_n854), .B2(new_n863), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n877), .A2(new_n866), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n867), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1064), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1080), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n875), .A2(new_n876), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n1086), .B2(new_n873), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1087), .B2(new_n867), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n681), .A2(new_n624), .A3(new_n787), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1077), .B1(new_n1089), .B2(new_n789), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n879), .B(new_n877), .C1(new_n1092), .C2(new_n862), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n797), .A2(new_n790), .A3(new_n863), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1088), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1084), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n721), .B1(new_n1087), .B2(new_n867), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n710), .B1(new_n341), .B2(new_n804), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n213), .A2(new_n746), .B1(new_n752), .B2(new_n215), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n281), .B1(new_n470), .B2(new_n735), .C1(new_n731), .C2(new_n500), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n761), .A2(new_n751), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n807), .A2(new_n350), .B1(new_n326), .B2(new_n750), .ZN(new_n1103));
  OR4_X1    g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n742), .A2(new_n747), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n752), .A2(new_n255), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT54), .B(G143), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n286), .B1(new_n735), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G132), .B2(new_n730), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1107), .B(new_n1110), .C1(new_n1111), .C2(new_n761), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n805), .A2(G159), .B1(new_n905), .B2(G50), .ZN(new_n1113));
  INV_X1    g0913(.A(G128), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1113), .B1(new_n819), .B2(new_n807), .C1(new_n742), .C2(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1104), .A2(new_n1105), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1099), .B1(new_n1116), .B2(new_n724), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1097), .A2(new_n709), .B1(new_n1098), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(G330), .B(new_n406), .C1(new_n700), .C2(new_n889), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n883), .A2(new_n593), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n863), .B1(new_n797), .B2(new_n790), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n854), .B1(new_n1121), .B2(new_n1064), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n790), .C1(new_n700), .C2(new_n889), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n862), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1092), .A2(new_n1094), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1120), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1084), .A2(new_n1095), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT116), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1084), .A2(new_n1095), .A3(new_n1126), .A4(KEYINPUT116), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT117), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1126), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n668), .B1(new_n1096), .B2(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1132), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1118), .B1(new_n1135), .B2(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(new_n1120), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1140));
  XNOR2_X1  g0940(.A(new_n303), .B(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n836), .A2(new_n267), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT118), .Z(new_n1143));
  XOR2_X1   g0943(.A(new_n1141), .B(new_n1143), .Z(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n896), .B2(new_n630), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(G330), .C1(new_n892), .C2(new_n895), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n881), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n881), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1139), .A2(KEYINPUT57), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1120), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n1150), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(new_n667), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1144), .A2(new_n721), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n710), .B1(G50), .B2(new_n804), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n286), .A2(G41), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G50), .B(new_n1159), .C1(new_n277), .C2(new_n271), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n807), .A2(new_n470), .B1(new_n746), .B2(new_n368), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n917), .B(new_n1161), .C1(G77), .C2(new_n769), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1159), .B1(new_n343), .B2(new_n735), .C1(new_n731), .C2(new_n350), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G283), .B2(new_n762), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(new_n500), .C2(new_n742), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT58), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1160), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n731), .A2(new_n1114), .B1(new_n735), .B2(new_n819), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G132), .B2(new_n755), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1108), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n805), .A2(G150), .B1(new_n769), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n1111), .C2(new_n742), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n762), .A2(G124), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G33), .B(G41), .C1(new_n905), .C2(G159), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1167), .B1(new_n1166), .B2(new_n1165), .C1(new_n1173), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1158), .B1(new_n1178), .B2(new_n724), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1151), .A2(new_n709), .B1(new_n1157), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1156), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(G375));
  AOI22_X1  g0982(.A1(new_n805), .A2(G50), .B1(new_n905), .B2(G58), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n371), .B2(new_n752), .C1(new_n807), .C2(new_n1108), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n281), .B1(new_n730), .B2(G137), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n255), .B2(new_n735), .C1(new_n761), .C2(new_n1114), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G132), .C2(new_n743), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n805), .A2(new_n928), .B1(new_n905), .B2(G77), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n470), .B2(new_n752), .C1(new_n500), .C2(new_n807), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n286), .B1(new_n736), .B2(G107), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n747), .B2(new_n731), .C1(new_n761), .C2(new_n753), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(G294), .C2(new_n743), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n724), .B1(new_n1187), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n711), .B1(new_n213), .B2(new_n803), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n863), .C2(new_n722), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n709), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1138), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT119), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT119), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1126), .A2(new_n963), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1198), .B1(new_n1202), .B2(new_n1203), .ZN(G381));
  NAND3_X1  g1004(.A1(new_n1023), .A2(new_n782), .A3(new_n1024), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(G384), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1118), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1206), .A2(new_n1208), .A3(G387), .A4(G381), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1209), .A2(new_n1062), .A3(new_n1060), .A4(new_n1181), .ZN(G407));
  INV_X1    g1010(.A(new_n1208), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1181), .A2(G213), .A3(new_n623), .A4(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(G407), .A2(new_n1212), .A3(G213), .ZN(G409));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n623), .A2(G213), .A3(G2897), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n668), .B1(new_n1199), .B2(KEYINPUT60), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT60), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1126), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1217), .B1(new_n1202), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(G384), .A3(new_n1198), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G384), .B1(new_n1220), .B2(new_n1198), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1216), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1223), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n1221), .A3(new_n1215), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1154), .A2(new_n963), .A3(new_n1150), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT120), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1180), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1154), .A2(new_n1150), .A3(KEYINPUT120), .A4(new_n963), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1211), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1156), .A2(G378), .A3(new_n1180), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n623), .A2(G213), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1227), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1214), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1237), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1232), .A2(new_n1233), .B1(G213), .B2(new_n623), .ZN(new_n1240));
  OAI211_X1 g1040(.A(KEYINPUT124), .B(new_n1239), .C1(new_n1240), .C2(new_n1227), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1234), .A2(new_n1235), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT62), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1240), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1238), .A2(new_n1241), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1205), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT121), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G390), .B2(new_n977), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1061), .B1(new_n1034), .B2(new_n1058), .ZN(new_n1253));
  AOI211_X1 g1053(.A(KEYINPUT114), .B(new_n1057), .C1(new_n1028), .C2(new_n1033), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1251), .B(new_n977), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1060), .A2(G387), .A3(new_n1062), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n977), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT122), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(KEYINPUT122), .B(new_n977), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(new_n1249), .A3(new_n1256), .A4(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1258), .A2(KEYINPUT125), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT125), .B1(new_n1258), .B2(new_n1263), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1247), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1243), .B(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1258), .A2(new_n1263), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1236), .A2(KEYINPUT61), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(G405));
  OAI21_X1  g1072(.A(KEYINPUT127), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1259), .A2(KEYINPUT121), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1249), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AND4_X1   g1077(.A1(new_n1249), .A2(new_n1261), .A3(new_n1256), .A4(new_n1262), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1274), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT127), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1258), .A2(KEYINPUT125), .A3(new_n1263), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1233), .B1(new_n1181), .B2(new_n1208), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1242), .A2(KEYINPUT126), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1242), .A2(KEYINPUT126), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1273), .A2(new_n1282), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1273), .B2(new_n1282), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G402));
endmodule


