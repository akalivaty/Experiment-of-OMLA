

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789;

  AND2_X2 U377 ( .A1(n643), .A2(n705), .ZN(n737) );
  NOR2_X1 U378 ( .A1(n788), .A2(n654), .ZN(n587) );
  BUF_X1 U379 ( .A(n661), .Z(n356) );
  NOR2_X1 U380 ( .A1(n588), .A2(n685), .ZN(n575) );
  XNOR2_X1 U381 ( .A(n524), .B(n523), .ZN(n661) );
  XOR2_X1 U382 ( .A(G128), .B(KEYINPUT24), .Z(n513) );
  XNOR2_X1 U383 ( .A(G146), .B(G125), .ZN(n455) );
  INV_X2 U384 ( .A(G953), .ZN(n780) );
  NAND2_X1 U385 ( .A1(n737), .A2(G475), .ZN(n733) );
  NOR2_X2 U386 ( .A1(G953), .A2(G237), .ZN(n496) );
  NAND2_X1 U387 ( .A1(n666), .A2(n665), .ZN(n547) );
  INV_X1 U388 ( .A(n568), .ZN(n673) );
  XNOR2_X1 U389 ( .A(n525), .B(KEYINPUT106), .ZN(n736) );
  NAND2_X1 U390 ( .A1(n398), .A2(n396), .ZN(n525) );
  NAND2_X1 U391 ( .A1(n397), .A2(KEYINPUT64), .ZN(n396) );
  AND2_X1 U392 ( .A1(n402), .A2(n399), .ZN(n398) );
  AND2_X1 U393 ( .A1(n412), .A2(n410), .ZN(n409) );
  NAND2_X1 U394 ( .A1(n377), .A2(KEYINPUT80), .ZN(n380) );
  XNOR2_X1 U395 ( .A(n470), .B(G134), .ZN(n485) );
  INV_X1 U396 ( .A(KEYINPUT75), .ZN(n360) );
  XNOR2_X1 U397 ( .A(n503), .B(n381), .ZN(n644) );
  BUF_X1 U398 ( .A(n736), .Z(n357) );
  BUF_X1 U399 ( .A(n526), .Z(n358) );
  NAND2_X1 U400 ( .A1(n634), .A2(KEYINPUT75), .ZN(n361) );
  NAND2_X1 U401 ( .A1(n359), .A2(n360), .ZN(n362) );
  NAND2_X1 U402 ( .A1(n361), .A2(n362), .ZN(n705) );
  INV_X1 U403 ( .A(n634), .ZN(n359) );
  NAND2_X1 U404 ( .A1(n714), .A2(n437), .ZN(n419) );
  XNOR2_X2 U405 ( .A(n769), .B(n428), .ZN(n432) );
  XNOR2_X2 U406 ( .A(n424), .B(n450), .ZN(n769) );
  OR2_X1 U407 ( .A1(n714), .A2(n417), .ZN(n416) );
  XNOR2_X2 U408 ( .A(n432), .B(n431), .ZN(n714) );
  NOR2_X1 U409 ( .A1(n415), .A2(n684), .ZN(n414) );
  XNOR2_X1 U410 ( .A(n486), .B(n485), .ZN(n778) );
  XOR2_X1 U411 ( .A(KEYINPUT4), .B(G131), .Z(n486) );
  XNOR2_X1 U412 ( .A(G137), .B(G140), .ZN(n509) );
  XNOR2_X1 U413 ( .A(n778), .B(G146), .ZN(n503) );
  XNOR2_X1 U414 ( .A(KEYINPUT65), .B(G101), .ZN(n489) );
  NOR2_X1 U415 ( .A1(n419), .A2(n439), .ZN(n411) );
  XOR2_X1 U416 ( .A(G137), .B(KEYINPUT91), .Z(n498) );
  XNOR2_X1 U417 ( .A(n469), .B(n468), .ZN(n511) );
  XOR2_X1 U418 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n468) );
  NAND2_X1 U419 ( .A1(n380), .A2(n379), .ZN(n469) );
  NAND2_X1 U420 ( .A1(n378), .A2(G234), .ZN(n379) );
  AND2_X1 U421 ( .A1(n477), .A2(n552), .ZN(n686) );
  NAND2_X1 U422 ( .A1(n376), .A2(n593), .ZN(n394) );
  NOR2_X1 U423 ( .A1(n661), .A2(n366), .ZN(n376) );
  INV_X1 U424 ( .A(n365), .ZN(n393) );
  INV_X1 U425 ( .A(KEYINPUT76), .ZN(n395) );
  OR2_X1 U426 ( .A1(n437), .A2(n433), .ZN(n417) );
  INV_X1 U427 ( .A(KEYINPUT0), .ZN(n388) );
  NAND2_X1 U428 ( .A1(n594), .A2(n446), .ZN(n389) );
  XNOR2_X1 U429 ( .A(n507), .B(n506), .ZN(n568) );
  NAND2_X1 U430 ( .A1(n644), .A2(n518), .ZN(n507) );
  XNOR2_X1 U431 ( .A(n593), .B(KEYINPUT1), .ZN(n666) );
  INV_X1 U432 ( .A(G104), .ZN(n421) );
  XNOR2_X1 U433 ( .A(G119), .B(KEYINPUT3), .ZN(n771) );
  XNOR2_X1 U434 ( .A(n363), .B(n503), .ZN(n721) );
  XNOR2_X1 U435 ( .A(KEYINPUT88), .B(KEYINPUT4), .ZN(n429) );
  NAND2_X1 U436 ( .A1(n683), .A2(n375), .ZN(n374) );
  INV_X1 U437 ( .A(n650), .ZN(n375) );
  NAND2_X1 U438 ( .A1(n372), .A2(n369), .ZN(n371) );
  NOR2_X1 U439 ( .A1(G953), .A2(KEYINPUT80), .ZN(n378) );
  NAND2_X1 U440 ( .A1(n780), .A2(G234), .ZN(n377) );
  NAND2_X1 U441 ( .A1(n621), .A2(n610), .ZN(n683) );
  INV_X1 U442 ( .A(G237), .ZN(n434) );
  XOR2_X1 U443 ( .A(G104), .B(G110), .Z(n487) );
  NOR2_X1 U444 ( .A1(n636), .A2(n639), .ZN(n638) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n440) );
  XNOR2_X1 U446 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U447 ( .A1(n409), .A2(n405), .ZN(n594) );
  NAND2_X1 U448 ( .A1(n408), .A2(n406), .ZN(n405) );
  XNOR2_X1 U449 ( .A(n464), .B(n463), .ZN(n551) );
  XNOR2_X1 U450 ( .A(n504), .B(n502), .ZN(n381) );
  XNOR2_X1 U451 ( .A(KEYINPUT97), .B(KEYINPUT11), .ZN(n447) );
  NOR2_X1 U452 ( .A1(n700), .A2(n534), .ZN(n536) );
  INV_X1 U453 ( .A(KEYINPUT104), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n394), .B(n395), .ZN(n572) );
  AND2_X1 U455 ( .A1(n400), .A2(n356), .ZN(n399) );
  NAND2_X1 U456 ( .A1(n401), .A2(KEYINPUT64), .ZN(n400) );
  INV_X1 U457 ( .A(n548), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n551), .B(KEYINPUT100), .ZN(n553) );
  XNOR2_X1 U459 ( .A(n494), .B(G469), .ZN(n382) );
  NOR2_X1 U460 ( .A1(n721), .A2(G902), .ZN(n383) );
  XNOR2_X1 U461 ( .A(n568), .B(KEYINPUT6), .ZN(n605) );
  XOR2_X1 U462 ( .A(KEYINPUT23), .B(G110), .Z(n514) );
  NOR2_X1 U463 ( .A1(n780), .A2(G952), .ZN(n745) );
  XNOR2_X1 U464 ( .A(n528), .B(KEYINPUT32), .ZN(n659) );
  NAND2_X1 U465 ( .A1(n387), .A2(n384), .ZN(n528) );
  XNOR2_X1 U466 ( .A(n386), .B(n385), .ZN(n384) );
  NOR2_X1 U467 ( .A1(n527), .A2(n605), .ZN(n387) );
  OR2_X1 U468 ( .A1(n553), .A2(n552), .ZN(n760) );
  XOR2_X1 U469 ( .A(n493), .B(n492), .Z(n363) );
  INV_X1 U470 ( .A(KEYINPUT19), .ZN(n439) );
  AND2_X1 U471 ( .A1(n626), .A2(n495), .ZN(n364) );
  AND2_X1 U472 ( .A1(n566), .A2(n695), .ZN(n365) );
  OR2_X1 U473 ( .A1(n531), .A2(n393), .ZN(n366) );
  AND2_X1 U474 ( .A1(n358), .A2(n626), .ZN(n367) );
  AND2_X1 U475 ( .A1(n416), .A2(n418), .ZN(n368) );
  OR2_X1 U476 ( .A1(n600), .A2(n599), .ZN(n369) );
  INV_X1 U477 ( .A(G107), .ZN(n488) );
  BUF_X2 U478 ( .A(n737), .Z(n741) );
  NAND2_X1 U479 ( .A1(n481), .A2(n420), .ZN(n484) );
  NOR2_X2 U480 ( .A1(n719), .A2(n745), .ZN(n720) );
  NOR2_X2 U481 ( .A1(n734), .A2(n745), .ZN(n735) );
  NOR2_X2 U482 ( .A1(n728), .A2(n745), .ZN(n729) );
  NOR2_X2 U483 ( .A1(n647), .A2(n745), .ZN(n649) );
  NAND2_X1 U484 ( .A1(n373), .A2(n370), .ZN(n602) );
  NAND2_X1 U485 ( .A1(n683), .A2(n371), .ZN(n370) );
  NAND2_X1 U486 ( .A1(n598), .A2(n597), .ZN(n372) );
  NAND2_X1 U487 ( .A1(n374), .A2(n601), .ZN(n373) );
  NAND2_X1 U488 ( .A1(n553), .A2(n552), .ZN(n610) );
  XNOR2_X2 U489 ( .A(n383), .B(n382), .ZN(n593) );
  NAND2_X1 U490 ( .A1(n614), .A2(n356), .ZN(n386) );
  INV_X1 U491 ( .A(n481), .ZN(n534) );
  XNOR2_X2 U492 ( .A(n389), .B(n388), .ZN(n481) );
  NAND2_X1 U493 ( .A1(n390), .A2(KEYINPUT105), .ZN(n392) );
  NAND2_X1 U494 ( .A1(n526), .A2(n626), .ZN(n390) );
  NAND2_X1 U495 ( .A1(n392), .A2(n391), .ZN(n404) );
  NAND2_X1 U496 ( .A1(n364), .A2(n526), .ZN(n391) );
  NAND2_X1 U497 ( .A1(n413), .A2(KEYINPUT19), .ZN(n412) );
  NOR2_X2 U498 ( .A1(n623), .A2(n611), .ZN(n612) );
  NOR2_X1 U499 ( .A1(n615), .A2(n713), .ZN(n616) );
  NOR2_X1 U500 ( .A1(n661), .A2(n531), .ZN(n665) );
  NAND2_X1 U501 ( .A1(n593), .A2(n665), .ZN(n567) );
  INV_X1 U502 ( .A(n404), .ZN(n397) );
  NAND2_X1 U503 ( .A1(n404), .A2(n403), .ZN(n402) );
  AND2_X1 U504 ( .A1(n548), .A2(n508), .ZN(n403) );
  NOR2_X1 U505 ( .A1(n407), .A2(KEYINPUT19), .ZN(n406) );
  INV_X1 U506 ( .A(n419), .ZN(n407) );
  INV_X1 U507 ( .A(n413), .ZN(n408) );
  INV_X1 U508 ( .A(n411), .ZN(n410) );
  NAND2_X1 U509 ( .A1(n368), .A2(n419), .ZN(n573) );
  NAND2_X1 U510 ( .A1(n416), .A2(n414), .ZN(n413) );
  INV_X1 U511 ( .A(n418), .ZN(n415) );
  NAND2_X1 U512 ( .A1(n437), .A2(n433), .ZN(n418) );
  AND2_X1 U513 ( .A1(n686), .A2(n662), .ZN(n420) );
  INV_X1 U514 ( .A(KEYINPUT116), .ZN(n667) );
  XNOR2_X1 U515 ( .A(n667), .B(KEYINPUT50), .ZN(n668) );
  XNOR2_X1 U516 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U517 ( .A(n677), .B(KEYINPUT51), .ZN(n678) );
  INV_X1 U518 ( .A(KEYINPUT84), .ZN(n529) );
  XNOR2_X1 U519 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U520 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n693) );
  XNOR2_X1 U521 ( .A(n694), .B(n693), .ZN(n696) );
  XNOR2_X1 U522 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U523 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X2 U524 ( .A(G122), .B(G113), .ZN(n422) );
  XNOR2_X2 U525 ( .A(n422), .B(n421), .ZN(n450) );
  XNOR2_X2 U526 ( .A(G116), .B(G107), .ZN(n471) );
  XNOR2_X1 U527 ( .A(KEYINPUT16), .B(G110), .ZN(n423) );
  XNOR2_X1 U528 ( .A(n471), .B(n423), .ZN(n424) );
  NAND2_X1 U529 ( .A1(n780), .A2(G224), .ZN(n426) );
  XNOR2_X1 U530 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n425) );
  XNOR2_X1 U531 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X2 U532 ( .A(G143), .B(G128), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n427), .B(n470), .ZN(n428) );
  XNOR2_X1 U534 ( .A(n489), .B(n771), .ZN(n501) );
  XNOR2_X1 U535 ( .A(n455), .B(n429), .ZN(n430) );
  XNOR2_X1 U536 ( .A(n501), .B(n430), .ZN(n431) );
  XNOR2_X1 U537 ( .A(G902), .B(KEYINPUT15), .ZN(n639) );
  INV_X1 U538 ( .A(n639), .ZN(n433) );
  INV_X1 U539 ( .A(G902), .ZN(n518) );
  NAND2_X1 U540 ( .A1(n518), .A2(n434), .ZN(n438) );
  NAND2_X1 U541 ( .A1(n438), .A2(G210), .ZN(n436) );
  INV_X1 U542 ( .A(KEYINPUT89), .ZN(n435) );
  XNOR2_X1 U543 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U544 ( .A1(n438), .A2(G214), .ZN(n604) );
  INV_X1 U545 ( .A(n604), .ZN(n684) );
  XOR2_X1 U546 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n441) );
  XNOR2_X1 U547 ( .A(n441), .B(n440), .ZN(n695) );
  INV_X1 U548 ( .A(G952), .ZN(n697) );
  NOR2_X1 U549 ( .A1(G953), .A2(n697), .ZN(n563) );
  NAND2_X1 U550 ( .A1(n695), .A2(n563), .ZN(n445) );
  OR2_X1 U551 ( .A1(n780), .A2(G898), .ZN(n774) );
  NOR2_X1 U552 ( .A1(n518), .A2(n774), .ZN(n442) );
  NAND2_X1 U553 ( .A1(n442), .A2(n695), .ZN(n443) );
  XNOR2_X1 U554 ( .A(n443), .B(KEYINPUT90), .ZN(n444) );
  NAND2_X1 U555 ( .A1(n445), .A2(n444), .ZN(n446) );
  XOR2_X1 U556 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n448) );
  XNOR2_X1 U557 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U558 ( .A(n450), .B(n449), .ZN(n454) );
  XOR2_X1 U559 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n452) );
  XNOR2_X1 U560 ( .A(G131), .B(KEYINPUT96), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U562 ( .A(n454), .B(n453), .ZN(n461) );
  XNOR2_X1 U563 ( .A(n455), .B(KEYINPUT10), .ZN(n510) );
  NAND2_X1 U564 ( .A1(G214), .A2(n496), .ZN(n456) );
  XNOR2_X1 U565 ( .A(n456), .B(G140), .ZN(n458) );
  XNOR2_X1 U566 ( .A(G143), .B(KEYINPUT95), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U568 ( .A(n510), .B(n459), .ZN(n460) );
  XNOR2_X1 U569 ( .A(n461), .B(n460), .ZN(n731) );
  NAND2_X1 U570 ( .A1(n731), .A2(n518), .ZN(n464) );
  XNOR2_X1 U571 ( .A(KEYINPUT13), .B(G475), .ZN(n462) );
  XNOR2_X1 U572 ( .A(n462), .B(KEYINPUT99), .ZN(n463) );
  INV_X1 U573 ( .A(n551), .ZN(n477) );
  XOR2_X1 U574 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n466) );
  XNOR2_X1 U575 ( .A(G122), .B(KEYINPUT101), .ZN(n465) );
  XNOR2_X1 U576 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U577 ( .A(n467), .B(KEYINPUT102), .Z(n475) );
  NAND2_X1 U578 ( .A1(n511), .A2(G217), .ZN(n473) );
  XNOR2_X1 U579 ( .A(n485), .B(n471), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n475), .B(n474), .ZN(n742) );
  NAND2_X1 U581 ( .A1(n742), .A2(n518), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n476), .B(G478), .ZN(n555) );
  INV_X1 U583 ( .A(n555), .ZN(n552) );
  NAND2_X1 U584 ( .A1(n639), .A2(G234), .ZN(n478) );
  XNOR2_X1 U585 ( .A(n478), .B(KEYINPUT20), .ZN(n519) );
  NAND2_X1 U586 ( .A1(G221), .A2(n519), .ZN(n480) );
  INV_X1 U587 ( .A(KEYINPUT21), .ZN(n479) );
  XNOR2_X1 U588 ( .A(n480), .B(n479), .ZN(n662) );
  INV_X1 U589 ( .A(KEYINPUT72), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n482), .B(KEYINPUT22), .ZN(n483) );
  XNOR2_X2 U591 ( .A(n484), .B(n483), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n509), .B(n487), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n491), .B(n490), .ZN(n493) );
  NAND2_X1 U594 ( .A1(G227), .A2(n780), .ZN(n492) );
  XNOR2_X1 U595 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n494) );
  INV_X1 U596 ( .A(n666), .ZN(n626) );
  INV_X1 U597 ( .A(KEYINPUT105), .ZN(n495) );
  NAND2_X1 U598 ( .A1(n496), .A2(G210), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U600 ( .A(n499), .B(KEYINPUT5), .Z(n504) );
  XNOR2_X1 U601 ( .A(G113), .B(G116), .ZN(n500) );
  INV_X1 U602 ( .A(KEYINPUT92), .ZN(n505) );
  XNOR2_X1 U603 ( .A(n505), .B(G472), .ZN(n506) );
  INV_X1 U604 ( .A(n673), .ZN(n548) );
  INV_X1 U605 ( .A(KEYINPUT64), .ZN(n508) );
  XNOR2_X1 U606 ( .A(n510), .B(n509), .ZN(n777) );
  AND2_X1 U607 ( .A1(n511), .A2(G221), .ZN(n512) );
  XNOR2_X1 U608 ( .A(n777), .B(n512), .ZN(n517) );
  XNOR2_X1 U609 ( .A(n513), .B(G119), .ZN(n515) );
  XNOR2_X1 U610 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U611 ( .A(n517), .B(n516), .ZN(n739) );
  NAND2_X1 U612 ( .A1(n739), .A2(n518), .ZN(n524) );
  NAND2_X1 U613 ( .A1(G217), .A2(n519), .ZN(n522) );
  INV_X1 U614 ( .A(KEYINPUT77), .ZN(n520) );
  XNOR2_X1 U615 ( .A(n520), .B(KEYINPUT25), .ZN(n521) );
  XNOR2_X1 U616 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n666), .B(KEYINPUT86), .ZN(n614) );
  INV_X1 U618 ( .A(n358), .ZN(n527) );
  NAND2_X1 U619 ( .A1(n736), .A2(n659), .ZN(n530) );
  XNOR2_X1 U620 ( .A(n530), .B(n529), .ZN(n543) );
  INV_X1 U621 ( .A(n662), .ZN(n531) );
  INV_X1 U622 ( .A(n547), .ZN(n532) );
  NAND2_X1 U623 ( .A1(n605), .A2(n532), .ZN(n533) );
  XOR2_X1 U624 ( .A(n533), .B(KEYINPUT33), .Z(n700) );
  XOR2_X1 U625 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n535) );
  XNOR2_X1 U626 ( .A(n536), .B(n535), .ZN(n537) );
  AND2_X1 U627 ( .A1(n555), .A2(n551), .ZN(n591) );
  NAND2_X1 U628 ( .A1(n537), .A2(n591), .ZN(n541) );
  XNOR2_X1 U629 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n539) );
  INV_X1 U630 ( .A(KEYINPUT83), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X2 U632 ( .A(n541), .B(n540), .ZN(n789) );
  INV_X1 U633 ( .A(n789), .ZN(n542) );
  NAND2_X1 U634 ( .A1(n543), .A2(n542), .ZN(n545) );
  INV_X1 U635 ( .A(KEYINPUT44), .ZN(n544) );
  XNOR2_X1 U636 ( .A(n545), .B(n544), .ZN(n559) );
  NOR2_X1 U637 ( .A1(n356), .A2(n605), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n367), .A2(n546), .ZN(n747) );
  OR2_X1 U639 ( .A1(n548), .A2(n547), .ZN(n660) );
  OR2_X1 U640 ( .A1(n534), .A2(n660), .ZN(n549) );
  XNOR2_X1 U641 ( .A(n549), .B(KEYINPUT31), .ZN(n759) );
  OR2_X1 U642 ( .A1(n673), .A2(n567), .ZN(n550) );
  NOR2_X1 U643 ( .A1(n534), .A2(n550), .ZN(n753) );
  OR2_X1 U644 ( .A1(n759), .A2(n753), .ZN(n556) );
  INV_X1 U645 ( .A(KEYINPUT103), .ZN(n554) );
  XNOR2_X1 U646 ( .A(n760), .B(n554), .ZN(n621) );
  NAND2_X1 U647 ( .A1(n556), .A2(n683), .ZN(n557) );
  AND2_X1 U648 ( .A1(n747), .A2(n557), .ZN(n558) );
  NAND2_X1 U649 ( .A1(n559), .A2(n558), .ZN(n561) );
  INV_X1 U650 ( .A(KEYINPUT45), .ZN(n560) );
  XNOR2_X2 U651 ( .A(n561), .B(n560), .ZN(n637) );
  NOR2_X1 U652 ( .A1(G900), .A2(n780), .ZN(n562) );
  NAND2_X1 U653 ( .A1(n562), .A2(G902), .ZN(n565) );
  INV_X1 U654 ( .A(n563), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U656 ( .A(KEYINPUT30), .ZN(n570) );
  NAND2_X1 U657 ( .A1(n673), .A2(n604), .ZN(n569) );
  XNOR2_X1 U658 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U659 ( .A1(n572), .A2(n571), .ZN(n588) );
  INV_X1 U660 ( .A(KEYINPUT38), .ZN(n574) );
  XNOR2_X1 U661 ( .A(n573), .B(n574), .ZN(n685) );
  XNOR2_X1 U662 ( .A(n575), .B(KEYINPUT39), .ZN(n622) );
  NOR2_X1 U663 ( .A1(n622), .A2(n610), .ZN(n578) );
  XNOR2_X1 U664 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n576) );
  XOR2_X1 U665 ( .A(n576), .B(KEYINPUT40), .Z(n577) );
  XNOR2_X1 U666 ( .A(n578), .B(n577), .ZN(n788) );
  AND2_X1 U667 ( .A1(n662), .A2(n365), .ZN(n579) );
  AND2_X1 U668 ( .A1(n661), .A2(n579), .ZN(n606) );
  NAND2_X1 U669 ( .A1(n673), .A2(n606), .ZN(n581) );
  INV_X1 U670 ( .A(KEYINPUT28), .ZN(n580) );
  XNOR2_X1 U671 ( .A(n581), .B(n580), .ZN(n598) );
  AND2_X1 U672 ( .A1(n598), .A2(n593), .ZN(n584) );
  NAND2_X1 U673 ( .A1(n686), .A2(n604), .ZN(n582) );
  OR2_X1 U674 ( .A1(n685), .A2(n582), .ZN(n583) );
  XNOR2_X1 U675 ( .A(n583), .B(KEYINPUT41), .ZN(n680) );
  NAND2_X1 U676 ( .A1(n584), .A2(n680), .ZN(n586) );
  INV_X1 U677 ( .A(KEYINPUT42), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n586), .B(n585), .ZN(n654) );
  XNOR2_X1 U679 ( .A(n587), .B(KEYINPUT46), .ZN(n618) );
  NOR2_X1 U680 ( .A1(n588), .A2(n573), .ZN(n590) );
  INV_X1 U681 ( .A(KEYINPUT109), .ZN(n589) );
  XNOR2_X1 U682 ( .A(n590), .B(n589), .ZN(n592) );
  NAND2_X1 U683 ( .A1(n592), .A2(n591), .ZN(n758) );
  AND2_X1 U684 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U685 ( .A1(n598), .A2(n596), .ZN(n650) );
  INV_X1 U686 ( .A(KEYINPUT79), .ZN(n599) );
  OR2_X1 U687 ( .A1(n650), .A2(n599), .ZN(n595) );
  AND2_X1 U688 ( .A1(n758), .A2(n595), .ZN(n603) );
  AND2_X1 U689 ( .A1(n596), .A2(KEYINPUT47), .ZN(n597) );
  INV_X1 U690 ( .A(KEYINPUT47), .ZN(n600) );
  NOR2_X1 U691 ( .A1(KEYINPUT79), .A2(KEYINPUT47), .ZN(n601) );
  NAND2_X1 U692 ( .A1(n603), .A2(n602), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n605), .A2(n604), .ZN(n608) );
  INV_X1 U694 ( .A(n606), .ZN(n607) );
  OR2_X1 U695 ( .A1(n608), .A2(n607), .ZN(n623) );
  INV_X1 U696 ( .A(KEYINPUT107), .ZN(n609) );
  XNOR2_X1 U697 ( .A(n610), .B(n609), .ZN(n656) );
  OR2_X1 U698 ( .A1(n573), .A2(n656), .ZN(n611) );
  XNOR2_X1 U699 ( .A(n612), .B(KEYINPUT36), .ZN(n613) );
  AND2_X1 U700 ( .A1(n614), .A2(n613), .ZN(n713) );
  XNOR2_X1 U701 ( .A(n616), .B(KEYINPUT68), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U703 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n619) );
  XNOR2_X1 U704 ( .A(n620), .B(n619), .ZN(n631) );
  OR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n763) );
  OR2_X1 U706 ( .A1(n656), .A2(n623), .ZN(n625) );
  INV_X1 U707 ( .A(KEYINPUT108), .ZN(n624) );
  XNOR2_X1 U708 ( .A(n625), .B(n624), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U710 ( .A(n628), .B(KEYINPUT43), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n629), .A2(n573), .ZN(n655) );
  AND2_X1 U712 ( .A1(n763), .A2(n655), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n635) );
  INV_X1 U714 ( .A(n635), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n632), .A2(KEYINPUT2), .ZN(n633) );
  NOR2_X2 U716 ( .A1(n637), .A2(n633), .ZN(n634) );
  XNOR2_X2 U717 ( .A(n635), .B(KEYINPUT82), .ZN(n779) );
  XNOR2_X1 U718 ( .A(n779), .B(KEYINPUT74), .ZN(n636) );
  BUF_X2 U719 ( .A(n637), .Z(n706) );
  INV_X2 U720 ( .A(n706), .ZN(n764) );
  NAND2_X1 U721 ( .A1(n638), .A2(n764), .ZN(n642) );
  XNOR2_X1 U722 ( .A(n639), .B(KEYINPUT81), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n737), .A2(G472), .ZN(n646) );
  XOR2_X1 U726 ( .A(KEYINPUT62), .B(n644), .Z(n645) );
  XNOR2_X1 U727 ( .A(n646), .B(n645), .ZN(n647) );
  INV_X1 U728 ( .A(KEYINPUT63), .ZN(n648) );
  XNOR2_X1 U729 ( .A(n649), .B(n648), .ZN(G57) );
  NOR2_X1 U730 ( .A1(n650), .A2(n656), .ZN(n651) );
  XOR2_X1 U731 ( .A(G146), .B(n651), .Z(G48) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT29), .Z(n653) );
  NOR2_X1 U733 ( .A1(n650), .A2(n760), .ZN(n652) );
  XOR2_X1 U734 ( .A(n653), .B(n652), .Z(G30) );
  XOR2_X1 U735 ( .A(G137), .B(n654), .Z(G39) );
  XNOR2_X1 U736 ( .A(n655), .B(G140), .ZN(G42) );
  XNOR2_X1 U737 ( .A(G113), .B(KEYINPUT115), .ZN(n658) );
  INV_X1 U738 ( .A(n656), .ZN(n749) );
  NAND2_X1 U739 ( .A1(n759), .A2(n749), .ZN(n657) );
  XOR2_X1 U740 ( .A(n658), .B(n657), .Z(G15) );
  XNOR2_X1 U741 ( .A(n659), .B(G119), .ZN(G21) );
  INV_X1 U742 ( .A(n660), .ZN(n676) );
  INV_X1 U743 ( .A(n356), .ZN(n663) );
  NOR2_X1 U744 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U745 ( .A(KEYINPUT49), .B(n664), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U749 ( .A(KEYINPUT117), .B(n674), .Z(n675) );
  NOR2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n679) );
  INV_X1 U751 ( .A(KEYINPUT118), .ZN(n677) );
  INV_X1 U752 ( .A(n680), .ZN(n699) );
  NOR2_X1 U753 ( .A1(n681), .A2(n699), .ZN(n692) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n682) );
  NAND2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  AND2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n700), .A2(n690), .ZN(n691) );
  NOR2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U765 ( .A(KEYINPUT120), .B(n703), .Z(n704) );
  NOR2_X1 U766 ( .A1(n704), .A2(G953), .ZN(n710) );
  NOR2_X1 U767 ( .A1(n706), .A2(n779), .ZN(n707) );
  OR2_X1 U768 ( .A1(n707), .A2(KEYINPUT2), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n705), .A2(n708), .ZN(n709) );
  NAND2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U771 ( .A(KEYINPUT53), .B(n711), .Z(G75) );
  XNOR2_X1 U772 ( .A(G125), .B(KEYINPUT37), .ZN(n712) );
  XNOR2_X1 U773 ( .A(n713), .B(n712), .ZN(G27) );
  NAND2_X1 U774 ( .A1(n737), .A2(G210), .ZN(n718) );
  XNOR2_X1 U775 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n715) );
  XNOR2_X1 U776 ( .A(n715), .B(KEYINPUT55), .ZN(n716) );
  XNOR2_X1 U777 ( .A(n714), .B(n716), .ZN(n717) );
  XNOR2_X1 U778 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U779 ( .A(n720), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U780 ( .A1(n737), .A2(G469), .ZN(n727) );
  XNOR2_X1 U781 ( .A(n721), .B(KEYINPUT122), .ZN(n725) );
  XOR2_X1 U782 ( .A(KEYINPUT121), .B(KEYINPUT123), .Z(n723) );
  XNOR2_X1 U783 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n722) );
  XNOR2_X1 U784 ( .A(n723), .B(n722), .ZN(n724) );
  XNOR2_X1 U785 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U786 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U787 ( .A(n729), .B(KEYINPUT124), .ZN(G54) );
  XOR2_X1 U788 ( .A(KEYINPUT87), .B(KEYINPUT59), .Z(n730) );
  XNOR2_X1 U789 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U790 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U791 ( .A(n735), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U792 ( .A(n357), .B(G110), .ZN(G12) );
  NAND2_X1 U793 ( .A1(n741), .A2(G217), .ZN(n738) );
  XOR2_X1 U794 ( .A(n739), .B(n738), .Z(n740) );
  NOR2_X1 U795 ( .A1(n740), .A2(n745), .ZN(G66) );
  NAND2_X1 U796 ( .A1(n741), .A2(G478), .ZN(n744) );
  XNOR2_X1 U797 ( .A(n742), .B(KEYINPUT125), .ZN(n743) );
  XNOR2_X1 U798 ( .A(n744), .B(n743), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n746), .A2(n745), .ZN(G63) );
  XNOR2_X1 U800 ( .A(G101), .B(KEYINPUT112), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n748), .B(n747), .ZN(G3) );
  XNOR2_X1 U802 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n753), .A2(n749), .ZN(n750) );
  XOR2_X1 U804 ( .A(n751), .B(n750), .Z(n752) );
  XNOR2_X1 U805 ( .A(G104), .B(n752), .ZN(G6) );
  INV_X1 U806 ( .A(n753), .ZN(n754) );
  NOR2_X1 U807 ( .A1(n754), .A2(n760), .ZN(n756) );
  XNOR2_X1 U808 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n755) );
  XNOR2_X1 U809 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U810 ( .A(G107), .B(n757), .ZN(G9) );
  XNOR2_X1 U811 ( .A(G143), .B(n758), .ZN(G45) );
  INV_X1 U812 ( .A(n759), .ZN(n761) );
  NOR2_X1 U813 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U814 ( .A(G116), .B(n762), .Z(G18) );
  XNOR2_X1 U815 ( .A(G134), .B(n763), .ZN(G36) );
  NAND2_X1 U816 ( .A1(n764), .A2(n780), .ZN(n768) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n765) );
  XNOR2_X1 U818 ( .A(KEYINPUT61), .B(n765), .ZN(n766) );
  NAND2_X1 U819 ( .A1(n766), .A2(G898), .ZN(n767) );
  NAND2_X1 U820 ( .A1(n768), .A2(n767), .ZN(n776) );
  XNOR2_X1 U821 ( .A(G101), .B(KEYINPUT126), .ZN(n770) );
  XNOR2_X1 U822 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U823 ( .A(n769), .B(n772), .ZN(n773) );
  NAND2_X1 U824 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U825 ( .A(n776), .B(n775), .Z(G69) );
  XNOR2_X1 U826 ( .A(n777), .B(n778), .ZN(n782) );
  XNOR2_X1 U827 ( .A(n779), .B(n782), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n781), .A2(n780), .ZN(n786) );
  XNOR2_X1 U829 ( .A(G227), .B(n782), .ZN(n783) );
  NAND2_X1 U830 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U831 ( .A1(G953), .A2(n784), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U833 ( .A(KEYINPUT127), .B(n787), .Z(G72) );
  XOR2_X1 U834 ( .A(n788), .B(G131), .Z(G33) );
  XOR2_X1 U835 ( .A(G122), .B(n789), .Z(G24) );
endmodule

