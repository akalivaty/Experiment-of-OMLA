

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737;

  NOR2_X1 U366 ( .A1(n597), .A2(n596), .ZN(n697) );
  INV_X1 U367 ( .A(n699), .ZN(n696) );
  XNOR2_X2 U368 ( .A(n362), .B(KEYINPUT45), .ZN(n650) );
  XNOR2_X2 U369 ( .A(n571), .B(n570), .ZN(n649) );
  XNOR2_X2 U370 ( .A(n464), .B(n463), .ZN(n726) );
  XNOR2_X2 U371 ( .A(n655), .B(KEYINPUT66), .ZN(n358) );
  NOR2_X1 U372 ( .A1(n671), .A2(n723), .ZN(n672) );
  BUF_X1 U373 ( .A(n708), .Z(n718) );
  NOR2_X1 U374 ( .A1(n537), .A2(n736), .ZN(n364) );
  XNOR2_X1 U375 ( .A(n519), .B(n518), .ZN(n648) );
  AND2_X1 U376 ( .A1(n520), .A2(n517), .ZN(n519) );
  AND2_X1 U377 ( .A1(n566), .A2(n565), .ZN(n604) );
  NOR2_X1 U378 ( .A1(n525), .A2(n512), .ZN(n513) );
  OR2_X1 U379 ( .A1(n529), .A2(n511), .ZN(n699) );
  XNOR2_X1 U380 ( .A(n447), .B(n446), .ZN(n572) );
  INV_X1 U381 ( .A(KEYINPUT76), .ZN(n374) );
  XNOR2_X1 U382 ( .A(G122), .B(G104), .ZN(n410) );
  NOR2_X1 U383 ( .A1(n706), .A2(n350), .ZN(n349) );
  XNOR2_X1 U384 ( .A(n354), .B(n584), .ZN(n353) );
  NAND2_X1 U385 ( .A1(n351), .A2(n602), .ZN(n350) );
  XNOR2_X1 U386 ( .A(n407), .B(n406), .ZN(n725) );
  XNOR2_X1 U387 ( .A(G125), .B(G140), .ZN(n407) );
  OR2_X1 U388 ( .A1(n666), .A2(n368), .ZN(n367) );
  NAND2_X1 U389 ( .A1(n369), .A2(n443), .ZN(n368) );
  NAND2_X1 U390 ( .A1(n396), .A2(n653), .ZN(n370) );
  XNOR2_X1 U391 ( .A(n475), .B(n474), .ZN(n526) );
  XNOR2_X1 U392 ( .A(n725), .B(n408), .ZN(n440) );
  INV_X1 U393 ( .A(G146), .ZN(n408) );
  AND2_X1 U394 ( .A1(n352), .A2(n601), .ZN(n351) );
  INV_X1 U395 ( .A(n695), .ZN(n352) );
  AND2_X1 U396 ( .A1(n348), .A2(n593), .ZN(n594) );
  NAND2_X1 U397 ( .A1(n737), .A2(n649), .ZN(n354) );
  XNOR2_X1 U398 ( .A(G119), .B(G128), .ZN(n435) );
  XNOR2_X1 U399 ( .A(n440), .B(n361), .ZN(n360) );
  NAND2_X1 U400 ( .A1(n365), .A2(n371), .ZN(n589) );
  AND2_X1 U401 ( .A1(n367), .A2(n346), .ZN(n365) );
  INV_X1 U402 ( .A(n614), .ZN(n366) );
  OR2_X1 U403 ( .A1(n576), .A2(n586), .ZN(n578) );
  NOR2_X1 U404 ( .A1(G902), .A2(n720), .ZN(n447) );
  XNOR2_X1 U405 ( .A(KEYINPUT1), .B(KEYINPUT68), .ZN(n472) );
  NAND2_X1 U406 ( .A1(n356), .A2(n355), .ZN(n359) );
  INV_X1 U407 ( .A(n358), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n599), .B(KEYINPUT82), .ZN(n348) );
  NAND2_X1 U409 ( .A1(n699), .A2(n704), .ZN(n599) );
  INV_X1 U410 ( .A(KEYINPUT46), .ZN(n584) );
  XNOR2_X1 U411 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U412 ( .A(n344), .B(n411), .ZN(n361) );
  XOR2_X1 U413 ( .A(KEYINPUT92), .B(G143), .Z(n411) );
  XNOR2_X1 U414 ( .A(n453), .B(n452), .ZN(n464) );
  AND2_X1 U415 ( .A1(n572), .A2(n575), .ZN(n541) );
  INV_X1 U416 ( .A(G953), .ZN(n504) );
  BUF_X1 U417 ( .A(n650), .Z(n636) );
  XNOR2_X1 U418 ( .A(G116), .B(G122), .ZN(n416) );
  XNOR2_X1 U419 ( .A(G101), .B(G107), .ZN(n375) );
  XNOR2_X1 U420 ( .A(G143), .B(G128), .ZN(n383) );
  INV_X1 U421 ( .A(KEYINPUT65), .ZN(n382) );
  XNOR2_X1 U422 ( .A(n496), .B(KEYINPUT116), .ZN(n497) );
  NAND2_X1 U423 ( .A1(n345), .A2(n371), .ZN(n621) );
  NOR2_X1 U424 ( .A1(n526), .A2(n543), .ZN(n528) );
  XNOR2_X1 U425 ( .A(n415), .B(G475), .ZN(n529) );
  NOR2_X1 U426 ( .A1(n659), .A2(G902), .ZN(n414) );
  XNOR2_X1 U427 ( .A(n576), .B(KEYINPUT6), .ZN(n585) );
  INV_X1 U428 ( .A(KEYINPUT64), .ZN(n387) );
  XNOR2_X1 U429 ( .A(n442), .B(n441), .ZN(n720) );
  XNOR2_X1 U430 ( .A(n439), .B(n438), .ZN(n442) );
  OR2_X1 U431 ( .A1(n732), .A2(G952), .ZN(n680) );
  XNOR2_X1 U432 ( .A(n583), .B(n582), .ZN(n737) );
  AND2_X1 U433 ( .A1(n592), .A2(n618), .ZN(n706) );
  XNOR2_X1 U434 ( .A(n359), .B(n670), .ZN(n671) );
  XNOR2_X1 U435 ( .A(n589), .B(KEYINPUT19), .ZN(n595) );
  XOR2_X1 U436 ( .A(n410), .B(n409), .Z(n344) );
  AND2_X1 U437 ( .A1(n367), .A2(n370), .ZN(n345) );
  AND2_X1 U438 ( .A1(n370), .A2(n366), .ZN(n346) );
  AND2_X1 U439 ( .A1(n553), .A2(n684), .ZN(n347) );
  XNOR2_X1 U440 ( .A(n412), .B(n360), .ZN(n659) );
  NAND2_X1 U441 ( .A1(n547), .A2(n348), .ZN(n553) );
  NAND2_X1 U442 ( .A1(n353), .A2(n349), .ZN(n612) );
  NOR2_X2 U443 ( .A1(n358), .A2(n658), .ZN(n708) );
  NOR2_X1 U444 ( .A1(n658), .A2(n357), .ZN(n356) );
  INV_X1 U445 ( .A(G210), .ZN(n357) );
  NAND2_X1 U446 ( .A1(n363), .A2(n347), .ZN(n362) );
  XNOR2_X1 U447 ( .A(n364), .B(KEYINPUT44), .ZN(n363) );
  INV_X1 U448 ( .A(n396), .ZN(n369) );
  NAND2_X1 U449 ( .A1(n666), .A2(n396), .ZN(n371) );
  NAND2_X2 U450 ( .A1(n625), .A2(n624), .ZN(n730) );
  BUF_X1 U451 ( .A(n525), .Z(n543) );
  XNOR2_X1 U452 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n478) );
  XNOR2_X1 U453 ( .A(n479), .B(n478), .ZN(n483) );
  XNOR2_X1 U454 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n488) );
  INV_X1 U455 ( .A(KEYINPUT52), .ZN(n496) );
  XNOR2_X1 U456 ( .A(n498), .B(n497), .ZN(n499) );
  INV_X1 U457 ( .A(KEYINPUT33), .ZN(n474) );
  XNOR2_X1 U458 ( .A(n445), .B(KEYINPUT25), .ZN(n446) );
  INV_X1 U459 ( .A(KEYINPUT34), .ZN(n527) );
  XNOR2_X1 U460 ( .A(n709), .B(n710), .ZN(n711) );
  XNOR2_X1 U461 ( .A(n722), .B(n721), .ZN(n724) );
  XNOR2_X1 U462 ( .A(n632), .B(n631), .ZN(G75) );
  NAND2_X1 U463 ( .A1(G237), .A2(G234), .ZN(n373) );
  INV_X1 U464 ( .A(KEYINPUT14), .ZN(n372) );
  XNOR2_X1 U465 ( .A(n373), .B(n372), .ZN(n506) );
  XNOR2_X1 U466 ( .A(n374), .B(G110), .ZN(n376) );
  XNOR2_X1 U467 ( .A(n376), .B(n375), .ZN(n467) );
  XNOR2_X1 U468 ( .A(n410), .B(KEYINPUT16), .ZN(n377) );
  XNOR2_X1 U469 ( .A(n467), .B(n377), .ZN(n381) );
  XNOR2_X1 U470 ( .A(G119), .B(G116), .ZN(n378) );
  XNOR2_X1 U471 ( .A(n378), .B(KEYINPUT3), .ZN(n380) );
  XNOR2_X1 U472 ( .A(G113), .B(KEYINPUT73), .ZN(n379) );
  XNOR2_X1 U473 ( .A(n380), .B(n379), .ZN(n459) );
  XNOR2_X1 U474 ( .A(n381), .B(n459), .ZN(n634) );
  XNOR2_X1 U475 ( .A(n382), .B(KEYINPUT79), .ZN(n384) );
  XNOR2_X1 U476 ( .A(n384), .B(n383), .ZN(n425) );
  XNOR2_X1 U477 ( .A(KEYINPUT4), .B(G146), .ZN(n451) );
  XNOR2_X1 U478 ( .A(G125), .B(KEYINPUT87), .ZN(n385) );
  XNOR2_X1 U479 ( .A(n451), .B(n385), .ZN(n386) );
  XNOR2_X1 U480 ( .A(n425), .B(n386), .ZN(n392) );
  XNOR2_X2 U481 ( .A(n387), .B(G953), .ZN(n732) );
  NAND2_X1 U482 ( .A1(n732), .A2(G224), .ZN(n390) );
  XNOR2_X1 U483 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n388) );
  XNOR2_X1 U484 ( .A(n388), .B(KEYINPUT88), .ZN(n389) );
  XNOR2_X1 U485 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U486 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U487 ( .A(n634), .B(n393), .ZN(n666) );
  XNOR2_X1 U488 ( .A(G902), .B(KEYINPUT15), .ZN(n443) );
  INV_X1 U489 ( .A(n443), .ZN(n653) );
  NOR2_X1 U490 ( .A1(G902), .A2(G237), .ZN(n394) );
  XNOR2_X1 U491 ( .A(KEYINPUT75), .B(n394), .ZN(n397) );
  NAND2_X1 U492 ( .A1(n397), .A2(G210), .ZN(n395) );
  XNOR2_X1 U493 ( .A(n395), .B(KEYINPUT80), .ZN(n396) );
  XNOR2_X1 U494 ( .A(n621), .B(KEYINPUT38), .ZN(n567) );
  INV_X1 U495 ( .A(n567), .ZN(n431) );
  NAND2_X1 U496 ( .A1(n397), .A2(G214), .ZN(n398) );
  XNOR2_X1 U497 ( .A(n398), .B(KEYINPUT89), .ZN(n614) );
  NAND2_X1 U498 ( .A1(n431), .A2(n614), .ZN(n430) );
  XOR2_X1 U499 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n400) );
  NOR2_X1 U500 ( .A1(G953), .A2(G237), .ZN(n454) );
  NAND2_X1 U501 ( .A1(G214), .A2(n454), .ZN(n399) );
  XNOR2_X1 U502 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U503 ( .A(n401), .B(KEYINPUT91), .Z(n412) );
  INV_X1 U504 ( .A(KEYINPUT70), .ZN(n402) );
  NAND2_X1 U505 ( .A1(n402), .A2(KEYINPUT10), .ZN(n405) );
  INV_X1 U506 ( .A(KEYINPUT10), .ZN(n403) );
  NAND2_X1 U507 ( .A1(n403), .A2(KEYINPUT70), .ZN(n404) );
  NAND2_X1 U508 ( .A1(n405), .A2(n404), .ZN(n406) );
  XNOR2_X1 U509 ( .A(G113), .B(G131), .ZN(n409) );
  XNOR2_X1 U510 ( .A(KEYINPUT13), .B(KEYINPUT93), .ZN(n413) );
  XNOR2_X1 U511 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U512 ( .A(KEYINPUT7), .B(G107), .Z(n417) );
  XNOR2_X1 U513 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U514 ( .A(KEYINPUT96), .B(KEYINPUT9), .Z(n419) );
  XNOR2_X1 U515 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n418) );
  XNOR2_X1 U516 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U517 ( .A(n421), .B(n420), .Z(n424) );
  NAND2_X1 U518 ( .A1(n732), .A2(G234), .ZN(n422) );
  XOR2_X1 U519 ( .A(KEYINPUT8), .B(n422), .Z(n434) );
  NAND2_X1 U520 ( .A1(G217), .A2(n434), .ZN(n423) );
  XNOR2_X1 U521 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U522 ( .A(n425), .B(G134), .ZN(n453) );
  XNOR2_X1 U523 ( .A(n426), .B(n453), .ZN(n714) );
  INV_X1 U524 ( .A(G902), .ZN(n427) );
  NAND2_X1 U525 ( .A1(n714), .A2(n427), .ZN(n429) );
  INV_X1 U526 ( .A(G478), .ZN(n428) );
  XNOR2_X1 U527 ( .A(n429), .B(n428), .ZN(n530) );
  AND2_X1 U528 ( .A1(n529), .A2(n530), .ZN(n491) );
  NAND2_X1 U529 ( .A1(n430), .A2(n491), .ZN(n433) );
  NOR2_X1 U530 ( .A1(n431), .A2(n614), .ZN(n490) );
  INV_X1 U531 ( .A(n530), .ZN(n511) );
  NAND2_X1 U532 ( .A1(n529), .A2(n511), .ZN(n704) );
  NAND2_X1 U533 ( .A1(n490), .A2(n599), .ZN(n432) );
  NAND2_X1 U534 ( .A1(n433), .A2(n432), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n434), .A2(G221), .ZN(n439) );
  XOR2_X1 U536 ( .A(KEYINPUT24), .B(G110), .Z(n436) );
  XNOR2_X1 U537 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U538 ( .A(n437), .B(KEYINPUT23), .Z(n438) );
  XOR2_X1 U539 ( .A(G137), .B(KEYINPUT71), .Z(n463) );
  XNOR2_X1 U540 ( .A(n463), .B(n440), .ZN(n441) );
  NAND2_X1 U541 ( .A1(G234), .A2(n443), .ZN(n444) );
  XNOR2_X1 U542 ( .A(KEYINPUT20), .B(n444), .ZN(n448) );
  NAND2_X1 U543 ( .A1(G217), .A2(n448), .ZN(n445) );
  AND2_X1 U544 ( .A1(n448), .A2(G221), .ZN(n450) );
  INV_X1 U545 ( .A(KEYINPUT21), .ZN(n449) );
  XNOR2_X1 U546 ( .A(n450), .B(n449), .ZN(n510) );
  INV_X1 U547 ( .A(n510), .ZN(n575) );
  XNOR2_X1 U548 ( .A(n451), .B(G131), .ZN(n452) );
  NAND2_X1 U549 ( .A1(n454), .A2(G210), .ZN(n455) );
  XNOR2_X1 U550 ( .A(n455), .B(G137), .ZN(n457) );
  XNOR2_X1 U551 ( .A(G101), .B(KEYINPUT5), .ZN(n456) );
  XNOR2_X1 U552 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U553 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U554 ( .A(n464), .B(n460), .ZN(n677) );
  OR2_X1 U555 ( .A1(n677), .A2(G902), .ZN(n462) );
  INV_X1 U556 ( .A(G472), .ZN(n461) );
  XNOR2_X2 U557 ( .A(n462), .B(n461), .ZN(n576) );
  AND2_X1 U558 ( .A1(n541), .A2(n585), .ZN(n473) );
  XOR2_X1 U559 ( .A(G104), .B(G140), .Z(n466) );
  NAND2_X1 U560 ( .A1(G227), .A2(n732), .ZN(n465) );
  XNOR2_X1 U561 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U562 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U563 ( .A(n726), .B(n469), .ZN(n709) );
  NOR2_X1 U564 ( .A1(n709), .A2(G902), .ZN(n471) );
  INV_X1 U565 ( .A(G469), .ZN(n470) );
  XNOR2_X2 U566 ( .A(n471), .B(n470), .ZN(n540) );
  XNOR2_X2 U567 ( .A(n540), .B(n472), .ZN(n618) );
  NAND2_X1 U568 ( .A1(n473), .A2(n618), .ZN(n475) );
  INV_X1 U569 ( .A(n526), .ZN(n501) );
  NAND2_X1 U570 ( .A1(n476), .A2(n501), .ZN(n495) );
  INV_X1 U571 ( .A(n618), .ZN(n522) );
  INV_X1 U572 ( .A(n541), .ZN(n477) );
  NAND2_X1 U573 ( .A1(n522), .A2(n477), .ZN(n479) );
  INV_X1 U574 ( .A(n572), .ZN(n550) );
  NAND2_X1 U575 ( .A1(n550), .A2(n510), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n480), .B(KEYINPUT112), .ZN(n481) );
  XNOR2_X1 U577 ( .A(KEYINPUT49), .B(n481), .ZN(n482) );
  NOR2_X1 U578 ( .A1(n483), .A2(n482), .ZN(n484) );
  NAND2_X1 U579 ( .A1(n484), .A2(n576), .ZN(n485) );
  XNOR2_X1 U580 ( .A(n485), .B(KEYINPUT114), .ZN(n487) );
  AND2_X1 U581 ( .A1(n618), .A2(n541), .ZN(n486) );
  INV_X1 U582 ( .A(n576), .ZN(n542) );
  NAND2_X1 U583 ( .A1(n486), .A2(n542), .ZN(n538) );
  NAND2_X1 U584 ( .A1(n487), .A2(n538), .ZN(n489) );
  NAND2_X1 U585 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U586 ( .A(n492), .B(KEYINPUT41), .ZN(n581) );
  NAND2_X1 U587 ( .A1(n493), .A2(n581), .ZN(n494) );
  NAND2_X1 U588 ( .A1(n495), .A2(n494), .ZN(n498) );
  NOR2_X1 U589 ( .A1(n506), .A2(n499), .ZN(n500) );
  NAND2_X1 U590 ( .A1(n500), .A2(G952), .ZN(n503) );
  NAND2_X1 U591 ( .A1(n501), .A2(n581), .ZN(n502) );
  NAND2_X1 U592 ( .A1(n503), .A2(n502), .ZN(n628) );
  NOR2_X1 U593 ( .A1(G898), .A2(n504), .ZN(n635) );
  NAND2_X1 U594 ( .A1(n635), .A2(G902), .ZN(n505) );
  NAND2_X1 U595 ( .A1(n504), .A2(G952), .ZN(n559) );
  NAND2_X1 U596 ( .A1(n505), .A2(n559), .ZN(n507) );
  INV_X1 U597 ( .A(n506), .ZN(n561) );
  AND2_X1 U598 ( .A1(n507), .A2(n561), .ZN(n508) );
  NAND2_X1 U599 ( .A1(n595), .A2(n508), .ZN(n509) );
  XNOR2_X1 U600 ( .A(n509), .B(KEYINPUT0), .ZN(n525) );
  OR2_X1 U601 ( .A1(n511), .A2(n510), .ZN(n512) );
  NAND2_X1 U602 ( .A1(n513), .A2(n529), .ZN(n515) );
  INV_X1 U603 ( .A(KEYINPUT22), .ZN(n514) );
  XNOR2_X1 U604 ( .A(n515), .B(n514), .ZN(n520) );
  NAND2_X1 U605 ( .A1(n618), .A2(n550), .ZN(n516) );
  NOR2_X1 U606 ( .A1(n516), .A2(n585), .ZN(n517) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(KEYINPUT32), .Z(n518) );
  INV_X1 U608 ( .A(n520), .ZN(n548) );
  NOR2_X1 U609 ( .A1(n572), .A2(n542), .ZN(n521) );
  NAND2_X1 U610 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U611 ( .A1(n548), .A2(n523), .ZN(n646) );
  NOR2_X1 U612 ( .A1(n648), .A2(n646), .ZN(n524) );
  XNOR2_X1 U613 ( .A(n524), .B(KEYINPUT85), .ZN(n537) );
  XNOR2_X1 U614 ( .A(n528), .B(n527), .ZN(n534) );
  INV_X1 U615 ( .A(KEYINPUT97), .ZN(n532) );
  OR2_X1 U616 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U617 ( .A(n532), .B(n531), .ZN(n607) );
  XNOR2_X1 U618 ( .A(n607), .B(KEYINPUT78), .ZN(n533) );
  NOR2_X1 U619 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U620 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n535) );
  XNOR2_X1 U621 ( .A(n536), .B(n535), .ZN(n736) );
  NOR2_X1 U622 ( .A1(n538), .A2(n543), .ZN(n539) );
  XNOR2_X1 U623 ( .A(n539), .B(KEYINPUT31), .ZN(n703) );
  NAND2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n555) );
  NOR2_X1 U625 ( .A1(n555), .A2(n542), .ZN(n545) );
  INV_X1 U626 ( .A(n543), .ZN(n544) );
  NAND2_X1 U627 ( .A1(n545), .A2(n544), .ZN(n688) );
  NAND2_X1 U628 ( .A1(n703), .A2(n688), .ZN(n546) );
  XNOR2_X1 U629 ( .A(n546), .B(KEYINPUT90), .ZN(n547) );
  OR2_X1 U630 ( .A1(n548), .A2(n585), .ZN(n549) );
  XOR2_X1 U631 ( .A(KEYINPUT84), .B(n549), .Z(n552) );
  NOR2_X1 U632 ( .A1(n618), .A2(n550), .ZN(n551) );
  NAND2_X1 U633 ( .A1(n552), .A2(n551), .ZN(n684) );
  INV_X1 U634 ( .A(KEYINPUT100), .ZN(n554) );
  XNOR2_X1 U635 ( .A(n555), .B(n554), .ZN(n566) );
  OR2_X1 U636 ( .A1(n576), .A2(n614), .ZN(n557) );
  XNOR2_X1 U637 ( .A(KEYINPUT101), .B(KEYINPUT30), .ZN(n556) );
  XNOR2_X1 U638 ( .A(n557), .B(n556), .ZN(n564) );
  NOR2_X1 U639 ( .A1(n732), .A2(G900), .ZN(n558) );
  NAND2_X1 U640 ( .A1(G902), .A2(n558), .ZN(n560) );
  NAND2_X1 U641 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U642 ( .A1(n562), .A2(n561), .ZN(n573) );
  INV_X1 U643 ( .A(n573), .ZN(n563) );
  AND2_X1 U644 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U645 ( .A1(n604), .A2(n567), .ZN(n568) );
  XNOR2_X1 U646 ( .A(n568), .B(KEYINPUT39), .ZN(n623) );
  NAND2_X1 U647 ( .A1(n623), .A2(n696), .ZN(n571) );
  INV_X1 U648 ( .A(KEYINPUT103), .ZN(n569) );
  XNOR2_X1 U649 ( .A(n569), .B(KEYINPUT40), .ZN(n570) );
  NOR2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U651 ( .A1(n575), .A2(n574), .ZN(n586) );
  INV_X1 U652 ( .A(KEYINPUT28), .ZN(n577) );
  XNOR2_X1 U653 ( .A(n578), .B(n577), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n540), .A2(n579), .ZN(n597) );
  INV_X1 U655 ( .A(n597), .ZN(n580) );
  AND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X1 U657 ( .A(KEYINPUT42), .ZN(n582) );
  INV_X1 U658 ( .A(n585), .ZN(n587) );
  NOR2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n696), .A2(n588), .ZN(n613) );
  XNOR2_X1 U661 ( .A(KEYINPUT104), .B(n613), .ZN(n590) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT36), .ZN(n592) );
  INV_X1 U664 ( .A(KEYINPUT47), .ZN(n593) );
  XNOR2_X1 U665 ( .A(KEYINPUT74), .B(n594), .ZN(n598) );
  INV_X1 U666 ( .A(n595), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n598), .A2(n697), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n697), .A2(n599), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n600), .A2(KEYINPUT47), .ZN(n601) );
  INV_X1 U670 ( .A(n621), .ZN(n603) );
  NAND2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n606) );
  INV_X1 U672 ( .A(KEYINPUT102), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n606), .B(n605), .ZN(n609) );
  INV_X1 U674 ( .A(n607), .ZN(n608) );
  AND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(n695) );
  INV_X1 U676 ( .A(KEYINPUT72), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(KEYINPUT48), .ZN(n611) );
  XNOR2_X1 U678 ( .A(n612), .B(n611), .ZN(n625) );
  INV_X1 U679 ( .A(KEYINPUT98), .ZN(n616) );
  NOR2_X1 U680 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U681 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X1 U682 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U683 ( .A(n619), .B(KEYINPUT43), .ZN(n620) );
  XNOR2_X1 U684 ( .A(n620), .B(KEYINPUT99), .ZN(n622) );
  AND2_X1 U685 ( .A1(n622), .A2(n621), .ZN(n673) );
  INV_X1 U686 ( .A(n704), .ZN(n691) );
  AND2_X1 U687 ( .A1(n623), .A2(n691), .ZN(n633) );
  NOR2_X1 U688 ( .A1(n673), .A2(n633), .ZN(n624) );
  INV_X1 U689 ( .A(n730), .ZN(n626) );
  NAND2_X1 U690 ( .A1(n636), .A2(n626), .ZN(n657) );
  XNOR2_X1 U691 ( .A(n657), .B(KEYINPUT2), .ZN(n627) );
  NOR2_X1 U692 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U693 ( .A(n629), .B(KEYINPUT117), .ZN(n630) );
  NOR2_X1 U694 ( .A1(G953), .A2(n630), .ZN(n632) );
  XNOR2_X1 U695 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n631) );
  XOR2_X1 U696 ( .A(G134), .B(n633), .Z(G36) );
  NOR2_X1 U697 ( .A1(n634), .A2(n635), .ZN(n645) );
  INV_X1 U698 ( .A(n636), .ZN(n637) );
  NOR2_X1 U699 ( .A1(n637), .A2(G953), .ZN(n643) );
  NAND2_X1 U700 ( .A1(G224), .A2(G953), .ZN(n638) );
  XNOR2_X1 U701 ( .A(n638), .B(KEYINPUT124), .ZN(n639) );
  XNOR2_X1 U702 ( .A(KEYINPUT61), .B(n639), .ZN(n640) );
  NAND2_X1 U703 ( .A1(n640), .A2(G898), .ZN(n641) );
  XNOR2_X1 U704 ( .A(n641), .B(KEYINPUT125), .ZN(n642) );
  NOR2_X1 U705 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U706 ( .A(n645), .B(n644), .Z(G69) );
  XOR2_X1 U707 ( .A(G110), .B(n646), .Z(G12) );
  XNOR2_X1 U708 ( .A(G119), .B(KEYINPUT127), .ZN(n647) );
  XNOR2_X1 U709 ( .A(n648), .B(n647), .ZN(G21) );
  XNOR2_X1 U710 ( .A(n649), .B(G131), .ZN(G33) );
  XNOR2_X1 U711 ( .A(n730), .B(KEYINPUT77), .ZN(n651) );
  NAND2_X1 U712 ( .A1(n651), .A2(n650), .ZN(n652) );
  INV_X1 U713 ( .A(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U714 ( .A1(n652), .A2(n656), .ZN(n654) );
  NAND2_X1 U715 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U716 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U717 ( .A1(n708), .A2(G475), .ZN(n662) );
  XOR2_X1 U718 ( .A(KEYINPUT69), .B(KEYINPUT59), .Z(n660) );
  XNOR2_X1 U719 ( .A(n659), .B(n660), .ZN(n661) );
  XNOR2_X1 U720 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U721 ( .A1(n663), .A2(n680), .ZN(n665) );
  XOR2_X1 U722 ( .A(KEYINPUT120), .B(KEYINPUT60), .Z(n664) );
  XNOR2_X1 U723 ( .A(n665), .B(n664), .ZN(G60) );
  XOR2_X1 U724 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n668) );
  XNOR2_X1 U725 ( .A(KEYINPUT55), .B(KEYINPUT81), .ZN(n667) );
  XNOR2_X1 U726 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U727 ( .A(n666), .B(n669), .ZN(n670) );
  INV_X1 U728 ( .A(n680), .ZN(n723) );
  XNOR2_X1 U729 ( .A(n672), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U730 ( .A(n673), .B(G140), .Z(G42) );
  NAND2_X1 U731 ( .A1(n708), .A2(G472), .ZN(n679) );
  XNOR2_X1 U732 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n675) );
  XNOR2_X1 U733 ( .A(KEYINPUT62), .B(KEYINPUT86), .ZN(n674) );
  XNOR2_X1 U734 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U735 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U737 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U738 ( .A(KEYINPUT107), .B(KEYINPUT63), .Z(n682) );
  XNOR2_X1 U739 ( .A(n683), .B(n682), .ZN(G57) );
  XNOR2_X1 U740 ( .A(G101), .B(n684), .ZN(G3) );
  NOR2_X1 U741 ( .A1(n688), .A2(n699), .ZN(n685) );
  XOR2_X1 U742 ( .A(G104), .B(n685), .Z(G6) );
  XOR2_X1 U743 ( .A(KEYINPUT26), .B(KEYINPUT108), .Z(n687) );
  XNOR2_X1 U744 ( .A(G107), .B(KEYINPUT27), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n687), .B(n686), .ZN(n690) );
  NOR2_X1 U746 ( .A1(n688), .A2(n704), .ZN(n689) );
  XOR2_X1 U747 ( .A(n690), .B(n689), .Z(G9) );
  XOR2_X1 U748 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n693) );
  NAND2_X1 U749 ( .A1(n697), .A2(n691), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(n694) );
  XOR2_X1 U751 ( .A(G128), .B(n694), .Z(G30) );
  XOR2_X1 U752 ( .A(G143), .B(n695), .Z(G45) );
  NAND2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(G146), .ZN(G48) );
  NOR2_X1 U755 ( .A1(n699), .A2(n703), .ZN(n701) );
  XNOR2_X1 U756 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U758 ( .A(G113), .B(n702), .ZN(G15) );
  NOR2_X1 U759 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U760 ( .A(G116), .B(n705), .Z(G18) );
  XNOR2_X1 U761 ( .A(G125), .B(n706), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U763 ( .A1(n718), .A2(G469), .ZN(n712) );
  XOR2_X1 U764 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n710) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n723), .A2(n713), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n718), .A2(G478), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n714), .B(KEYINPUT121), .ZN(n715) );
  XNOR2_X1 U769 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U770 ( .A1(n723), .A2(n717), .ZN(G63) );
  NAND2_X1 U771 ( .A1(n718), .A2(G217), .ZN(n722) );
  XOR2_X1 U772 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n724), .A2(n723), .ZN(G66) );
  XNOR2_X1 U775 ( .A(n726), .B(n725), .ZN(n731) );
  XOR2_X1 U776 ( .A(G227), .B(n731), .Z(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U778 ( .A1(G953), .A2(n728), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n729), .B(KEYINPUT126), .ZN(n735) );
  XOR2_X1 U780 ( .A(n731), .B(n730), .Z(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n735), .A2(n734), .ZN(G72) );
  XOR2_X1 U783 ( .A(n736), .B(G122), .Z(G24) );
  XNOR2_X1 U784 ( .A(G137), .B(n737), .ZN(G39) );
endmodule

