

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770;

  NOR2_X2 U378 ( .A1(G953), .A2(G237), .ZN(n449) );
  INV_X1 U379 ( .A(G953), .ZN(n747) );
  NOR2_X1 U380 ( .A1(n673), .A2(n609), .ZN(n664) );
  NOR2_X2 U381 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X2 U382 ( .A(n756), .B(G146), .ZN(n496) );
  XNOR2_X2 U383 ( .A(n484), .B(n483), .ZN(n756) );
  NOR2_X2 U384 ( .A1(n746), .A2(n758), .ZN(n668) );
  NOR2_X1 U385 ( .A1(n611), .A2(n607), .ZN(n608) );
  NAND2_X1 U386 ( .A1(n407), .A2(n403), .ZN(n588) );
  NOR2_X1 U387 ( .A1(n646), .A2(n736), .ZN(n647) );
  NOR2_X1 U388 ( .A1(n639), .A2(n736), .ZN(n641) );
  NOR2_X1 U389 ( .A1(n630), .A2(n736), .ZN(n632) );
  AND2_X1 U390 ( .A1(n394), .A2(n363), .ZN(n392) );
  XNOR2_X1 U391 ( .A(n520), .B(KEYINPUT32), .ZN(n768) );
  XNOR2_X1 U392 ( .A(n369), .B(n564), .ZN(n618) );
  AND2_X1 U393 ( .A1(n410), .A2(n408), .ZN(n407) );
  NOR2_X2 U394 ( .A1(n673), .A2(n672), .ZN(n528) );
  OR2_X1 U395 ( .A1(n534), .A2(n376), .ZN(n374) );
  XNOR2_X1 U396 ( .A(n461), .B(n460), .ZN(n536) );
  AND2_X1 U397 ( .A1(n406), .A2(n404), .ZN(n403) );
  XNOR2_X1 U398 ( .A(n514), .B(n365), .ZN(n540) );
  XNOR2_X1 U399 ( .A(n496), .B(n489), .ZN(n718) );
  XNOR2_X1 U400 ( .A(n739), .B(n426), .ZN(n493) );
  XNOR2_X1 U401 ( .A(n427), .B(G116), .ZN(n465) );
  XNOR2_X1 U402 ( .A(n359), .B(n424), .ZN(n739) );
  INV_X1 U403 ( .A(G107), .ZN(n427) );
  INV_X2 U404 ( .A(G143), .ZN(n418) );
  XNOR2_X1 U405 ( .A(KEYINPUT72), .B(G110), .ZN(n485) );
  XNOR2_X1 U406 ( .A(G146), .B(G125), .ZN(n448) );
  XOR2_X1 U407 ( .A(G137), .B(G140), .Z(n498) );
  NOR2_X2 U408 ( .A1(n658), .A2(n661), .ZN(n695) );
  INV_X2 U409 ( .A(n537), .ZN(n661) );
  NAND2_X1 U410 ( .A1(n436), .A2(n432), .ZN(n415) );
  XNOR2_X1 U411 ( .A(n486), .B(n498), .ZN(n390) );
  NAND2_X1 U412 ( .A1(n413), .A2(n619), .ZN(n412) );
  NAND2_X1 U413 ( .A1(n588), .A2(KEYINPUT0), .ZN(n381) );
  NAND2_X1 U414 ( .A1(n379), .A2(n377), .ZN(n375) );
  NOR2_X1 U415 ( .A1(n378), .A2(KEYINPUT0), .ZN(n377) );
  INV_X1 U416 ( .A(n588), .ZN(n379) );
  INV_X1 U417 ( .A(n417), .ZN(n378) );
  NOR2_X1 U418 ( .A1(n613), .A2(n396), .ZN(n395) );
  NAND2_X1 U419 ( .A1(n604), .A2(KEYINPUT19), .ZN(n409) );
  XNOR2_X1 U420 ( .A(G116), .B(G137), .ZN(n494) );
  XNOR2_X1 U421 ( .A(n482), .B(G134), .ZN(n484) );
  XNOR2_X1 U422 ( .A(G110), .B(KEYINPUT24), .ZN(n502) );
  XNOR2_X1 U423 ( .A(n448), .B(KEYINPUT10), .ZN(n500) );
  XNOR2_X1 U424 ( .A(KEYINPUT66), .B(G131), .ZN(n482) );
  XNOR2_X1 U425 ( .A(n485), .B(n389), .ZN(n388) );
  XNOR2_X1 U426 ( .A(n427), .B(G104), .ZN(n389) );
  INV_X1 U427 ( .A(KEYINPUT64), .ZN(n425) );
  XNOR2_X1 U428 ( .A(G122), .B(G104), .ZN(n455) );
  NAND2_X1 U429 ( .A1(n405), .A2(n440), .ZN(n404) );
  INV_X1 U430 ( .A(n416), .ZN(n400) );
  INV_X1 U431 ( .A(KEYINPUT0), .ZN(n380) );
  INV_X1 U432 ( .A(n482), .ZN(n481) );
  NAND2_X1 U433 ( .A1(n562), .A2(n563), .ZN(n369) );
  NAND2_X1 U434 ( .A1(n606), .A2(n605), .ZN(n611) );
  NOR2_X1 U435 ( .A1(n602), .A2(n386), .ZN(n603) );
  INV_X1 U436 ( .A(KEYINPUT101), .ZN(n396) );
  AND2_X1 U437 ( .A1(n531), .A2(n540), .ZN(n560) );
  NAND2_X1 U438 ( .A1(n372), .A2(n375), .ZN(n480) );
  AND2_X1 U439 ( .A1(n373), .A2(n381), .ZN(n372) );
  NOR2_X1 U440 ( .A1(n374), .A2(n536), .ZN(n373) );
  INV_X1 U441 ( .A(G237), .ZN(n433) );
  XNOR2_X1 U442 ( .A(n500), .B(n499), .ZN(n757) );
  XOR2_X1 U443 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n451) );
  NAND2_X1 U444 ( .A1(n361), .A2(n567), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n496), .B(n382), .ZN(n636) );
  XNOR2_X1 U446 ( .A(n383), .B(n493), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n492), .B(n357), .ZN(n383) );
  XNOR2_X1 U448 ( .A(KEYINPUT68), .B(KEYINPUT3), .ZN(n424) );
  XNOR2_X1 U449 ( .A(n504), .B(n503), .ZN(n506) );
  XOR2_X1 U450 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n503) );
  XNOR2_X1 U451 ( .A(n502), .B(n501), .ZN(n504) );
  XNOR2_X1 U452 ( .A(G128), .B(G119), .ZN(n505) );
  XNOR2_X1 U453 ( .A(n390), .B(n388), .ZN(n488) );
  XNOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n421) );
  INV_X1 U455 ( .A(KEYINPUT74), .ZN(n625) );
  XNOR2_X1 U456 ( .A(n560), .B(n370), .ZN(n581) );
  INV_X1 U457 ( .A(KEYINPUT104), .ZN(n370) );
  XNOR2_X1 U458 ( .A(n513), .B(KEYINPUT25), .ZN(n365) );
  XNOR2_X1 U459 ( .A(G143), .B(G113), .ZN(n447) );
  AND2_X1 U460 ( .A1(n629), .A2(G953), .ZN(n736) );
  XNOR2_X1 U461 ( .A(n565), .B(KEYINPUT40), .ZN(n769) );
  NOR2_X1 U462 ( .A1(n364), .A2(n543), .ZN(n520) );
  XNOR2_X1 U463 ( .A(n385), .B(KEYINPUT76), .ZN(n364) );
  NOR2_X1 U464 ( .A1(n589), .A2(n588), .ZN(n655) );
  AND2_X2 U465 ( .A1(n392), .A2(n391), .ZN(n521) );
  XNOR2_X1 U466 ( .A(n521), .B(n371), .ZN(G12) );
  INV_X1 U467 ( .A(G110), .ZN(n371) );
  NOR2_X1 U468 ( .A1(n533), .A2(n532), .ZN(n356) );
  XOR2_X1 U469 ( .A(n495), .B(n494), .Z(n357) );
  NOR2_X1 U470 ( .A1(n543), .A2(n542), .ZN(n358) );
  XOR2_X1 U471 ( .A(G113), .B(G119), .Z(n359) );
  AND2_X1 U472 ( .A1(n367), .A2(n601), .ZN(n360) );
  OR2_X1 U473 ( .A1(n417), .A2(n380), .ZN(n361) );
  AND2_X1 U474 ( .A1(n381), .A2(n361), .ZN(n362) );
  AND2_X1 U475 ( .A1(n393), .A2(n515), .ZN(n363) );
  XNOR2_X1 U476 ( .A(n519), .B(KEYINPUT100), .ZN(n387) );
  NAND2_X1 U477 ( .A1(n366), .A2(KEYINPUT44), .ZN(n384) );
  NAND2_X1 U478 ( .A1(n767), .A2(n548), .ZN(n366) );
  AND2_X1 U479 ( .A1(n600), .A2(n368), .ZN(n367) );
  INV_X1 U480 ( .A(n664), .ZN(n368) );
  NOR2_X1 U481 ( .A1(n536), .A2(n534), .ZN(n693) );
  NAND2_X1 U482 ( .A1(n362), .A2(n375), .ZN(n533) );
  INV_X1 U483 ( .A(n539), .ZN(n386) );
  AND2_X2 U484 ( .A1(n528), .A2(n539), .ZN(n522) );
  NAND2_X1 U485 ( .A1(n545), .A2(n384), .ZN(n546) );
  XNOR2_X2 U486 ( .A(n527), .B(n526), .ZN(n767) );
  NOR2_X2 U487 ( .A1(n768), .A2(n521), .ZN(n548) );
  NAND2_X1 U488 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U489 ( .A(n543), .ZN(n397) );
  XNOR2_X2 U490 ( .A(n480), .B(KEYINPUT22), .ZN(n543) );
  NAND2_X1 U491 ( .A1(n543), .A2(n396), .ZN(n391) );
  NAND2_X1 U492 ( .A1(n613), .A2(n396), .ZN(n393) );
  NAND2_X1 U493 ( .A1(n397), .A2(n395), .ZN(n394) );
  INV_X1 U494 ( .A(n402), .ZN(n414) );
  NAND2_X1 U495 ( .A1(n416), .A2(n415), .ZN(n402) );
  NAND2_X1 U496 ( .A1(n398), .A2(n411), .ZN(n410) );
  NOR2_X1 U497 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X1 U498 ( .A1(n415), .A2(n440), .ZN(n399) );
  NAND2_X1 U499 ( .A1(n402), .A2(n401), .ZN(n408) );
  INV_X1 U500 ( .A(n409), .ZN(n401) );
  NAND2_X1 U501 ( .A1(n414), .A2(n411), .ZN(n615) );
  INV_X1 U502 ( .A(n604), .ZN(n405) );
  OR2_X1 U503 ( .A1(n411), .A2(n409), .ZN(n406) );
  OR2_X1 U504 ( .A1(n643), .A2(n412), .ZN(n411) );
  INV_X1 U505 ( .A(n436), .ZN(n413) );
  NAND2_X1 U506 ( .A1(n643), .A2(n436), .ZN(n416) );
  XNOR2_X2 U507 ( .A(n553), .B(KEYINPUT45), .ZN(n746) );
  NOR2_X2 U508 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U509 ( .A1(n446), .A2(n558), .ZN(n417) );
  INV_X1 U510 ( .A(KEYINPUT80), .ZN(n591) );
  INV_X1 U511 ( .A(KEYINPUT48), .ZN(n610) );
  INV_X1 U512 ( .A(KEYINPUT69), .ZN(n501) );
  AND2_X1 U513 ( .A1(n658), .A2(n604), .ZN(n605) );
  XNOR2_X1 U514 ( .A(n508), .B(n507), .ZN(n511) );
  INV_X1 U515 ( .A(n582), .ZN(n563) );
  XNOR2_X1 U516 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X2 U517 ( .A(n418), .B(G128), .ZN(n464) );
  INV_X1 U518 ( .A(KEYINPUT4), .ZN(n419) );
  XNOR2_X2 U519 ( .A(n464), .B(n419), .ZN(n483) );
  NAND2_X1 U520 ( .A1(n747), .A2(G224), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U522 ( .A(n448), .B(n422), .ZN(n423) );
  XNOR2_X1 U523 ( .A(n483), .B(n423), .ZN(n431) );
  XNOR2_X1 U524 ( .A(n425), .B(G101), .ZN(n486) );
  INV_X1 U525 ( .A(n486), .ZN(n426) );
  XNOR2_X1 U526 ( .A(n465), .B(n485), .ZN(n429) );
  XNOR2_X1 U527 ( .A(n455), .B(KEYINPUT16), .ZN(n428) );
  XNOR2_X1 U528 ( .A(n429), .B(n428), .ZN(n741) );
  XNOR2_X1 U529 ( .A(n493), .B(n741), .ZN(n430) );
  XNOR2_X1 U530 ( .A(n431), .B(n430), .ZN(n643) );
  XNOR2_X1 U531 ( .A(KEYINPUT15), .B(G902), .ZN(n619) );
  INV_X1 U532 ( .A(n619), .ZN(n432) );
  INV_X1 U533 ( .A(G902), .ZN(n497) );
  NAND2_X1 U534 ( .A1(n497), .A2(n433), .ZN(n437) );
  NAND2_X1 U535 ( .A1(n437), .A2(G210), .ZN(n435) );
  INV_X1 U536 ( .A(KEYINPUT88), .ZN(n434) );
  XNOR2_X1 U537 ( .A(n435), .B(n434), .ZN(n436) );
  NAND2_X1 U538 ( .A1(n437), .A2(G214), .ZN(n439) );
  INV_X1 U539 ( .A(KEYINPUT89), .ZN(n438) );
  XNOR2_X1 U540 ( .A(n439), .B(n438), .ZN(n604) );
  INV_X1 U541 ( .A(KEYINPUT19), .ZN(n440) );
  NOR2_X1 U542 ( .A1(G898), .A2(n747), .ZN(n441) );
  XNOR2_X1 U543 ( .A(KEYINPUT91), .B(n441), .ZN(n743) );
  NAND2_X1 U544 ( .A1(G237), .A2(G234), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n442), .B(KEYINPUT14), .ZN(n443) );
  NAND2_X1 U546 ( .A1(G902), .A2(n443), .ZN(n555) );
  OR2_X1 U547 ( .A1(n743), .A2(n555), .ZN(n446) );
  NAND2_X1 U548 ( .A1(G952), .A2(n443), .ZN(n707) );
  NOR2_X1 U549 ( .A1(G953), .A2(n707), .ZN(n445) );
  INV_X1 U550 ( .A(KEYINPUT90), .ZN(n444) );
  XNOR2_X1 U551 ( .A(n445), .B(n444), .ZN(n558) );
  XNOR2_X1 U552 ( .A(n447), .B(n481), .ZN(n459) );
  XOR2_X1 U553 ( .A(KEYINPUT73), .B(n449), .Z(n491) );
  NAND2_X1 U554 ( .A1(n491), .A2(G214), .ZN(n453) );
  XNOR2_X1 U555 ( .A(KEYINPUT96), .B(KEYINPUT11), .ZN(n450) );
  XNOR2_X1 U556 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U557 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U558 ( .A(n500), .B(n454), .Z(n457) );
  XOR2_X1 U559 ( .A(n455), .B(G140), .Z(n456) );
  XNOR2_X1 U560 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U561 ( .A(n459), .B(n458), .ZN(n728) );
  NOR2_X1 U562 ( .A1(G902), .A2(n728), .ZN(n461) );
  XNOR2_X1 U563 ( .A(KEYINPUT13), .B(G475), .ZN(n460) );
  XOR2_X1 U564 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n463) );
  XNOR2_X1 U565 ( .A(G122), .B(G134), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n463), .B(n462), .ZN(n469) );
  XOR2_X1 U567 ( .A(n465), .B(n464), .Z(n467) );
  XNOR2_X1 U568 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n466) );
  XNOR2_X1 U569 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U570 ( .A(n469), .B(n468), .Z(n472) );
  NAND2_X1 U571 ( .A1(G234), .A2(n747), .ZN(n470) );
  XOR2_X1 U572 ( .A(KEYINPUT8), .B(n470), .Z(n509) );
  NAND2_X1 U573 ( .A1(G217), .A2(n509), .ZN(n471) );
  XNOR2_X1 U574 ( .A(n472), .B(n471), .ZN(n627) );
  NOR2_X1 U575 ( .A1(n627), .A2(G902), .ZN(n473) );
  INV_X1 U576 ( .A(n473), .ZN(n474) );
  XNOR2_X1 U577 ( .A(G478), .B(n474), .ZN(n534) );
  XOR2_X1 U578 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n476) );
  NAND2_X1 U579 ( .A1(G234), .A2(n619), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n476), .B(n475), .ZN(n512) );
  NAND2_X1 U581 ( .A1(n512), .A2(G221), .ZN(n479) );
  INV_X1 U582 ( .A(KEYINPUT94), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n477), .B(KEYINPUT21), .ZN(n478) );
  XNOR2_X1 U584 ( .A(n479), .B(n478), .ZN(n567) );
  NAND2_X1 U585 ( .A1(G227), .A2(n747), .ZN(n487) );
  XNOR2_X1 U586 ( .A(n488), .B(n487), .ZN(n489) );
  NOR2_X2 U587 ( .A1(G902), .A2(n718), .ZN(n490) );
  XNOR2_X2 U588 ( .A(n490), .B(G469), .ZN(n572) );
  XNOR2_X2 U589 ( .A(n572), .B(KEYINPUT1), .ZN(n673) );
  INV_X1 U590 ( .A(n673), .ZN(n613) );
  AND2_X1 U591 ( .A1(n491), .A2(G210), .ZN(n492) );
  XOR2_X1 U592 ( .A(KEYINPUT71), .B(KEYINPUT5), .Z(n495) );
  NAND2_X1 U593 ( .A1(n636), .A2(n497), .ZN(n517) );
  XNOR2_X1 U594 ( .A(KEYINPUT95), .B(G472), .ZN(n516) );
  XNOR2_X1 U595 ( .A(n517), .B(n516), .ZN(n570) );
  INV_X1 U596 ( .A(n498), .ZN(n499) );
  INV_X1 U597 ( .A(n757), .ZN(n508) );
  XNOR2_X1 U598 ( .A(n506), .B(n505), .ZN(n507) );
  NAND2_X1 U599 ( .A1(G221), .A2(n509), .ZN(n510) );
  XNOR2_X1 U600 ( .A(n511), .B(n510), .ZN(n735) );
  NOR2_X1 U601 ( .A1(G902), .A2(n735), .ZN(n514) );
  NAND2_X1 U602 ( .A1(n512), .A2(G217), .ZN(n513) );
  INV_X1 U603 ( .A(n540), .ZN(n676) );
  AND2_X1 U604 ( .A1(n570), .A2(n676), .ZN(n515) );
  XOR2_X1 U605 ( .A(n517), .B(n516), .Z(n682) );
  INV_X1 U606 ( .A(KEYINPUT6), .ZN(n518) );
  XNOR2_X1 U607 ( .A(n682), .B(n518), .ZN(n539) );
  NOR2_X1 U608 ( .A1(n673), .A2(n540), .ZN(n519) );
  NAND2_X1 U609 ( .A1(n540), .A2(n567), .ZN(n672) );
  XNOR2_X2 U610 ( .A(n522), .B(KEYINPUT33), .ZN(n690) );
  NOR2_X1 U611 ( .A1(n690), .A2(n533), .ZN(n523) );
  XNOR2_X1 U612 ( .A(n523), .B(KEYINPUT34), .ZN(n525) );
  NAND2_X1 U613 ( .A1(n536), .A2(n534), .ZN(n583) );
  XNOR2_X1 U614 ( .A(n583), .B(KEYINPUT75), .ZN(n524) );
  NAND2_X1 U615 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U616 ( .A(KEYINPUT35), .ZN(n526) );
  INV_X1 U617 ( .A(n528), .ZN(n529) );
  OR2_X1 U618 ( .A1(n570), .A2(n529), .ZN(n684) );
  OR2_X1 U619 ( .A1(n684), .A2(n533), .ZN(n530) );
  XNOR2_X1 U620 ( .A(n530), .B(KEYINPUT31), .ZN(n662) );
  INV_X1 U621 ( .A(n567), .ZN(n675) );
  NOR2_X1 U622 ( .A1(n572), .A2(n675), .ZN(n531) );
  NAND2_X1 U623 ( .A1(n570), .A2(n560), .ZN(n532) );
  NOR2_X1 U624 ( .A1(n662), .A2(n356), .ZN(n538) );
  INV_X1 U625 ( .A(n534), .ZN(n535) );
  AND2_X1 U626 ( .A1(n536), .A2(n535), .ZN(n658) );
  OR2_X1 U627 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U628 ( .A(n695), .B(KEYINPUT81), .Z(n594) );
  NOR2_X1 U629 ( .A1(n538), .A2(n594), .ZN(n544) );
  AND2_X1 U630 ( .A1(n673), .A2(n540), .ZN(n541) );
  NAND2_X1 U631 ( .A1(n386), .A2(n541), .ZN(n542) );
  NOR2_X1 U632 ( .A1(n544), .A2(n358), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n546), .B(KEYINPUT84), .ZN(n552) );
  INV_X1 U634 ( .A(KEYINPUT44), .ZN(n547) );
  NAND2_X1 U635 ( .A1(n767), .A2(n547), .ZN(n550) );
  XNOR2_X1 U636 ( .A(n548), .B(KEYINPUT85), .ZN(n549) );
  NOR2_X1 U637 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U638 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n564) );
  NOR2_X1 U639 ( .A1(n405), .A2(n570), .ZN(n554) );
  XNOR2_X1 U640 ( .A(n554), .B(KEYINPUT30), .ZN(n559) );
  NOR2_X1 U641 ( .A1(G900), .A2(n555), .ZN(n556) );
  NAND2_X1 U642 ( .A1(G953), .A2(n556), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n558), .A2(n557), .ZN(n566) );
  NAND2_X1 U644 ( .A1(n559), .A2(n566), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n561) );
  XNOR2_X1 U646 ( .A(n615), .B(n561), .ZN(n691) );
  NOR2_X1 U647 ( .A1(n581), .A2(n691), .ZN(n562) );
  NAND2_X1 U648 ( .A1(n618), .A2(n658), .ZN(n565) );
  XOR2_X1 U649 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n578) );
  NAND2_X1 U650 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U651 ( .A(KEYINPUT67), .B(n568), .ZN(n569) );
  NAND2_X1 U652 ( .A1(n569), .A2(n676), .ZN(n602) );
  NOR2_X1 U653 ( .A1(n602), .A2(n570), .ZN(n571) );
  XNOR2_X1 U654 ( .A(n571), .B(KEYINPUT28), .ZN(n574) );
  INV_X1 U655 ( .A(n572), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n574), .A2(n573), .ZN(n589) );
  INV_X1 U657 ( .A(n589), .ZN(n576) );
  NOR2_X1 U658 ( .A1(n691), .A2(n405), .ZN(n697) );
  NAND2_X1 U659 ( .A1(n693), .A2(n697), .ZN(n575) );
  XNOR2_X1 U660 ( .A(n575), .B(KEYINPUT41), .ZN(n709) );
  NAND2_X1 U661 ( .A1(n576), .A2(n709), .ZN(n577) );
  XNOR2_X1 U662 ( .A(n578), .B(n577), .ZN(n770) );
  NAND2_X1 U663 ( .A1(n769), .A2(n770), .ZN(n580) );
  XOR2_X1 U664 ( .A(KEYINPUT46), .B(KEYINPUT82), .Z(n579) );
  XNOR2_X1 U665 ( .A(n580), .B(n579), .ZN(n601) );
  OR2_X1 U666 ( .A1(n582), .A2(n581), .ZN(n584) );
  NOR2_X1 U667 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U668 ( .A1(n585), .A2(n615), .ZN(n634) );
  NAND2_X1 U669 ( .A1(KEYINPUT47), .A2(n695), .ZN(n586) );
  NAND2_X1 U670 ( .A1(n634), .A2(n586), .ZN(n587) );
  XNOR2_X1 U671 ( .A(n587), .B(KEYINPUT78), .ZN(n599) );
  INV_X1 U672 ( .A(KEYINPUT47), .ZN(n590) );
  NOR2_X1 U673 ( .A1(n655), .A2(n590), .ZN(n592) );
  XNOR2_X1 U674 ( .A(n592), .B(n591), .ZN(n597) );
  XOR2_X1 U675 ( .A(KEYINPUT47), .B(KEYINPUT65), .Z(n593) );
  NOR2_X1 U676 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n655), .A2(n595), .ZN(n596) );
  NAND2_X1 U678 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U680 ( .A(n603), .B(KEYINPUT102), .ZN(n606) );
  INV_X1 U681 ( .A(n615), .ZN(n607) );
  XOR2_X1 U682 ( .A(n608), .B(KEYINPUT36), .Z(n609) );
  XNOR2_X1 U683 ( .A(n360), .B(n610), .ZN(n617) );
  XOR2_X1 U684 ( .A(KEYINPUT103), .B(n611), .Z(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT43), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n633) );
  NOR2_X2 U688 ( .A1(n617), .A2(n633), .ZN(n623) );
  NAND2_X1 U689 ( .A1(n618), .A2(n661), .ZN(n667) );
  NAND2_X1 U690 ( .A1(n623), .A2(n667), .ZN(n758) );
  NOR2_X1 U691 ( .A1(n668), .A2(KEYINPUT2), .ZN(n620) );
  NOR2_X2 U692 ( .A1(n620), .A2(n619), .ZN(n725) );
  NAND2_X1 U693 ( .A1(n667), .A2(KEYINPUT2), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT77), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X2 U696 ( .A1(n746), .A2(n624), .ZN(n626) );
  XNOR2_X2 U697 ( .A(n626), .B(n625), .ZN(n724) );
  AND2_X2 U698 ( .A1(n725), .A2(n724), .ZN(n733) );
  NAND2_X1 U699 ( .A1(n733), .A2(G478), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(n627), .ZN(n630) );
  INV_X1 U701 ( .A(G952), .ZN(n629) );
  INV_X1 U702 ( .A(KEYINPUT121), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(G63) );
  XOR2_X1 U704 ( .A(G140), .B(n633), .Z(G42) );
  XNOR2_X1 U705 ( .A(n634), .B(G143), .ZN(G45) );
  NAND2_X1 U706 ( .A1(n733), .A2(G472), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT86), .B(KEYINPUT62), .Z(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(G57) );
  NAND2_X1 U712 ( .A1(n733), .A2(G210), .ZN(n645) );
  XOR2_X1 U713 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U717 ( .A(G101), .B(n358), .Z(G3) );
  NAND2_X1 U718 ( .A1(n356), .A2(n658), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n648), .B(G104), .ZN(G6) );
  XNOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .ZN(n652) );
  XOR2_X1 U721 ( .A(KEYINPUT106), .B(KEYINPUT26), .Z(n650) );
  NAND2_X1 U722 ( .A1(n356), .A2(n661), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(G9) );
  XOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .Z(n654) );
  NAND2_X1 U726 ( .A1(n655), .A2(n661), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(G30) );
  XOR2_X1 U728 ( .A(G146), .B(KEYINPUT107), .Z(n657) );
  NAND2_X1 U729 ( .A1(n655), .A2(n658), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(G48) );
  NAND2_X1 U731 ( .A1(n662), .A2(n658), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT108), .ZN(n660) );
  XNOR2_X1 U733 ( .A(G113), .B(n660), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(G116), .ZN(G18) );
  XNOR2_X1 U736 ( .A(G125), .B(n664), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U738 ( .A(G134), .B(KEYINPUT109), .Z(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(G36) );
  INV_X1 U740 ( .A(n724), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT2), .B(KEYINPUT79), .Z(n669) );
  NOR2_X1 U742 ( .A1(n668), .A2(n669), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n715) );
  NAND2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U745 ( .A(KEYINPUT50), .B(n674), .ZN(n680) );
  XOR2_X1 U746 ( .A(KEYINPUT49), .B(KEYINPUT110), .Z(n678) );
  NAND2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n683), .B(KEYINPUT111), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n687) );
  XOR2_X1 U753 ( .A(KEYINPUT51), .B(KEYINPUT112), .Z(n686) );
  XNOR2_X1 U754 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n709), .A2(n688), .ZN(n689) );
  XNOR2_X1 U756 ( .A(KEYINPUT113), .B(n689), .ZN(n704) );
  NAND2_X1 U757 ( .A1(n691), .A2(n405), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U759 ( .A(n694), .B(KEYINPUT114), .ZN(n699) );
  INV_X1 U760 ( .A(n695), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U763 ( .A(KEYINPUT115), .B(n700), .ZN(n701) );
  NOR2_X1 U764 ( .A1(n690), .A2(n701), .ZN(n702) );
  XNOR2_X1 U765 ( .A(n702), .B(KEYINPUT116), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U767 ( .A(n705), .B(KEYINPUT52), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U769 ( .A(n708), .B(KEYINPUT117), .ZN(n712) );
  INV_X1 U770 ( .A(n690), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n713), .B(KEYINPUT118), .ZN(n714) );
  NOR2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n747), .A2(n716), .ZN(n717) );
  XOR2_X1 U776 ( .A(KEYINPUT53), .B(n717), .Z(G75) );
  NAND2_X1 U777 ( .A1(n733), .A2(G469), .ZN(n722) );
  XNOR2_X1 U778 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n718), .B(KEYINPUT57), .ZN(n719) );
  XNOR2_X1 U780 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U781 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U782 ( .A1(n736), .A2(n723), .ZN(G54) );
  AND2_X1 U783 ( .A1(n724), .A2(G475), .ZN(n726) );
  NAND2_X1 U784 ( .A1(n726), .A2(n725), .ZN(n730) );
  XOR2_X1 U785 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n727) );
  XNOR2_X1 U786 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n736), .A2(n731), .ZN(n732) );
  XNOR2_X1 U788 ( .A(KEYINPUT60), .B(n732), .ZN(G60) );
  NAND2_X1 U789 ( .A1(n733), .A2(G217), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n735), .B(n734), .ZN(n737) );
  XNOR2_X1 U791 ( .A(n738), .B(KEYINPUT122), .ZN(G66) );
  XNOR2_X1 U792 ( .A(n739), .B(KEYINPUT124), .ZN(n740) );
  XOR2_X1 U793 ( .A(n741), .B(n740), .Z(n742) );
  XNOR2_X1 U794 ( .A(G101), .B(n742), .ZN(n744) );
  NAND2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U796 ( .A(n745), .B(KEYINPUT125), .ZN(n755) );
  INV_X1 U797 ( .A(n746), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n748), .A2(n747), .ZN(n753) );
  XOR2_X1 U799 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n750) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U804 ( .A(n755), .B(n754), .ZN(G69) );
  XOR2_X1 U805 ( .A(n756), .B(n757), .Z(n762) );
  XOR2_X1 U806 ( .A(n758), .B(n762), .Z(n759) );
  XNOR2_X1 U807 ( .A(KEYINPUT126), .B(n759), .ZN(n760) );
  NOR2_X1 U808 ( .A1(G953), .A2(n760), .ZN(n761) );
  XNOR2_X1 U809 ( .A(n761), .B(KEYINPUT127), .ZN(n766) );
  XNOR2_X1 U810 ( .A(G227), .B(n762), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(G900), .ZN(n764) );
  NAND2_X1 U812 ( .A1(G953), .A2(n764), .ZN(n765) );
  NAND2_X1 U813 ( .A1(n766), .A2(n765), .ZN(G72) );
  XNOR2_X1 U814 ( .A(n767), .B(G122), .ZN(G24) );
  XOR2_X1 U815 ( .A(G119), .B(n768), .Z(G21) );
  XNOR2_X1 U816 ( .A(n769), .B(G131), .ZN(G33) );
  XNOR2_X1 U817 ( .A(G137), .B(n770), .ZN(G39) );
endmodule

