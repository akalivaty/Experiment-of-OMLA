

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U559 ( .A1(n953), .A2(n845), .ZN(n526) );
  XNOR2_X1 U560 ( .A(n704), .B(KEYINPUT99), .ZN(n705) );
  XNOR2_X1 U561 ( .A(n706), .B(n705), .ZN(n708) );
  INV_X1 U562 ( .A(KEYINPUT28), .ZN(n709) );
  NOR2_X1 U563 ( .A1(n831), .A2(n526), .ZN(n832) );
  XOR2_X1 U564 ( .A(G2443), .B(G2446), .Z(n528) );
  XNOR2_X1 U565 ( .A(G2427), .B(G2451), .ZN(n527) );
  XNOR2_X1 U566 ( .A(n528), .B(n527), .ZN(n534) );
  XOR2_X1 U567 ( .A(G2430), .B(G2454), .Z(n530) );
  XNOR2_X1 U568 ( .A(G1348), .B(G1341), .ZN(n529) );
  XNOR2_X1 U569 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U570 ( .A(G2435), .B(G2438), .Z(n531) );
  XNOR2_X1 U571 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U572 ( .A(n534), .B(n533), .Z(n535) );
  AND2_X1 U573 ( .A1(G14), .A2(n535), .ZN(G401) );
  INV_X1 U574 ( .A(G57), .ZN(G237) );
  INV_X1 U575 ( .A(G132), .ZN(G219) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n650) );
  XNOR2_X1 U577 ( .A(G651), .B(KEYINPUT67), .ZN(n538) );
  NOR2_X1 U578 ( .A1(n650), .A2(n538), .ZN(n656) );
  NAND2_X1 U579 ( .A1(G75), .A2(n656), .ZN(n537) );
  NOR2_X1 U580 ( .A1(G543), .A2(G651), .ZN(n658) );
  NAND2_X1 U581 ( .A1(G88), .A2(n658), .ZN(n536) );
  NAND2_X1 U582 ( .A1(n537), .A2(n536), .ZN(n544) );
  NOR2_X1 U583 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n539), .Z(n662) );
  NAND2_X1 U585 ( .A1(n662), .A2(G62), .ZN(n542) );
  NOR2_X1 U586 ( .A1(G651), .A2(n650), .ZN(n540) );
  XNOR2_X1 U587 ( .A(KEYINPUT64), .B(n540), .ZN(n659) );
  NAND2_X1 U588 ( .A1(G50), .A2(n659), .ZN(n541) );
  NAND2_X1 U589 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U590 ( .A1(n544), .A2(n543), .ZN(G166) );
  INV_X1 U591 ( .A(G2104), .ZN(n546) );
  NOR2_X1 U592 ( .A1(G2105), .A2(n546), .ZN(n905) );
  NAND2_X1 U593 ( .A1(n905), .A2(G102), .ZN(n545) );
  XNOR2_X1 U594 ( .A(n545), .B(KEYINPUT90), .ZN(n555) );
  INV_X1 U595 ( .A(G2105), .ZN(n547) );
  NOR2_X1 U596 ( .A1(n547), .A2(n546), .ZN(n910) );
  NAND2_X1 U597 ( .A1(G114), .A2(n910), .ZN(n549) );
  NOR2_X1 U598 ( .A1(G2104), .A2(n547), .ZN(n913) );
  NAND2_X1 U599 ( .A1(G126), .A2(n913), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n553) );
  NOR2_X1 U601 ( .A1(G2105), .A2(G2104), .ZN(n550) );
  XOR2_X2 U602 ( .A(KEYINPUT17), .B(n550), .Z(n906) );
  NAND2_X1 U603 ( .A1(G138), .A2(n906), .ZN(n551) );
  XNOR2_X1 U604 ( .A(KEYINPUT91), .B(n551), .ZN(n552) );
  NOR2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U607 ( .A(n556), .B(KEYINPUT92), .Z(G164) );
  NAND2_X1 U608 ( .A1(G89), .A2(n658), .ZN(n557) );
  XNOR2_X1 U609 ( .A(n557), .B(KEYINPUT76), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U611 ( .A1(G76), .A2(n656), .ZN(n559) );
  NAND2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U613 ( .A(n561), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U614 ( .A1(n662), .A2(G63), .ZN(n563) );
  NAND2_X1 U615 ( .A1(G51), .A2(n659), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U619 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G94), .A2(G452), .ZN(n568) );
  XNOR2_X1 U622 ( .A(n568), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U624 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n850) );
  NAND2_X1 U626 ( .A1(n850), .A2(G567), .ZN(n570) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U628 ( .A1(n659), .A2(G43), .ZN(n580) );
  NAND2_X1 U629 ( .A1(n662), .A2(G56), .ZN(n571) );
  XNOR2_X1 U630 ( .A(KEYINPUT14), .B(n571), .ZN(n577) );
  NAND2_X1 U631 ( .A1(n658), .A2(G81), .ZN(n572) );
  XNOR2_X1 U632 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G68), .A2(n656), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(n575), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U637 ( .A(KEYINPUT73), .B(n578), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n580), .A2(n579), .ZN(n615) );
  INV_X1 U639 ( .A(n615), .ZN(n994) );
  NAND2_X1 U640 ( .A1(n994), .A2(G860), .ZN(G153) );
  NAND2_X1 U641 ( .A1(n662), .A2(G64), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G52), .A2(n659), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G77), .A2(n656), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G90), .A2(n658), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT9), .B(n585), .Z(n586) );
  NOR2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U649 ( .A(KEYINPUT70), .B(n588), .ZN(G171) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(n662), .A2(G66), .ZN(n595) );
  NAND2_X1 U652 ( .A1(G79), .A2(n656), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G92), .A2(n658), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U655 ( .A1(n659), .A2(G54), .ZN(n591) );
  XOR2_X1 U656 ( .A(KEYINPUT74), .B(n591), .Z(n592) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U658 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n596), .Z(n995) );
  INV_X1 U660 ( .A(n995), .ZN(n631) );
  NOR2_X1 U661 ( .A1(n631), .A2(G868), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n597), .B(KEYINPUT75), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U665 ( .A1(n662), .A2(G65), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G53), .A2(n659), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U668 ( .A1(G78), .A2(n656), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G91), .A2(n658), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U671 ( .A1(n605), .A2(n604), .ZN(n711) );
  INV_X1 U672 ( .A(n711), .ZN(G299) );
  INV_X1 U673 ( .A(G868), .ZN(n612) );
  NOR2_X1 U674 ( .A1(G286), .A2(n612), .ZN(n607) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U677 ( .A(KEYINPUT77), .B(n608), .Z(G297) );
  INV_X1 U678 ( .A(G860), .ZN(n634) );
  NAND2_X1 U679 ( .A1(n634), .A2(G559), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n609), .A2(n631), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT16), .ZN(n611) );
  XNOR2_X1 U682 ( .A(KEYINPUT78), .B(n611), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G559), .A2(n612), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n631), .A2(n613), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n614), .B(KEYINPUT79), .ZN(n617) );
  NOR2_X1 U686 ( .A1(n615), .A2(G868), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G135), .A2(n906), .ZN(n626) );
  NAND2_X1 U689 ( .A1(G123), .A2(n913), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(KEYINPUT18), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G111), .A2(n910), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n619), .B(KEYINPUT80), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G99), .A2(n905), .ZN(n622) );
  XNOR2_X1 U695 ( .A(KEYINPUT81), .B(n622), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(KEYINPUT82), .ZN(n933) );
  XNOR2_X1 U699 ( .A(n933), .B(G2096), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT83), .ZN(n630) );
  INV_X1 U701 ( .A(G2100), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n630), .A2(n629), .ZN(G156) );
  NAND2_X1 U703 ( .A1(G559), .A2(n631), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT84), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n994), .B(n633), .ZN(n676) );
  NAND2_X1 U706 ( .A1(n634), .A2(n676), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n662), .A2(G67), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G55), .A2(n659), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U710 ( .A1(G80), .A2(n656), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G93), .A2(n658), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n679) );
  XOR2_X1 U714 ( .A(n641), .B(n679), .Z(G145) );
  NAND2_X1 U715 ( .A1(G47), .A2(n659), .ZN(n648) );
  NAND2_X1 U716 ( .A1(G72), .A2(n656), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G85), .A2(n658), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n662), .A2(G60), .ZN(n644) );
  XOR2_X1 U720 ( .A(KEYINPUT68), .B(n644), .Z(n645) );
  NOR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U723 ( .A(KEYINPUT69), .B(n649), .Z(G290) );
  NAND2_X1 U724 ( .A1(G87), .A2(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U727 ( .A1(n662), .A2(n653), .ZN(n655) );
  NAND2_X1 U728 ( .A1(G49), .A2(n659), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(G288) );
  NAND2_X1 U730 ( .A1(n656), .A2(G73), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(KEYINPUT2), .ZN(n667) );
  NAND2_X1 U732 ( .A1(G86), .A2(n658), .ZN(n661) );
  NAND2_X1 U733 ( .A1(G48), .A2(n659), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U735 ( .A1(G61), .A2(n662), .ZN(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT85), .B(n663), .ZN(n664) );
  NOR2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(G305) );
  XOR2_X1 U739 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n669) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U742 ( .A(n679), .B(n670), .Z(n671) );
  XNOR2_X1 U743 ( .A(G288), .B(n671), .ZN(n672) );
  XNOR2_X1 U744 ( .A(G290), .B(n672), .ZN(n674) );
  XNOR2_X1 U745 ( .A(G166), .B(n711), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U747 ( .A(n675), .B(G305), .ZN(n856) );
  XNOR2_X1 U748 ( .A(n856), .B(n676), .ZN(n677) );
  NAND2_X1 U749 ( .A1(n677), .A2(G868), .ZN(n678) );
  XOR2_X1 U750 ( .A(KEYINPUT89), .B(n678), .Z(n681) );
  OR2_X1 U751 ( .A1(n679), .A2(G868), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U759 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U762 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U763 ( .A1(G96), .A2(n688), .ZN(n854) );
  NAND2_X1 U764 ( .A1(n854), .A2(G2106), .ZN(n692) );
  NAND2_X1 U765 ( .A1(G120), .A2(G69), .ZN(n689) );
  NOR2_X1 U766 ( .A1(G237), .A2(n689), .ZN(n690) );
  NAND2_X1 U767 ( .A1(G108), .A2(n690), .ZN(n855) );
  NAND2_X1 U768 ( .A1(n855), .A2(G567), .ZN(n691) );
  NAND2_X1 U769 ( .A1(n692), .A2(n691), .ZN(n932) );
  NAND2_X1 U770 ( .A1(G483), .A2(G661), .ZN(n693) );
  NOR2_X1 U771 ( .A1(n932), .A2(n693), .ZN(n853) );
  NAND2_X1 U772 ( .A1(n853), .A2(G36), .ZN(G176) );
  NAND2_X1 U773 ( .A1(G113), .A2(n910), .ZN(n695) );
  NAND2_X1 U774 ( .A1(G125), .A2(n913), .ZN(n694) );
  NAND2_X1 U775 ( .A1(n695), .A2(n694), .ZN(n702) );
  NAND2_X1 U776 ( .A1(G101), .A2(n905), .ZN(n696) );
  XNOR2_X1 U777 ( .A(n696), .B(KEYINPUT65), .ZN(n697) );
  XNOR2_X1 U778 ( .A(KEYINPUT23), .B(n697), .ZN(n700) );
  NAND2_X1 U779 ( .A1(G137), .A2(n906), .ZN(n698) );
  XNOR2_X1 U780 ( .A(n698), .B(KEYINPUT66), .ZN(n699) );
  NAND2_X1 U781 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U782 ( .A1(n702), .A2(n701), .ZN(G160) );
  INV_X1 U783 ( .A(G166), .ZN(G303) );
  INV_X1 U784 ( .A(KEYINPUT103), .ZN(n772) );
  NOR2_X1 U785 ( .A1(G1384), .A2(G164), .ZN(n799) );
  NAND2_X1 U786 ( .A1(G160), .A2(G40), .ZN(n798) );
  INV_X1 U787 ( .A(n798), .ZN(n703) );
  NAND2_X1 U788 ( .A1(n799), .A2(n703), .ZN(n745) );
  NAND2_X1 U789 ( .A1(G8), .A2(n745), .ZN(n794) );
  INV_X1 U790 ( .A(n745), .ZN(n717) );
  NAND2_X1 U791 ( .A1(G2072), .A2(n717), .ZN(n706) );
  INV_X1 U792 ( .A(KEYINPUT27), .ZN(n704) );
  INV_X1 U793 ( .A(G1956), .ZN(n1006) );
  NOR2_X1 U794 ( .A1(n717), .A2(n1006), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U796 ( .A1(n712), .A2(n711), .ZN(n710) );
  XNOR2_X1 U797 ( .A(n710), .B(n709), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n727) );
  INV_X1 U799 ( .A(G1996), .ZN(n960) );
  NOR2_X1 U800 ( .A1(n745), .A2(n960), .ZN(n714) );
  XOR2_X1 U801 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n713) );
  XNOR2_X1 U802 ( .A(n714), .B(n713), .ZN(n716) );
  NAND2_X1 U803 ( .A1(n745), .A2(G1341), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n722) );
  NAND2_X1 U805 ( .A1(G1348), .A2(n745), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n717), .A2(G2067), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U808 ( .A1(n995), .A2(n723), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n994), .A2(n720), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n725) );
  NOR2_X1 U811 ( .A1(n723), .A2(n995), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U814 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U815 ( .A(KEYINPUT29), .B(n730), .Z(n734) );
  INV_X1 U816 ( .A(G1961), .ZN(n1025) );
  NAND2_X1 U817 ( .A1(n745), .A2(n1025), .ZN(n732) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n967) );
  NAND2_X1 U819 ( .A1(n717), .A2(n967), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n741) );
  NAND2_X1 U821 ( .A1(G171), .A2(n741), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n761) );
  INV_X1 U823 ( .A(G8), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n750), .A2(G1966), .ZN(n735) );
  AND2_X1 U825 ( .A1(n735), .A2(n745), .ZN(n736) );
  XOR2_X1 U826 ( .A(KEYINPUT98), .B(n736), .Z(n763) );
  NOR2_X1 U827 ( .A1(G2084), .A2(n745), .ZN(n758) );
  NOR2_X1 U828 ( .A1(n750), .A2(n758), .ZN(n737) );
  AND2_X1 U829 ( .A1(n763), .A2(n737), .ZN(n739) );
  XNOR2_X1 U830 ( .A(KEYINPUT30), .B(KEYINPUT101), .ZN(n738) );
  XNOR2_X1 U831 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U832 ( .A1(G168), .A2(n740), .ZN(n743) );
  NOR2_X1 U833 ( .A1(G171), .A2(n741), .ZN(n742) );
  NOR2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U835 ( .A(KEYINPUT31), .B(n744), .Z(n760) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n794), .ZN(n747) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n745), .ZN(n746) );
  NOR2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n748), .A2(G303), .ZN(n749) );
  OR2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n752) );
  AND2_X1 U841 ( .A1(n760), .A2(n752), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n761), .A2(n751), .ZN(n756) );
  INV_X1 U843 ( .A(n752), .ZN(n754) );
  AND2_X1 U844 ( .A1(G286), .A2(G8), .ZN(n753) );
  OR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n757), .B(KEYINPUT32), .ZN(n767) );
  NAND2_X1 U848 ( .A1(G8), .A2(n758), .ZN(n759) );
  XOR2_X1 U849 ( .A(KEYINPUT97), .B(n759), .Z(n765) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n777) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n768) );
  NAND2_X1 U855 ( .A1(G8), .A2(n768), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n777), .A2(n769), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n794), .A2(n770), .ZN(n771) );
  XNOR2_X1 U858 ( .A(n772), .B(n771), .ZN(n791) );
  NOR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n987) );
  NOR2_X1 U860 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n987), .A2(n773), .ZN(n775) );
  INV_X1 U862 ( .A(KEYINPUT33), .ZN(n774) );
  AND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n781) );
  INV_X1 U865 ( .A(KEYINPUT102), .ZN(n782) );
  NOR2_X1 U866 ( .A1(n794), .A2(n782), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n988) );
  AND2_X1 U868 ( .A1(n778), .A2(n988), .ZN(n779) );
  OR2_X1 U869 ( .A1(KEYINPUT33), .A2(n779), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n788) );
  NAND2_X1 U871 ( .A1(n782), .A2(n987), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n987), .A2(KEYINPUT33), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n783), .A2(KEYINPUT102), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U875 ( .A1(n794), .A2(n786), .ZN(n787) );
  NOR2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U877 ( .A(G1981), .B(G305), .Z(n982) );
  NAND2_X1 U878 ( .A1(n789), .A2(n982), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n796) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XOR2_X1 U881 ( .A(n792), .B(KEYINPUT24), .Z(n793) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n797) );
  INV_X1 U884 ( .A(n797), .ZN(n833) );
  NOR2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n845) );
  NOR2_X1 U886 ( .A1(G1986), .A2(G290), .ZN(n834) );
  INV_X1 U887 ( .A(n834), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n991) );
  NAND2_X1 U890 ( .A1(n845), .A2(n991), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n802), .B(KEYINPUT93), .ZN(n831) );
  NAND2_X1 U892 ( .A1(G141), .A2(n906), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G117), .A2(n910), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n905), .A2(G105), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(n805), .Z(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n913), .A2(G129), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n899) );
  NAND2_X1 U900 ( .A1(G1996), .A2(n899), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n810), .B(KEYINPUT96), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G95), .A2(n905), .ZN(n812) );
  NAND2_X1 U903 ( .A1(G131), .A2(n906), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n816) );
  NAND2_X1 U905 ( .A1(G107), .A2(n910), .ZN(n814) );
  NAND2_X1 U906 ( .A1(G119), .A2(n913), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n900) );
  NAND2_X1 U909 ( .A1(G1991), .A2(n900), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n836) );
  INV_X1 U911 ( .A(n836), .ZN(n830) );
  NAND2_X1 U912 ( .A1(n910), .A2(G116), .ZN(n819) );
  XOR2_X1 U913 ( .A(KEYINPUT95), .B(n819), .Z(n821) );
  NAND2_X1 U914 ( .A1(n913), .A2(G128), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n822), .B(KEYINPUT35), .ZN(n827) );
  NAND2_X1 U917 ( .A1(G104), .A2(n905), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G140), .A2(n906), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U920 ( .A(KEYINPUT34), .B(n825), .Z(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U922 ( .A(n828), .B(KEYINPUT36), .Z(n921) );
  XOR2_X1 U923 ( .A(G2067), .B(KEYINPUT37), .Z(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT94), .B(n829), .Z(n842) );
  OR2_X1 U925 ( .A1(n921), .A2(n842), .ZN(n839) );
  NAND2_X1 U926 ( .A1(n830), .A2(n839), .ZN(n953) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n848) );
  NOR2_X1 U928 ( .A1(G1996), .A2(n899), .ZN(n948) );
  NOR2_X1 U929 ( .A1(G1991), .A2(n900), .ZN(n936) );
  NOR2_X1 U930 ( .A1(n834), .A2(n936), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U932 ( .A1(n948), .A2(n837), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n838), .B(KEYINPUT39), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n841), .B(KEYINPUT104), .ZN(n843) );
  NAND2_X1 U936 ( .A1(n842), .A2(n921), .ZN(n937) );
  NAND2_X1 U937 ( .A1(n843), .A2(n937), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U939 ( .A(KEYINPUT105), .B(n846), .Z(n847) );
  NAND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U941 ( .A(KEYINPUT40), .B(n849), .ZN(G329) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U946 ( .A1(n853), .A2(n852), .ZN(G188) );
  XOR2_X1 U947 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  NOR2_X1 U951 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U953 ( .A(n995), .B(n856), .ZN(n858) );
  XNOR2_X1 U954 ( .A(G301), .B(n994), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U956 ( .A(G286), .B(n859), .Z(n860) );
  NOR2_X1 U957 ( .A1(G37), .A2(n860), .ZN(G397) );
  XOR2_X1 U958 ( .A(KEYINPUT109), .B(G1991), .Z(n862) );
  XNOR2_X1 U959 ( .A(G1976), .B(G1996), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n863), .B(KEYINPUT110), .Z(n865) );
  XNOR2_X1 U962 ( .A(G1971), .B(G1961), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U964 ( .A(G1986), .B(G1956), .Z(n867) );
  XNOR2_X1 U965 ( .A(G1981), .B(G1966), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U968 ( .A(G2474), .B(KEYINPUT41), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(G229) );
  XOR2_X1 U970 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n873) );
  XNOR2_X1 U971 ( .A(G2678), .B(KEYINPUT43), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n877) );
  XOR2_X1 U973 ( .A(KEYINPUT42), .B(G2090), .Z(n875) );
  XNOR2_X1 U974 ( .A(G2072), .B(G2067), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U976 ( .A(n877), .B(n876), .Z(n879) );
  XNOR2_X1 U977 ( .A(G2096), .B(G2100), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n881) );
  XOR2_X1 U979 ( .A(G2078), .B(G2084), .Z(n880) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(G227) );
  NAND2_X1 U981 ( .A1(G124), .A2(n913), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n882), .B(KEYINPUT44), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G136), .A2(n906), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT111), .B(n883), .Z(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G100), .A2(n905), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G112), .A2(n910), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(G162) );
  NAND2_X1 U990 ( .A1(G103), .A2(n905), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G139), .A2(n906), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n897) );
  NAND2_X1 U993 ( .A1(n913), .A2(G127), .ZN(n892) );
  XOR2_X1 U994 ( .A(KEYINPUT113), .B(n892), .Z(n894) );
  NAND2_X1 U995 ( .A1(n910), .A2(G115), .ZN(n893) );
  NAND2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n939) );
  XOR2_X1 U999 ( .A(G160), .B(G162), .Z(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n900), .B(KEYINPUT114), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1004 ( .A(n904), .B(n903), .Z(n919) );
  NAND2_X1 U1005 ( .A1(G106), .A2(n905), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n906), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n909), .B(KEYINPUT45), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(G118), .A2(n910), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n916) );
  NAND2_X1 U1011 ( .A1(n913), .A2(G130), .ZN(n914) );
  XOR2_X1 U1012 ( .A(KEYINPUT112), .B(n914), .Z(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n933), .B(n917), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n939), .B(n920), .ZN(n923) );
  XOR2_X1 U1017 ( .A(G164), .B(n921), .Z(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n924), .ZN(n925) );
  XOR2_X1 U1020 ( .A(KEYINPUT115), .B(n925), .Z(G395) );
  NOR2_X1 U1021 ( .A1(G401), .A2(n932), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(G229), .A2(G227), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT49), .B(n926), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G397), .A2(n927), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n930), .A2(G395), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1028 ( .A(G308), .ZN(G225) );
  INV_X1 U1029 ( .A(n932), .ZN(G319) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n945) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n942) );
  XOR2_X1 U1036 ( .A(n939), .B(KEYINPUT118), .Z(n940) );
  XNOR2_X1 U1037 ( .A(G2072), .B(n940), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n943), .Z(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G162), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(n946), .B(KEYINPUT117), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1044 ( .A(KEYINPUT51), .B(n949), .Z(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1047 ( .A(KEYINPUT52), .B(n954), .Z(n955) );
  NOR2_X1 U1048 ( .A1(KEYINPUT55), .A2(n955), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT119), .B(n956), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G29), .ZN(n1038) );
  XNOR2_X1 U1051 ( .A(G2072), .B(G33), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G1991), .B(G25), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(G32), .B(n960), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n961), .A2(G28), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT120), .B(G2067), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G26), .B(n962), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1060 ( .A(G27), .B(n967), .Z(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n970), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n971), .B(KEYINPUT121), .ZN(n975) );
  XOR2_X1 U1064 ( .A(G34), .B(KEYINPUT122), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G2084), .B(KEYINPUT54), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G35), .B(G2090), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT55), .B(n978), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n979), .B(KEYINPUT123), .ZN(n980) );
  OR2_X1 U1072 ( .A1(G29), .A2(n980), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n981), .ZN(n1036) );
  XNOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .ZN(n1005) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G168), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(n984), .B(KEYINPUT57), .ZN(n1003) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G166), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n985), .B(KEYINPUT124), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G299), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(n994), .B(G1341), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(n995), .B(G1348), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G301), .B(G1961), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1034) );
  INV_X1 U1093 ( .A(G16), .ZN(n1032) );
  XNOR2_X1 U1094 ( .A(G20), .B(n1006), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT59), .B(G1348), .Z(n1011) );
  XNOR2_X1 U1100 ( .A(G4), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(n1015), .B(n1014), .ZN(n1024) );
  XOR2_X1 U1104 ( .A(G1971), .B(G22), .Z(n1018) );
  XOR2_X1 U1105 ( .A(G23), .B(KEYINPUT126), .Z(n1016) );
  XNOR2_X1 U1106 ( .A(n1016), .B(G1976), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(KEYINPUT127), .B(G1986), .Z(n1019) );
  XNOR2_X1 U1109 ( .A(G24), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(G1966), .B(G21), .Z(n1027) );
  XNOR2_X1 U1114 ( .A(n1025), .B(G5), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1039), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

