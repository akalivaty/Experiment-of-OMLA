//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT69), .B(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n468), .B2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n474), .A3(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(KEYINPUT70), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G137), .A3(new_n461), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n467), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n465), .B1(new_n478), .B2(new_n485), .ZN(G160));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n461), .C2(G112), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n466), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n472), .A2(new_n474), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT72), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G124), .ZN(new_n495));
  OR3_X1    g070(.A1(new_n494), .A2(KEYINPUT73), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT73), .B1(new_n494), .B2(new_n495), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(G162));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT74), .B(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n481), .B2(new_n482), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT74), .A2(G114), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT74), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2105), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n500), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n503), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n469), .B2(new_n470), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(new_n512), .A3(KEYINPUT75), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n472), .A2(new_n474), .A3(G138), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT4), .B1(new_n471), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n472), .A2(new_n474), .A3(G138), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(new_n462), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n505), .A2(new_n513), .B1(new_n515), .B2(new_n518), .ZN(G164));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(G62), .ZN(new_n523));
  AND2_X1   g098(.A1(G75), .A2(G543), .ZN(new_n524));
  OAI21_X1  g099(.A(G651), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT76), .B1(new_n526), .B2(KEYINPUT6), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n529), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n531), .A2(G50), .A3(G543), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n531), .A2(G88), .A3(new_n532), .A4(new_n522), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n525), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G166));
  XNOR2_X1  g111(.A(new_n522), .B(KEYINPUT77), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n531), .A2(new_n532), .A3(new_n522), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n531), .A2(G543), .A3(new_n532), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n541), .A2(new_n542), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n538), .A2(new_n544), .A3(new_n546), .A4(new_n540), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT78), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(G168));
  AOI22_X1  g125(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n526), .ZN(new_n552));
  AOI22_X1  g127(.A1(G52), .A2(new_n545), .B1(new_n543), .B2(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(new_n537), .A2(G56), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n526), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n545), .A2(G43), .ZN(new_n559));
  INV_X1    g134(.A(new_n543), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n545), .A2(G53), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n545), .A2(new_n571), .A3(G53), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  XOR2_X1   g149(.A(KEYINPUT5), .B(G543), .Z(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n543), .A2(G91), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND2_X1  g155(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n525), .A2(new_n582), .A3(new_n533), .A4(new_n534), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(G303));
  NAND2_X1  g159(.A1(new_n543), .A2(G87), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n545), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n575), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n522), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(G74), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n585), .B(new_n586), .C1(new_n526), .C2(new_n590), .ZN(G288));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n520), .B2(new_n521), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n531), .A2(G48), .A3(G543), .A4(new_n532), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n531), .A2(G86), .A3(new_n532), .A4(new_n522), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n537), .A2(G60), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n526), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n545), .A2(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n560), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G171), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n543), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n575), .ZN(new_n614));
  AOI22_X1  g189(.A1(G54), .A2(new_n545), .B1(new_n614), .B2(G651), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT81), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n607), .B1(new_n618), .B2(G868), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT82), .ZN(G284));
  XNOR2_X1  g195(.A(new_n619), .B(KEYINPUT83), .ZN(G321));
  NOR2_X1   g196(.A1(G299), .A2(G868), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g198(.A(new_n622), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n617), .B1(new_n625), .B2(G860), .ZN(G148));
  OAI21_X1  g201(.A(G868), .B1(new_n618), .B2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI221_X1 g204(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n461), .C2(G111), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n489), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n493), .B2(G123), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n480), .A2(KEYINPUT3), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n479), .A2(G2104), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n466), .A2(G2104), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n641), .B(new_n642), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT13), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n636), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT87), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT86), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT14), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n659), .B2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT91), .B(KEYINPUT17), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT89), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT92), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n665), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(new_n672), .C1(new_n667), .C2(new_n670), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n665), .A3(new_n672), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n674), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n683), .A3(new_n684), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n683), .A2(new_n684), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n694), .C1(new_n690), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G24), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT96), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n605), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1986), .ZN(new_n708));
  NOR2_X1   g283(.A1(G25), .A2(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n493), .A2(G119), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n489), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n461), .A2(G107), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n713), .A2(G131), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n709), .B1(new_n718), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n708), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n704), .A2(G23), .ZN(new_n723));
  INV_X1    g298(.A(G288), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n704), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT33), .B(G1976), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n725), .B(new_n726), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n704), .A2(G22), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G166), .B2(new_n704), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1971), .ZN(new_n730));
  MUX2_X1   g305(.A(G6), .B(G305), .S(G16), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XOR2_X1   g307(.A(new_n731), .B(new_n732), .Z(new_n733));
  NOR3_X1   g308(.A1(new_n727), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n722), .B1(new_n719), .B2(new_n721), .C1(new_n735), .C2(KEYINPUT34), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(KEYINPUT34), .B2(new_n735), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT36), .Z(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT104), .B(KEYINPUT29), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2090), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n635), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT102), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n704), .A2(G20), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT23), .Z(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G299), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1956), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n704), .A2(G4), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n617), .B2(new_n704), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1348), .ZN(new_n755));
  NAND2_X1  g330(.A1(G160), .A2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT24), .B(G34), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(new_n745), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT99), .ZN(new_n759));
  AOI21_X1  g334(.A(G2084), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n756), .A2(G2084), .A3(new_n759), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n745), .B1(new_n763), .B2(G28), .ZN(new_n764));
  AOI21_X1  g339(.A(KEYINPUT103), .B1(new_n763), .B2(G28), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n763), .A2(KEYINPUT103), .A3(G28), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  NOR2_X1   g345(.A1(G164), .A2(new_n745), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G27), .B2(new_n745), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n760), .B(new_n769), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n563), .B2(G16), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G1341), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(G1341), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n772), .A2(new_n770), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n773), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n744), .A2(new_n752), .A3(new_n755), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G16), .A2(G21), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G168), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT101), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1966), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n745), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  INV_X1    g362(.A(G139), .ZN(new_n788));
  OAI21_X1  g363(.A(KEYINPUT97), .B1(new_n489), .B2(new_n788), .ZN(new_n789));
  OR3_X1    g364(.A1(new_n489), .A2(KEYINPUT97), .A3(new_n788), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT98), .Z(new_n792));
  AOI22_X1  g367(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n461), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n785), .B1(new_n795), .B2(new_n745), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(G2072), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n745), .A2(G32), .ZN(new_n798));
  INV_X1    g373(.A(G141), .ZN(new_n799));
  INV_X1    g374(.A(G105), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n489), .A2(new_n799), .B1(new_n800), .B2(new_n640), .ZN(new_n801));
  AND3_X1   g376(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT100), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT26), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n801), .B(new_n804), .C1(G129), .C2(new_n493), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n798), .B1(new_n805), .B2(new_n745), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n806), .B(new_n807), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n745), .A2(G26), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT28), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n493), .A2(G128), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n461), .A2(G116), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n713), .A2(G140), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(G29), .ZN(new_n817));
  INV_X1    g392(.A(G2067), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n808), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n796), .A2(G2072), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n704), .A2(G5), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G171), .B2(new_n704), .ZN(new_n823));
  INV_X1    g398(.A(G1961), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  AND4_X1   g400(.A1(new_n797), .A2(new_n820), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  AND4_X1   g401(.A1(new_n738), .A2(new_n780), .A3(new_n784), .A4(new_n826), .ZN(G311));
  NAND4_X1  g402(.A1(new_n738), .A2(new_n780), .A3(new_n784), .A4(new_n826), .ZN(G150));
  XOR2_X1   g403(.A(KEYINPUT106), .B(G55), .Z(new_n829));
  AOI22_X1  g404(.A1(G93), .A2(new_n543), .B1(new_n545), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n537), .A2(G67), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n526), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI211_X1 g410(.A(KEYINPUT105), .B(new_n526), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G860), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n617), .A2(G559), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT107), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n837), .A2(new_n563), .ZN(new_n844));
  INV_X1    g419(.A(new_n563), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n835), .B2(new_n836), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n838), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n840), .B1(new_n850), .B2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n635), .B(KEYINPUT108), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G160), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n713), .A2(G142), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT109), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n493), .A2(G130), .ZN(new_n858));
  OAI221_X1 g433(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n461), .C2(G118), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n718), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n805), .B(new_n816), .ZN(new_n862));
  INV_X1    g437(.A(new_n643), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n816), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n805), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n643), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n795), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n712), .A2(new_n717), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n860), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n864), .A3(new_n867), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n870), .B1(new_n869), .B2(new_n873), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n483), .A2(new_n511), .B1(new_n508), .B2(new_n509), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n517), .B1(new_n516), .B2(new_n483), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n514), .A2(new_n639), .A3(KEYINPUT4), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n875), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n510), .A2(new_n512), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n515), .B2(new_n518), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n869), .A2(new_n873), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n795), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n883), .B1(new_n885), .B2(new_n874), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n855), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n880), .B1(new_n875), .B2(new_n876), .ZN(new_n889));
  INV_X1    g464(.A(new_n855), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n883), .A3(new_n874), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g469(.A(new_n847), .B(KEYINPUT110), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n618), .A2(G559), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n616), .A2(G299), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n616), .A2(G299), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(KEYINPUT41), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n899), .B2(new_n900), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n898), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n901), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT111), .B1(new_n906), .B2(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n897), .A2(new_n901), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n605), .B(G305), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G288), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(KEYINPUT42), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n915), .B(new_n916), .Z(new_n917));
  AND3_X1   g492(.A1(new_n909), .A2(new_n910), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n909), .B2(new_n910), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g496(.A(new_n920), .B1(G868), .B2(new_n837), .ZN(G331));
  AOI21_X1  g497(.A(G301), .B1(G168), .B2(KEYINPUT113), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(G168), .A2(KEYINPUT113), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n847), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n847), .A2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(G168), .A2(KEYINPUT113), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n848), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n847), .A2(new_n925), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n923), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n908), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n928), .A2(new_n932), .A3(new_n906), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n913), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(new_n888), .ZN(new_n937));
  INV_X1    g512(.A(new_n935), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n928), .A2(new_n932), .B1(new_n905), .B2(new_n907), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT114), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT114), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n934), .A2(new_n941), .A3(new_n935), .ZN(new_n942));
  INV_X1    g517(.A(new_n913), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT43), .B1(new_n937), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n902), .A2(new_n904), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n928), .B2(new_n932), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n943), .B1(new_n938), .B2(new_n947), .ZN(new_n948));
  AND4_X1   g523(.A1(KEYINPUT43), .A2(new_n948), .A3(new_n936), .A4(new_n888), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT44), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n937), .B2(new_n944), .ZN(new_n953));
  AND4_X1   g528(.A1(new_n952), .A2(new_n948), .A3(new_n936), .A4(new_n888), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n955), .ZN(G397));
  INV_X1    g531(.A(KEYINPUT127), .ZN(new_n957));
  INV_X1    g532(.A(G40), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n958), .B(new_n465), .C1(new_n478), .C2(new_n485), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT116), .B1(new_n883), .B2(G1384), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n880), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1981), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g542(.A1(G305), .A2(G1981), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(KEYINPUT49), .A3(new_n966), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT49), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n964), .A2(G8), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(G288), .A2(G1976), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(G8), .B(new_n964), .C1(new_n975), .C2(KEYINPUT121), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(KEYINPUT121), .B2(new_n975), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n724), .A2(G1976), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n964), .A2(G8), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT52), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT118), .ZN(new_n981));
  INV_X1    g556(.A(G1976), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(G288), .B2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n964), .A2(G8), .A3(new_n978), .A4(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n979), .A2(new_n986), .A3(KEYINPUT52), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n981), .A2(new_n985), .A3(KEYINPUT119), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n465), .ZN(new_n993));
  INV_X1    g568(.A(new_n485), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT71), .B1(new_n484), .B2(new_n467), .ZN(new_n995));
  OAI211_X1 g570(.A(G40), .B(new_n993), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n515), .A2(new_n518), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n502), .A2(new_n499), .A3(new_n504), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT75), .B1(new_n510), .B2(new_n512), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n962), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n960), .A2(new_n1003), .A3(new_n963), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n743), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(G164), .B2(G1384), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n880), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n959), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1971), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n581), .A2(G8), .A3(new_n583), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n977), .B1(new_n992), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n505), .A2(new_n513), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n1019), .B2(new_n997), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n996), .B1(new_n1003), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n880), .A2(new_n961), .A3(new_n962), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n961), .B1(new_n880), .B2(new_n962), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT50), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1956), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n573), .B2(new_n578), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n573), .A2(new_n1026), .A3(new_n578), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT56), .B(G2072), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1007), .A2(new_n959), .A3(new_n1008), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1025), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT123), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1348), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n964), .A2(G2067), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1348), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1022), .A2(new_n1023), .A3(KEYINPUT50), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n959), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1022), .A2(new_n996), .A3(new_n1023), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n818), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(KEYINPUT123), .A3(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1038), .A2(new_n1046), .A3(new_n610), .A4(new_n615), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1030), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1034), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1036), .A2(new_n1037), .A3(new_n1035), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT123), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT60), .B(new_n616), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1956), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1003), .B1(new_n960), .B2(new_n963), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1000), .A2(new_n1003), .A3(new_n962), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n959), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1029), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n1027), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1059), .A3(new_n1032), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1048), .A2(KEYINPUT61), .A3(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1007), .A2(new_n959), .A3(new_n1008), .ZN(new_n1062));
  INV_X1    g637(.A(G1996), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT58), .B(G1341), .Z(new_n1064));
  AOI22_X1  g639(.A1(new_n1062), .A2(new_n1063), .B1(new_n964), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT59), .B1(new_n1065), .B2(new_n845), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1064), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n1044), .A2(new_n1067), .B1(new_n1009), .B2(G1996), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n563), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1059), .B1(new_n1057), .B2(new_n1032), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1034), .B2(new_n1073), .ZN(new_n1074));
  AND4_X1   g649(.A1(new_n1052), .A2(new_n1061), .A3(new_n1071), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n616), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1038), .A2(new_n1046), .A3(new_n1076), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1049), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G8), .ZN(new_n1082));
  INV_X1    g657(.A(G1966), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n959), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT45), .B1(new_n960), .B2(new_n963), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1002), .A2(new_n1087), .A3(new_n1004), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1082), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n547), .A2(G8), .A3(new_n549), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT124), .A4(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1089), .A2(new_n1094), .A3(KEYINPUT51), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n824), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1009), .B2(G2078), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n996), .B1(KEYINPUT45), .B2(new_n1020), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1006), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1102), .A2(G2078), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G171), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT45), .B1(new_n880), .B2(new_n962), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n996), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(KEYINPUT125), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n996), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1008), .B(new_n1106), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(G301), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1109), .A2(new_n1116), .A3(KEYINPUT126), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(G301), .A4(new_n1115), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(G301), .A3(new_n1107), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1119), .A2(new_n1115), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT54), .B(new_n1123), .C1(new_n1124), .C2(G301), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1021), .A2(new_n1024), .A3(new_n743), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1082), .B1(new_n1126), .B2(new_n1011), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1016), .B1(new_n1015), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(new_n988), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1100), .A2(new_n1122), .A3(new_n1125), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1018), .B1(new_n1081), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1082), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1089), .B(G168), .C1(new_n1133), .C2(new_n1015), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1016), .A2(KEYINPUT63), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n992), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n992), .B2(new_n1136), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1089), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(G286), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT63), .B1(new_n1129), .B2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n957), .B1(new_n1131), .B2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1100), .A2(new_n1129), .A3(new_n1125), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1079), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1145), .A2(new_n1077), .A3(new_n616), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1052), .A2(new_n1071), .A3(new_n1074), .A4(new_n1061), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1146), .A2(new_n1147), .B1(new_n1148), .B2(new_n1034), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1144), .A2(new_n1149), .A3(new_n1122), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1141), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n992), .A2(new_n1136), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT122), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n992), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1150), .A2(new_n1155), .A3(KEYINPUT127), .A4(new_n1018), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1109), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1157), .A2(new_n1129), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1143), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n959), .A2(new_n1110), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT115), .Z(new_n1163));
  NOR2_X1   g738(.A1(new_n718), .A2(new_n720), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n871), .A2(new_n721), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n816), .B(new_n818), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1063), .B2(new_n805), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1162), .A2(G1996), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1163), .A2(new_n1168), .B1(new_n805), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1162), .ZN(new_n1172));
  INV_X1    g747(.A(G1986), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n605), .B(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1161), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1163), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1170), .A2(new_n1165), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n865), .A2(new_n818), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1169), .B(KEYINPUT46), .Z(new_n1181));
  AND2_X1   g756(.A1(new_n1167), .A2(new_n805), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT47), .Z(new_n1184));
  INV_X1    g759(.A(new_n1171), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1172), .A2(new_n1173), .A3(new_n605), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT48), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1180), .B(new_n1184), .C1(new_n1185), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1176), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(G319), .ZN(new_n1191));
  OR2_X1    g765(.A1(G227), .A2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g766(.A1(G401), .A2(G229), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1193), .A2(new_n893), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1195), .ZN(G308));
  OAI211_X1 g770(.A(new_n1193), .B(new_n893), .C1(new_n953), .C2(new_n954), .ZN(G225));
endmodule


