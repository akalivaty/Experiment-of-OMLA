//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT0), .B(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G101), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n210), .A2(G101), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n205), .A2(new_n208), .A3(new_n214), .A4(new_n209), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n203), .B(new_n212), .C1(new_n213), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n196), .A2(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n194), .A2(G143), .ZN(new_n220));
  OAI211_X1 g034(.A(G128), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n195), .B(new_n197), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n204), .A2(G107), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n207), .A2(G104), .ZN(new_n226));
  OAI21_X1  g040(.A(G101), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n215), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n228), .A3(KEYINPUT10), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n221), .A2(new_n215), .A3(new_n227), .A4(new_n223), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n234), .A2(new_n235), .A3(G137), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT65), .A2(G134), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT65), .A2(G134), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n237), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n235), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT65), .A2(G134), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n242), .A3(G137), .A4(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(G137), .B1(new_n245), .B2(new_n246), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(KEYINPUT11), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n243), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n245), .A2(G137), .A3(new_n246), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n236), .B1(new_n251), .B2(KEYINPUT66), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n240), .B1(new_n238), .B2(new_n239), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n234), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n252), .A2(new_n253), .A3(new_n247), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n193), .B1(new_n233), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n221), .A2(new_n223), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n215), .A2(new_n227), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n230), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT12), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n257), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n256), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n241), .A2(new_n242), .B1(new_n254), .B2(new_n234), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n253), .B1(new_n268), .B2(new_n252), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n230), .B(KEYINPUT10), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n217), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n233), .A2(new_n257), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n193), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n187), .B(new_n188), .C1(new_n266), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n233), .A2(new_n257), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n233), .A2(new_n257), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n192), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n257), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n272), .B(new_n193), .C1(new_n281), .C2(new_n263), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT81), .A3(new_n187), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n272), .B1(new_n281), .B2(new_n263), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n192), .ZN(new_n287));
  INV_X1    g101(.A(new_n258), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n273), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n286), .A2(new_n192), .B1(new_n288), .B2(new_n273), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT80), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n285), .B1(new_n295), .B2(new_n187), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT90), .ZN(new_n297));
  INV_X1    g111(.A(G237), .ZN(new_n298));
  INV_X1    g112(.A(G953), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(G214), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n196), .ZN(new_n301));
  NOR2_X1   g115(.A1(G237), .A2(G953), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G131), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT17), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n253), .A3(new_n303), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(KEYINPUT75), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(G125), .A3(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(KEYINPUT16), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n310), .B2(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n194), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n316), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n304), .A2(KEYINPUT17), .A3(G131), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n308), .A2(new_n317), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G113), .B(G122), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(new_n204), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT89), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n301), .A2(new_n303), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT18), .A2(G131), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n194), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n311), .A2(G146), .A3(new_n313), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n327), .A2(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n328), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n304), .A2(KEYINPUT88), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT88), .B1(new_n304), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n321), .A2(new_n326), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n188), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n326), .B1(new_n321), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n297), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n321), .A2(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n325), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n343), .A2(KEYINPUT90), .A3(new_n188), .A4(new_n338), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(G475), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n305), .A2(new_n307), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n311), .A2(new_n313), .ZN(new_n347));
  MUX2_X1   g161(.A(new_n329), .B(new_n347), .S(KEYINPUT19), .Z(new_n348));
  OAI211_X1 g162(.A(new_n346), .B(new_n319), .C1(new_n348), .C2(G146), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n337), .A3(new_n324), .ZN(new_n350));
  NOR2_X1   g164(.A1(G475), .A2(G902), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n319), .A2(new_n320), .A3(new_n317), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n327), .B2(new_n328), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n334), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n308), .A2(new_n352), .B1(new_n355), .B2(new_n332), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n350), .B(new_n351), .C1(new_n356), .C2(new_n324), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT20), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n342), .A2(new_n323), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n350), .A4(new_n351), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n345), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G478), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT15), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT13), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT91), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT13), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n367), .A2(new_n369), .A3(G128), .A4(new_n196), .ZN(new_n370));
  XNOR2_X1  g184(.A(G128), .B(G143), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n370), .B(G134), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G122), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G116), .ZN(new_n376));
  INV_X1    g190(.A(G116), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G122), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n378), .A3(new_n207), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(new_n245), .A3(new_n246), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n385));
  INV_X1    g199(.A(new_n381), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n245), .A2(new_n246), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n372), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n383), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n377), .A2(KEYINPUT14), .A3(G122), .ZN(new_n390));
  OAI211_X1 g204(.A(G107), .B(new_n390), .C1(new_n379), .C2(KEYINPUT14), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n384), .A2(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n374), .A2(new_n382), .A3(KEYINPUT92), .A4(new_n383), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT9), .B(G234), .ZN(new_n394));
  INV_X1    g208(.A(G217), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n394), .A2(new_n395), .A3(G953), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n365), .B1(new_n399), .B2(G902), .ZN(new_n400));
  OAI221_X1 g214(.A(new_n188), .B1(KEYINPUT15), .B2(new_n364), .C1(new_n397), .C2(new_n398), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(G234), .A2(G237), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n403), .A2(G952), .A3(new_n299), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(G902), .A3(G953), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n405), .B(KEYINPUT93), .Z(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT21), .B(G898), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n363), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G221), .B1(new_n394), .B2(G902), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n410), .B(KEYINPUT78), .Z(new_n411));
  XOR2_X1   g225(.A(new_n411), .B(KEYINPUT79), .Z(new_n412));
  OAI21_X1  g226(.A(G214), .B1(G237), .B2(G902), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT82), .Z(new_n414));
  OAI21_X1  g228(.A(G210), .B1(G237), .B2(G902), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT2), .B(G113), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OR2_X1    g231(.A1(KEYINPUT68), .A2(G119), .ZN(new_n418));
  NAND2_X1  g232(.A1(KEYINPUT68), .A2(G119), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n377), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(G116), .A2(G119), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n417), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n421), .ZN(new_n423));
  INV_X1    g237(.A(new_n419), .ZN(new_n424));
  NOR2_X1   g238(.A1(KEYINPUT68), .A2(G119), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n416), .B(new_n423), .C1(new_n426), .C2(new_n377), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n210), .A2(G101), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n430), .A3(new_n212), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT5), .B1(new_n420), .B2(new_n421), .ZN(new_n432));
  INV_X1    g246(.A(G113), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n426), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n422), .A3(new_n228), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n431), .A2(new_n437), .A3(KEYINPUT83), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G122), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n299), .A2(G224), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(KEYINPUT85), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n449));
  AOI21_X1  g263(.A(G125), .B1(new_n221), .B2(new_n223), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n202), .A2(G125), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n449), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n448), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(KEYINPUT0), .A2(G128), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n198), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n219), .B2(new_n220), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n310), .B1(new_n459), .B2(new_n199), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT84), .B1(new_n460), .B2(new_n450), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n447), .A3(new_n454), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n431), .A2(new_n437), .A3(KEYINPUT83), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT83), .B1(new_n431), .B2(new_n437), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n464), .A2(new_n465), .A3(new_n443), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n431), .A2(new_n437), .A3(new_n443), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n445), .B(new_n463), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT68), .B(G119), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n471));
  OAI21_X1  g285(.A(G113), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(KEYINPUT86), .B(G113), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n432), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n476), .A2(new_n477), .A3(new_n422), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n476), .B2(new_n422), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n228), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n443), .B(KEYINPUT8), .Z(new_n481));
  AND2_X1   g295(.A1(new_n436), .A2(new_n422), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n260), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n461), .A2(KEYINPUT7), .A3(new_n447), .A4(new_n454), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n447), .A2(KEYINPUT7), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n460), .B2(new_n450), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n485), .A2(new_n467), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n415), .B1(new_n469), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n469), .A2(new_n489), .A3(new_n415), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n414), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND4_X1   g307(.A1(new_n296), .A2(new_n409), .A3(new_n412), .A4(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n203), .B1(new_n267), .B2(new_n269), .ZN(new_n495));
  INV_X1    g309(.A(new_n428), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n240), .A2(G134), .ZN(new_n497));
  OAI21_X1  g311(.A(G131), .B1(new_n248), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n256), .A2(new_n498), .A3(new_n224), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT26), .B(G101), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n302), .A2(G210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n502), .A2(KEYINPUT29), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n202), .B1(new_n250), .B2(new_n256), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n256), .A2(new_n498), .A3(new_n224), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n428), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n495), .A2(KEYINPUT72), .A3(new_n496), .A4(new_n499), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n509), .B1(KEYINPUT28), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT73), .B1(new_n517), .B2(G902), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n512), .A2(new_n513), .A3(new_n428), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT28), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n507), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n256), .A2(new_n523), .A3(new_n498), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n256), .B2(new_n498), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n524), .A2(new_n525), .A3(new_n259), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n202), .B(KEYINPUT64), .Z(new_n527));
  AND2_X1   g341(.A1(new_n527), .A2(new_n257), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n522), .B(new_n428), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n256), .A2(new_n498), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT67), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n256), .A2(new_n523), .A3(new_n498), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n224), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n257), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n496), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n521), .B1(new_n530), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n541), .A3(new_n535), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT30), .B1(new_n512), .B2(new_n513), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n496), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n507), .B1(new_n544), .B2(new_n519), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n539), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n515), .A2(new_n514), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n501), .B1(new_n548), .B2(new_n511), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n547), .B(new_n188), .C1(new_n549), .C2(new_n509), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n518), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G472), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT31), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n500), .A2(new_n555), .A3(new_n508), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n500), .B2(new_n508), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n554), .B1(new_n558), .B2(new_n544), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n542), .A2(new_n543), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n428), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT70), .B1(new_n519), .B2(new_n507), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n500), .A2(new_n555), .A3(new_n508), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n564), .A3(KEYINPUT31), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n502), .B1(new_n530), .B2(new_n538), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n559), .A2(new_n565), .B1(new_n566), .B2(new_n507), .ZN(new_n567));
  NOR2_X1   g381(.A1(G472), .A2(G902), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n553), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n558), .A2(new_n554), .A3(new_n544), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT31), .B1(new_n561), .B2(new_n564), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n428), .B1(new_n526), .B2(new_n528), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT71), .A3(new_n500), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n501), .B1(new_n536), .B2(new_n522), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n520), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n571), .A2(new_n572), .B1(new_n576), .B2(new_n508), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n568), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n552), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n418), .A2(G128), .A3(new_n419), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n222), .A2(G119), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT23), .B1(new_n470), .B2(new_n222), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT76), .B(G110), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n581), .A2(new_n582), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT24), .B(G110), .Z(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n319), .B(new_n330), .C1(new_n586), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n319), .A2(new_n317), .ZN(new_n591));
  OAI21_X1  g405(.A(G110), .B1(new_n583), .B2(new_n584), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(new_n588), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT22), .B(G137), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n299), .A2(G221), .A3(G234), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n590), .A2(new_n594), .A3(new_n598), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT77), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT25), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n600), .A2(new_n608), .A3(new_n601), .A4(new_n604), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n395), .B1(G234), .B2(new_n188), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT74), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n600), .A2(new_n601), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n494), .A2(new_n579), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  OAI21_X1  g432(.A(G472), .B1(new_n567), .B2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n577), .A2(new_n568), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n296), .A2(new_n616), .A3(new_n412), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n492), .B1(new_n490), .B2(KEYINPUT94), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n469), .A2(new_n489), .A3(new_n627), .A4(new_n415), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n414), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n408), .ZN(new_n630));
  INV_X1    g444(.A(new_n363), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n399), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT33), .B1(new_n397), .B2(new_n398), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(G478), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n364), .A2(new_n188), .ZN(new_n636));
  INV_X1    g450(.A(new_n398), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(new_n639), .B2(new_n364), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n629), .A2(new_n630), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n358), .A2(new_n647), .A3(new_n361), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n357), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n402), .A2(new_n648), .A3(new_n345), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n408), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n629), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n625), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n599), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n595), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n614), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n612), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n622), .A2(new_n494), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  AND3_X1   g476(.A1(new_n296), .A2(new_n412), .A3(new_n659), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT96), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n406), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n404), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n664), .B1(new_n650), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n648), .A2(new_n649), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n344), .A2(G475), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n670), .A2(new_n341), .B1(new_n400), .B2(new_n401), .ZN(new_n671));
  INV_X1    g485(.A(new_n667), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n669), .A2(new_n671), .A3(KEYINPUT96), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n579), .A2(new_n663), .A3(new_n629), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  NAND2_X1  g491(.A1(new_n491), .A2(new_n492), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n363), .A2(new_n402), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n659), .A3(new_n414), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n667), .B(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n296), .A2(new_n412), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n683), .B1(new_n686), .B2(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n561), .A2(new_n564), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n516), .A2(new_n507), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n690), .B2(G902), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n570), .A2(new_n578), .A3(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n687), .B(new_n692), .C1(KEYINPUT40), .C2(new_n686), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  NOR3_X1   g508(.A1(new_n631), .A2(new_n641), .A3(new_n667), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n629), .A2(KEYINPUT99), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT99), .B1(new_n629), .B2(new_n695), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n579), .B(new_n663), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NAND2_X1  g513(.A1(new_n280), .A2(new_n282), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n187), .B1(new_n700), .B2(new_n188), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n411), .B(new_n701), .C1(new_n277), .C2(new_n284), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(new_n616), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n643), .A2(new_n579), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND3_X1  g520(.A1(new_n579), .A2(new_n652), .A3(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  AND2_X1   g522(.A1(new_n409), .A2(new_n659), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n629), .A2(new_n710), .A3(new_n702), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n710), .B1(new_n629), .B2(new_n702), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n579), .B(new_n709), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NAND2_X1  g528(.A1(new_n577), .A2(new_n188), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n507), .B1(new_n549), .B2(new_n520), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n571), .B2(new_n572), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n715), .A2(G472), .B1(new_n568), .B2(new_n717), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n414), .B(new_n681), .C1(new_n626), .C2(new_n628), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n285), .B1(new_n187), .B2(new_n283), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n411), .A3(new_n408), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n616), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n568), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n619), .A2(new_n724), .A3(new_n659), .A4(new_n695), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n711), .B2(new_n712), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  INV_X1    g541(.A(new_n492), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n728), .A2(new_n490), .A3(new_n414), .ZN(new_n729));
  OAI21_X1  g543(.A(G469), .B1(new_n293), .B2(G902), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n275), .A2(new_n276), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT81), .B1(new_n283), .B2(new_n187), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n411), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n695), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n579), .A2(new_n737), .A3(new_n616), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n577), .A2(KEYINPUT101), .A3(KEYINPUT32), .A4(new_n568), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT101), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n742), .B1(new_n567), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n552), .A3(new_n570), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(KEYINPUT42), .A3(new_n616), .A4(new_n737), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n740), .A2(KEYINPUT102), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n253), .ZN(G33));
  NOR2_X1   g566(.A1(new_n674), .A2(new_n735), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n579), .A3(new_n616), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  OAI21_X1  g570(.A(G469), .B1(new_n290), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n292), .A2(new_n294), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(new_n756), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n187), .A2(new_n188), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT103), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n761), .A2(new_n762), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n285), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n734), .A3(new_n685), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT104), .ZN(new_n770));
  INV_X1    g584(.A(new_n641), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n631), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(KEYINPUT106), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(new_n772), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT106), .B1(new_n772), .B2(new_n773), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n621), .A3(new_n659), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  INV_X1    g597(.A(new_n414), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n491), .A2(new_n784), .A3(new_n492), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n779), .A2(new_n781), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT107), .Z(new_n788));
  NAND4_X1  g602(.A1(new_n770), .A2(new_n782), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NOR4_X1   g604(.A1(new_n579), .A2(new_n616), .A3(new_n736), .A4(new_n785), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n768), .A2(new_n734), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n768), .A2(KEYINPUT47), .A3(new_n734), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n309), .ZN(G42));
  XNOR2_X1  g612(.A(new_n720), .B(KEYINPUT49), .ZN(new_n799));
  INV_X1    g613(.A(new_n772), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n616), .A3(new_n412), .A4(new_n784), .ZN(new_n801));
  OR4_X1    g615(.A1(new_n692), .A2(new_n799), .A3(new_n680), .A4(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n803));
  OAI211_X1 g617(.A(new_n795), .B(new_n796), .C1(new_n412), .C2(new_n720), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n616), .A2(new_n778), .A3(new_n404), .A4(new_n718), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n729), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n404), .A2(new_n778), .A3(new_n702), .A4(new_n729), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n718), .A2(new_n659), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n702), .A2(new_n616), .A3(new_n404), .A4(new_n729), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n692), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n771), .A2(new_n363), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n809), .A2(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n680), .A2(new_n784), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n805), .A2(new_n702), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT50), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT118), .Z(new_n821));
  OAI21_X1  g635(.A(new_n803), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n809), .A2(new_n616), .A3(new_n745), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT48), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n805), .B1(new_n711), .B2(new_n712), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n299), .A2(G952), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n813), .B2(new_n642), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n816), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n822), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n659), .A2(new_n667), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n733), .A2(new_n734), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n733), .A2(new_n834), .A3(new_n837), .A4(new_n734), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n719), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n570), .A2(new_n578), .A3(new_n691), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT113), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n681), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n838), .A2(new_n629), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n692), .A4(new_n836), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n726), .A2(new_n698), .A3(new_n676), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT52), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n726), .A2(new_n698), .A3(new_n676), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n841), .A2(new_n845), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n713), .A2(new_n617), .A3(new_n704), .A4(new_n707), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT109), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n631), .A2(new_n630), .A3(new_n402), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n784), .B1(new_n728), .B2(new_n490), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n402), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n363), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n493), .A2(KEYINPUT109), .A3(new_n630), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n493), .A2(new_n642), .A3(new_n630), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n622), .A3(new_n623), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n660), .A3(new_n722), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n737), .A2(new_n718), .A3(new_n659), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n754), .A2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n859), .A2(new_n345), .A3(new_n672), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n729), .A3(new_n870), .A4(new_n669), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n669), .A2(new_n345), .A3(new_n859), .A4(new_n672), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT110), .B1(new_n872), .B2(new_n785), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n579), .A3(new_n663), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT111), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n874), .A2(new_n579), .A3(new_n663), .A4(KEYINPUT111), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n868), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n866), .A2(new_n749), .A3(new_n750), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n853), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n853), .B2(new_n880), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n833), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n890), .B(new_n881), .C1(new_n853), .C2(new_n880), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n747), .A4(new_n879), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n853), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n833), .A2(new_n889), .A3(new_n891), .A4(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n832), .A2(new_n888), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n802), .B1(new_n896), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n299), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n893), .B1(new_n885), .B2(KEYINPUT116), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n188), .B1(new_n901), .B2(new_n891), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n902), .B2(G210), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n445), .B1(new_n466), .B2(new_n468), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n463), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n903), .B2(new_n906), .ZN(G51));
  NAND3_X1  g722(.A1(new_n889), .A2(new_n891), .A3(new_n894), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n901), .A2(new_n833), .A3(new_n891), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n760), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n700), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n902), .A2(new_n759), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n899), .B1(new_n916), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n359), .A2(new_n350), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n899), .ZN(G60));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n633), .A2(new_n634), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT120), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n636), .B(KEYINPUT59), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n833), .B1(new_n901), .B2(new_n891), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n924), .B(new_n928), .C1(new_n895), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n900), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n924), .B1(new_n912), .B2(new_n928), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT122), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n928), .B1(new_n895), .B2(new_n929), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n936), .A3(new_n900), .A4(new_n930), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n888), .A2(new_n895), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n926), .B1(new_n938), .B2(new_n927), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n933), .A2(new_n937), .A3(new_n939), .ZN(G63));
  XNOR2_X1  g754(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT60), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n909), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n613), .B(KEYINPUT124), .Z(new_n945));
  AOI21_X1  g759(.A(new_n899), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n909), .A2(new_n657), .A3(new_n943), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n941), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  XNOR2_X1  g767(.A(new_n866), .B(KEYINPUT126), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n299), .ZN(new_n955));
  INV_X1    g769(.A(G224), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n407), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n904), .B1(G898), .B2(new_n299), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  NAND2_X1  g774(.A1(new_n579), .A2(new_n616), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n729), .B1(new_n642), .B2(new_n860), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n686), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n797), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n693), .A2(new_n849), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n789), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n299), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n560), .B(new_n348), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(G900), .B2(G953), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n770), .A2(new_n616), .A3(new_n719), .A4(new_n745), .ZN(new_n972));
  INV_X1    g786(.A(new_n754), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n797), .A2(new_n973), .A3(new_n847), .ZN(new_n974));
  INV_X1    g788(.A(new_n751), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n789), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n971), .B1(new_n976), .B2(G953), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n190), .B2(new_n665), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n970), .B(new_n977), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n978), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n976), .B2(new_n954), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n544), .A2(new_n519), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n507), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n984), .B1(new_n967), .B2(new_n954), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n986), .A2(new_n507), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n899), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n884), .A2(new_n887), .ZN(new_n992));
  INV_X1    g806(.A(new_n984), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n688), .B2(new_n545), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n992), .B2(new_n994), .ZN(G57));
endmodule


