//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n651, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G210), .B1(G237), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G122), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT73), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(new_n194), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n195), .A2(new_n198), .A3(new_n202), .A4(new_n199), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G116), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n214), .A3(G101), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n194), .A2(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n197), .A2(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n203), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT5), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(G113), .C1(KEYINPUT5), .C2(new_n206), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n211), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n193), .B1(new_n216), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n224), .A2(KEYINPUT6), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(new_n223), .A3(new_n192), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT74), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT74), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n216), .A2(new_n228), .A3(new_n223), .A4(new_n192), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT6), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n225), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G146), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n233), .A2(KEYINPUT64), .A3(G143), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n244));
  INV_X1    g058(.A(G125), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n236), .A2(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n234), .A2(new_n246), .A3(new_n247), .A4(G128), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n236), .A2(G146), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT64), .B1(new_n233), .B2(G143), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n235), .A2(new_n236), .A3(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n245), .B(new_n248), .C1(new_n253), .C2(new_n241), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT75), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n234), .A2(new_n246), .A3(new_n256), .ZN(new_n261));
  OAI21_X1  g075(.A(G125), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n249), .A2(new_n255), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G224), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n263), .B(new_n265), .Z(new_n266));
  AND2_X1   g080(.A1(new_n232), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(KEYINPUT7), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n222), .A2(new_n211), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n203), .A2(new_n219), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n223), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n192), .B(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n249), .A2(new_n255), .A3(new_n262), .A4(new_n265), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT76), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n277), .A2(new_n278), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n263), .A2(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n227), .A2(new_n229), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n191), .B1(new_n267), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n232), .A2(new_n266), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(new_n287), .A3(new_n190), .A4(new_n286), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n189), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G128), .B(G143), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n236), .A2(G128), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n295), .A2(KEYINPUT13), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n294), .A2(G134), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G134), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G122), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n207), .A2(G122), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n197), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n197), .B1(new_n301), .B2(new_n302), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT14), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n301), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G107), .B1(new_n302), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n240), .A2(G143), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n295), .A2(new_n311), .A3(new_n298), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n298), .B1(new_n295), .B2(new_n311), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI22_X1  g128(.A1(new_n297), .A2(new_n306), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  OAI221_X1 g134(.A(new_n318), .B1(new_n310), .B2(new_n314), .C1(new_n297), .C2(new_n306), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT80), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n323), .A3(new_n319), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n287), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G478), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT15), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n327), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n322), .A2(new_n287), .A3(new_n324), .A4(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G475), .ZN(new_n332));
  INV_X1    g146(.A(G131), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT65), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G131), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G237), .A2(G953), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n338), .A2(G143), .A3(G214), .ZN(new_n339));
  AOI21_X1  g153(.A(G143), .B1(new_n338), .B2(G214), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n342));
  INV_X1    g156(.A(G237), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n264), .A3(G214), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n236), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n334), .A2(new_n336), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n338), .A2(G143), .A3(G214), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n341), .A2(new_n342), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n345), .B2(new_n347), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT17), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT16), .ZN(new_n352));
  INV_X1    g166(.A(G140), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G125), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n245), .A2(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(G146), .B(new_n354), .C1(new_n357), .C2(new_n352), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n354), .B1(new_n357), .B2(new_n352), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n233), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n349), .A2(new_n351), .A3(new_n358), .A4(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G113), .B(G122), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT77), .B(G104), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n362), .A2(new_n363), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n363), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n355), .A2(new_n356), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n233), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n357), .A2(G146), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n345), .A2(new_n347), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT18), .B(G131), .C1(new_n339), .C2(new_n340), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n361), .A2(new_n371), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n341), .A2(new_n348), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT19), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n372), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n357), .A2(KEYINPUT19), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n381), .B(new_n358), .C1(G146), .C2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n371), .B1(new_n379), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n332), .B(new_n287), .C1(new_n380), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT20), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n361), .A2(new_n371), .A3(new_n379), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n386), .A2(new_n379), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(new_n371), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT20), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n332), .A4(new_n287), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n361), .A2(new_n379), .ZN(new_n396));
  INV_X1    g210(.A(new_n371), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT79), .A3(new_n390), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n400), .A3(new_n397), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n287), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G475), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n264), .A2(G952), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(G234), .B2(G237), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI211_X1 g220(.A(new_n287), .B(new_n264), .C1(G234), .C2(G237), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT21), .B(G898), .Z(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n410), .B(KEYINPUT81), .Z(new_n411));
  NAND4_X1  g225(.A1(new_n331), .A2(new_n395), .A3(new_n403), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n389), .A2(new_n394), .B1(new_n402), .B2(G475), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(KEYINPUT82), .A3(new_n331), .A4(new_n411), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G469), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n261), .B1(new_n239), .B2(new_n258), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n204), .A2(new_n419), .A3(new_n215), .ZN(new_n420));
  INV_X1    g234(.A(new_n248), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT1), .B1(new_n236), .B2(G146), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n422), .A2(G128), .B1(new_n234), .B2(new_n246), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n203), .B(new_n219), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n298), .B2(G137), .ZN(new_n428));
  INV_X1    g242(.A(G137), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT11), .A3(G134), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n298), .A2(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G131), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n346), .A2(new_n430), .A3(new_n431), .A4(new_n428), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n248), .B1(new_n253), .B2(new_n241), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n220), .A2(new_n437), .A3(KEYINPUT10), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n420), .A2(new_n426), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n264), .A2(G227), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(G140), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT71), .B(G110), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n424), .B1(new_n437), .B2(new_n220), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT12), .A3(new_n435), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  INV_X1    g261(.A(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n448), .B2(new_n436), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n444), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n420), .A2(new_n426), .A3(new_n438), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n435), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n443), .B1(new_n452), .B2(new_n439), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n418), .B(new_n287), .C1(new_n450), .C2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n439), .A3(new_n443), .ZN(new_n455));
  INV_X1    g269(.A(new_n451), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n449), .A2(new_n446), .B1(new_n456), .B2(new_n436), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n455), .B(G469), .C1(new_n457), .C2(new_n443), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n418), .A2(new_n287), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n454), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G221), .ZN(new_n462));
  INV_X1    g276(.A(new_n316), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n287), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n292), .A2(new_n417), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n205), .A2(G128), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT23), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT23), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n205), .B2(G128), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G119), .B(G128), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT24), .B(G110), .Z(new_n478));
  OAI22_X1  g292(.A1(new_n476), .A2(G110), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n358), .A3(new_n373), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT70), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n360), .A2(new_n358), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n477), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n476), .B(KEYINPUT69), .ZN(new_n485));
  INV_X1    g299(.A(G110), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n480), .A2(new_n481), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT22), .B(G137), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n482), .A2(new_n487), .A3(new_n488), .A4(new_n492), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n471), .B1(new_n496), .B2(G902), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(KEYINPUT25), .A3(new_n287), .A4(new_n495), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n317), .B1(G234), .B2(new_n287), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n419), .A2(new_n435), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n429), .A2(G134), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n333), .B1(new_n506), .B2(new_n431), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(new_n346), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n437), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n505), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n505), .B2(new_n510), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n213), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT26), .B(G101), .Z(new_n515));
  NAND2_X1  g329(.A1(new_n338), .A2(G210), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n435), .A2(new_n419), .B1(new_n509), .B2(new_n437), .ZN(new_n520));
  INV_X1    g334(.A(new_n213), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n514), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT31), .ZN(new_n524));
  INV_X1    g338(.A(new_n519), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n213), .B1(new_n520), .B2(KEYINPUT67), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n505), .A2(new_n510), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT28), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n213), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n522), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n525), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n514), .A2(new_n535), .A3(new_n519), .A4(new_n522), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G472), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n287), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT68), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OR3_X1    g358(.A1(new_n530), .A2(new_n533), .A3(new_n525), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n514), .A2(new_n522), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n545), .B(new_n546), .C1(new_n519), .C2(new_n547), .ZN(new_n548));
  OR4_X1    g362(.A1(new_n546), .A2(new_n530), .A3(new_n533), .A4(new_n525), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n287), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G472), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n504), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n292), .A2(new_n417), .A3(KEYINPUT83), .A4(new_n467), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n470), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G101), .ZN(G3));
  NAND2_X1  g369(.A1(new_n537), .A2(new_n287), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G472), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n539), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n504), .A2(new_n466), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n322), .A2(new_n560), .A3(new_n324), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT33), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT85), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(G478), .A4(new_n287), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n325), .A2(new_n326), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n561), .A2(G478), .A3(new_n287), .A4(new_n562), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT85), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n415), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT86), .ZN(new_n572));
  INV_X1    g386(.A(new_n187), .ZN(new_n573));
  INV_X1    g387(.A(new_n291), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n289), .A2(KEYINPUT84), .A3(new_n291), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n411), .A2(new_n559), .A3(new_n572), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT34), .B(G104), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G6));
  NAND2_X1  g396(.A1(new_n328), .A2(new_n330), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n415), .A2(new_n583), .A3(new_n411), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n559), .A3(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G107), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G9));
  OR2_X1    g401(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n489), .B(new_n588), .Z(new_n589));
  AOI22_X1  g403(.A1(new_n499), .A2(new_n500), .B1(new_n502), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n558), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n470), .A2(new_n553), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT37), .B(G110), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G12));
  OAI21_X1  g408(.A(new_n406), .B1(new_n408), .B2(G900), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n415), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n331), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OR3_X1    g412(.A1(new_n578), .A2(KEYINPUT87), .A3(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n539), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT32), .B1(new_n539), .B2(KEYINPUT68), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n551), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n590), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n602), .A2(new_n467), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT87), .B1(new_n578), .B2(new_n598), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G128), .ZN(G30));
  NAND2_X1  g421(.A1(new_n289), .A2(new_n291), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT38), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n415), .A2(new_n331), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n595), .B(KEYINPUT39), .Z(new_n612));
  NOR2_X1   g426(.A1(new_n466), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(KEYINPUT40), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n547), .A2(new_n525), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n532), .A2(new_n522), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n287), .B1(new_n619), .B2(new_n519), .ZN(new_n620));
  OAI21_X1  g434(.A(G472), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n544), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n603), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n573), .B1(new_n614), .B2(KEYINPUT40), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n616), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G143), .ZN(G45));
  AND3_X1   g440(.A1(new_n569), .A2(new_n570), .A3(new_n595), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n576), .A2(new_n627), .A3(new_n577), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT88), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n590), .B1(new_n544), .B2(new_n551), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT88), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n576), .A2(new_n627), .A3(new_n577), .A4(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n629), .A2(new_n630), .A3(new_n467), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT89), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT89), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n604), .A2(new_n635), .A3(new_n632), .A4(new_n629), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G146), .ZN(G48));
  NOR2_X1   g452(.A1(new_n450), .A2(new_n453), .ZN(new_n639));
  OAI21_X1  g453(.A(G469), .B1(new_n639), .B2(G902), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(new_n454), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(new_n465), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n578), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n552), .A3(new_n411), .A4(new_n572), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT90), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT41), .B(G113), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G15));
  NAND3_X1  g462(.A1(new_n644), .A2(new_n552), .A3(new_n584), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G116), .ZN(G18));
  NAND3_X1  g464(.A1(new_n644), .A2(new_n630), .A3(new_n417), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G119), .ZN(G21));
  AND3_X1   g466(.A1(new_n576), .A2(new_n577), .A3(new_n611), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n504), .A2(new_n558), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(new_n411), .A3(new_n654), .A4(new_n642), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G122), .ZN(G24));
  NOR3_X1   g470(.A1(new_n558), .A2(new_n590), .A3(KEYINPUT91), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT91), .B1(new_n558), .B2(new_n590), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n627), .A3(new_n644), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G125), .ZN(G27));
  INV_X1    g476(.A(new_n504), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n537), .A2(KEYINPUT32), .A3(new_n538), .A4(new_n287), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT94), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(KEYINPUT94), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n551), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n539), .A2(new_n541), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT95), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n539), .A2(KEYINPUT95), .A3(new_n541), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n663), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT96), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(KEYINPUT96), .B(new_n663), .C1(new_n667), .C2(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n289), .A2(new_n291), .A3(new_n187), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT92), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n461), .B2(new_n465), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n461), .A2(new_n679), .A3(new_n465), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n677), .A2(KEYINPUT42), .A3(new_n627), .A4(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n602), .A3(new_n663), .A4(new_n627), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT93), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT93), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G131), .ZN(G33));
  NAND3_X1  g506(.A1(new_n552), .A2(new_n597), .A3(new_n682), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT97), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G134), .ZN(G36));
  OAI21_X1  g509(.A(new_n455), .B1(new_n457), .B2(new_n443), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n455), .B(KEYINPUT45), .C1(new_n457), .C2(new_n443), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(G469), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT98), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT98), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n459), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(KEYINPUT99), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n454), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n703), .B2(KEYINPUT46), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT99), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n703), .B2(KEYINPUT46), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n706), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n711), .A2(new_n465), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n415), .B(KEYINPUT101), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n569), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n567), .B(new_n564), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n570), .B1(new_n715), .B2(new_n566), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n714), .B(KEYINPUT43), .C1(new_n716), .C2(KEYINPUT100), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n720), .A3(new_n558), .A4(new_n603), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n612), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n712), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n678), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n721), .A2(new_n727), .A3(new_n722), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n727), .B1(new_n721), .B2(new_n722), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT103), .B(G137), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT104), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n731), .B(new_n733), .ZN(G39));
  AND3_X1   g548(.A1(new_n711), .A2(KEYINPUT47), .A3(new_n465), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n711), .B2(new_n465), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n627), .B(new_n726), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n544), .A2(new_n551), .A3(new_n504), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n353), .ZN(G42));
  NOR2_X1   g554(.A1(new_n643), .A2(new_n678), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n622), .A2(new_n741), .A3(new_n663), .A4(new_n405), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n570), .A3(new_n569), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n717), .A2(new_n405), .A3(new_n720), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(new_n654), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n573), .A2(new_n745), .A3(new_n610), .A4(new_n642), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n746), .A2(KEYINPUT50), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(KEYINPUT50), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n744), .A2(new_n660), .A3(new_n741), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n735), .A2(new_n736), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT114), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n641), .A2(new_n464), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT115), .Z(new_n754));
  NOR2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n745), .A2(new_n726), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT113), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n749), .B(new_n750), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n677), .A2(new_n744), .A3(new_n741), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT48), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n404), .B(KEYINPUT116), .ZN(new_n762));
  INV_X1    g576(.A(new_n572), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n742), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n745), .B2(new_n644), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT117), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(KEYINPUT117), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n758), .A2(new_n759), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n623), .A2(new_n467), .A3(new_n595), .A4(new_n653), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n637), .A2(new_n606), .A3(new_n661), .A4(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n660), .A2(new_n627), .A3(new_n644), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n634), .B2(new_n636), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(KEYINPUT52), .A3(new_n606), .A4(new_n771), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n770), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n645), .A2(new_n651), .A3(new_n649), .A4(new_n655), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n415), .B1(new_n715), .B2(new_n566), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n608), .A2(new_n780), .A3(new_n411), .A4(new_n188), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT105), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT105), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n292), .A2(new_n783), .A3(new_n411), .A4(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n559), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n328), .A2(KEYINPUT106), .A3(new_n330), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT106), .B1(new_n328), .B2(new_n330), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n570), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n559), .A2(new_n411), .A3(new_n292), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n554), .A2(new_n592), .A3(new_n785), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n681), .A2(new_n680), .ZN(new_n793));
  INV_X1    g607(.A(new_n659), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n627), .B(new_n793), .C1(new_n794), .C2(new_n657), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n596), .A2(new_n788), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT107), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n602), .A3(new_n467), .A4(new_n603), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n678), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n779), .A2(new_n792), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n691), .A3(new_n694), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n778), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n772), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n801), .B1(new_n777), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n803), .B(new_n805), .C1(KEYINPUT53), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n777), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n802), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n813), .A2(new_n770), .B1(new_n778), .B2(new_n802), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(KEYINPUT112), .A3(new_n805), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT108), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n801), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n774), .A2(new_n777), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n800), .A2(new_n691), .A3(KEYINPUT108), .A4(new_n694), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n770), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n824));
  AOI211_X1 g638(.A(KEYINPUT110), .B(new_n817), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(KEYINPUT54), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n769), .B(new_n816), .C1(new_n825), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n749), .A2(new_n750), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n757), .B1(new_n751), .B2(new_n753), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n759), .A3(new_n831), .ZN(new_n832));
  OAI22_X1  g646(.A1(new_n829), .A2(new_n832), .B1(G952), .B2(G953), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n641), .B(KEYINPUT49), .Z(new_n834));
  NOR4_X1   g648(.A1(new_n609), .A2(new_n834), .A3(new_n504), .A4(new_n189), .ZN(new_n835));
  INV_X1    g649(.A(new_n714), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n465), .A3(new_n622), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(G75));
  XOR2_X1   g652(.A(new_n266), .B(KEYINPUT55), .Z(new_n839));
  OAI21_X1  g653(.A(new_n803), .B1(KEYINPUT53), .B2(new_n808), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(G210), .A3(G902), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n232), .B(KEYINPUT118), .Z(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n843), .B1(new_n841), .B2(new_n842), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n839), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n846), .ZN(new_n848));
  INV_X1    g662(.A(new_n839), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n264), .A2(G952), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n847), .A2(new_n850), .A3(new_n852), .ZN(G51));
  NAND2_X1  g667(.A1(new_n460), .A2(KEYINPUT57), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n460), .A2(KEYINPUT57), .ZN(new_n855));
  INV_X1    g669(.A(new_n809), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n814), .A2(new_n805), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n453), .B2(new_n450), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n840), .A2(G902), .A3(new_n701), .A4(new_n702), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(G54));
  AND4_X1   g675(.A1(KEYINPUT58), .A2(new_n840), .A3(G475), .A4(G902), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n392), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n392), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n851), .ZN(G60));
  OAI21_X1  g679(.A(new_n816), .B1(new_n828), .B2(new_n825), .ZN(new_n866));
  NAND2_X1  g680(.A1(G478), .A2(G902), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT59), .Z(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n563), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n563), .B1(new_n856), .B2(new_n857), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n868), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n851), .A3(new_n872), .ZN(G63));
  NAND2_X1  g687(.A1(G217), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT60), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n814), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  INV_X1    g691(.A(new_n875), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n778), .A2(new_n802), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n812), .B2(new_n802), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n876), .A2(new_n496), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n882), .A2(new_n852), .ZN(new_n883));
  INV_X1    g697(.A(new_n589), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n876), .B2(new_n881), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n883), .B(new_n886), .C1(KEYINPUT120), .C2(KEYINPUT61), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n882), .A2(KEYINPUT120), .A3(new_n852), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n852), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n885), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(G66));
  NOR2_X1   g706(.A1(new_n779), .A2(new_n792), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(G953), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n264), .B1(new_n409), .B2(G224), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT121), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(KEYINPUT121), .B2(new_n895), .ZN(new_n897));
  INV_X1    g711(.A(new_n843), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(G898), .B2(new_n264), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n897), .B(new_n899), .ZN(G69));
  NOR2_X1   g714(.A1(new_n512), .A2(new_n513), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n385), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n614), .A2(new_n678), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n552), .B(new_n903), .C1(new_n780), .C2(new_n790), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n737), .A2(new_n738), .B1(new_n730), .B2(new_n725), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n776), .A2(new_n606), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n776), .A2(new_n909), .A3(new_n606), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n625), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n905), .B(new_n906), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n902), .B1(new_n915), .B2(new_n264), .ZN(new_n916));
  NAND3_X1  g730(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(G227), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(G900), .A3(G953), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT123), .B1(new_n691), .B2(new_n694), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n906), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n691), .A2(KEYINPUT123), .A3(new_n694), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n712), .A2(new_n724), .A3(new_n653), .A4(new_n677), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n908), .A2(new_n910), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n922), .A2(KEYINPUT124), .A3(new_n923), .A4(new_n925), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n902), .B(new_n920), .C1(new_n930), .C2(G953), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n918), .A2(new_n931), .ZN(G72));
  INV_X1    g746(.A(new_n617), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n538), .A2(new_n287), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n547), .A2(new_n525), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n827), .A2(new_n933), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n936), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n915), .B2(new_n893), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n852), .B(new_n938), .C1(new_n940), .C2(new_n933), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n928), .A2(new_n893), .A3(new_n929), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n942), .A2(KEYINPUT126), .A3(new_n936), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT126), .B1(new_n942), .B2(new_n936), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n937), .B(KEYINPUT127), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(G57));
endmodule


