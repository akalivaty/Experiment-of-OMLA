//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G43gat), .ZN(new_n205));
  INV_X1    g004(.A(G43gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G50gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(KEYINPUT88), .A3(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT15), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT14), .B(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n213), .A2(new_n214), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n214), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n219), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n223), .A2(KEYINPUT89), .A3(new_n211), .A4(new_n210), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G22gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G15gat), .ZN(new_n228));
  INV_X1    g027(.A(G15gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G22gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT91), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT16), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G8gat), .ZN(new_n239));
  INV_X1    g038(.A(G8gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n233), .A2(new_n235), .A3(new_n240), .A4(new_n237), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT17), .B1(new_n220), .B2(new_n225), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n222), .A2(new_n224), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n214), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n210), .A2(new_n211), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT89), .B1(new_n250), .B2(new_n223), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n222), .B1(new_n251), .B2(new_n221), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n242), .B1(new_n226), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n244), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G229gat), .A2(G233gat), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT18), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT92), .B1(new_n253), .B2(KEYINPUT17), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n246), .B(new_n263), .C1(new_n249), .C2(new_n252), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n258), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT18), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(G229gat), .B2(G233gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n243), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT93), .B1(new_n226), .B2(new_n242), .ZN(new_n269));
  INV_X1    g068(.A(new_n242), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n253), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n272), .A3(new_n243), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n260), .B(KEYINPUT13), .Z(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G113gat), .B(G141gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G197gat), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT11), .B(G169gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n280), .B(KEYINPUT12), .Z(new_n281));
  NOR3_X1   g080(.A1(new_n261), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n259), .A2(new_n267), .B1(new_n274), .B2(new_n273), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n265), .A2(new_n260), .A3(new_n243), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n266), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n202), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n281), .B1(new_n261), .B2(new_n276), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n284), .A2(new_n286), .A3(new_n283), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT94), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G141gat), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT78), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n302));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n298), .A2(new_n300), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n308), .A2(KEYINPUT79), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n313), .A2(new_n316), .A3(new_n320), .A4(new_n317), .ZN(new_n321));
  AOI211_X1 g120(.A(KEYINPUT80), .B(KEYINPUT3), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n305), .B1(new_n299), .B2(new_n306), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n298), .A2(new_n303), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT79), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n313), .B1(new_n316), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n321), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n322), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G134gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G127gat), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G134gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n333), .A2(KEYINPUT71), .A3(G127gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G120gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G113gat), .ZN(new_n342));
  INV_X1    g141(.A(G113gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G120gat), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT1), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT72), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n338), .A4(new_n339), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n334), .A2(new_n336), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n330), .B2(new_n329), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT81), .B1(new_n332), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n330), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT80), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n329), .A2(new_n323), .A3(new_n330), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n346), .A2(new_n349), .B1(new_n345), .B2(new_n351), .ZN(new_n360));
  INV_X1    g159(.A(new_n329), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(KEYINPUT3), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n329), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n360), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n365), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n353), .A2(new_n361), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n367), .ZN(new_n376));
  INV_X1    g175(.A(new_n366), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G1gat), .B(G29gat), .Z(new_n381));
  XNOR2_X1  g180(.A(G57gat), .B(G85gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n365), .A2(KEYINPUT5), .A3(new_n366), .A4(new_n372), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n380), .A2(KEYINPUT6), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  AOI211_X1 g187(.A(new_n377), .B(new_n371), .C1(new_n355), .C2(new_n364), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n387), .B(new_n386), .C1(new_n389), .C2(new_n378), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n380), .B2(new_n387), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(G211gat), .B(G218gat), .Z(new_n395));
  NAND2_X1  g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(G197gat), .A2(G204gat), .ZN(new_n399));
  AND2_X1   g198(.A1(G197gat), .A2(G204gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n395), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n395), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(KEYINPUT74), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  AND2_X1   g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(KEYINPUT23), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n413));
  OR2_X1    g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT23), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n411), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n417));
  OAI211_X1 g216(.A(KEYINPUT25), .B(new_n412), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT67), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  INV_X1    g221(.A(G183gat), .ZN(new_n423));
  INV_X1    g222(.A(G190gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n421), .A2(new_n422), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n418), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT66), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT25), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT64), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n425), .B(new_n426), .C1(new_n419), .C2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n419), .A2(new_n433), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n429), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(KEYINPUT66), .B(new_n431), .C1(new_n432), .C2(new_n436), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT27), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G183gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n423), .A2(KEYINPUT27), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(G190gat), .B1(new_n442), .B2(KEYINPUT68), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n440), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT28), .A4(new_n424), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT70), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n440), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n423), .A2(KEYINPUT27), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n424), .B1(new_n453), .B2(new_n445), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT68), .B1(new_n442), .B2(new_n443), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n449), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n423), .A2(new_n424), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT26), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n460), .B(new_n461), .C1(KEYINPUT26), .C2(new_n411), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n438), .A2(new_n439), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n409), .B1(new_n463), .B2(KEYINPUT29), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n437), .A2(new_n430), .ZN(new_n465));
  INV_X1    g264(.A(new_n429), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n439), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n456), .A2(new_n457), .A3(new_n449), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n457), .B1(new_n456), .B2(new_n449), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n409), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT76), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT76), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n474), .B(new_n409), .C1(new_n467), .C2(new_n470), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n408), .B(new_n464), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n472), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n409), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n407), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G8gat), .B(G36gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT77), .ZN(new_n484));
  XNOR2_X1  g283(.A(G64gat), .B(G92gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n486), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n476), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n476), .A2(new_n481), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n488), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n394), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n477), .B1(new_n357), .B2(new_n358), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(new_n408), .ZN(new_n497));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT29), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT3), .B1(new_n408), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n501), .B2(new_n329), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n477), .B1(new_n405), .B2(new_n401), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n402), .A2(new_n395), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT3), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n496), .A2(new_n408), .B1(new_n329), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n509), .B2(new_n498), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n329), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n478), .B1(new_n322), .B2(new_n331), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n407), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n499), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n227), .B(new_n504), .C1(new_n510), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n516));
  XNOR2_X1  g315(.A(G78gat), .B(G106gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G50gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n509), .A2(new_n505), .A3(new_n498), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT83), .B1(new_n513), .B2(new_n499), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n503), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT85), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n227), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n519), .A2(KEYINPUT84), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n522), .B2(new_n227), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n504), .B1(new_n510), .B2(new_n514), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G22gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n522), .A2(new_n227), .A3(new_n526), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n495), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT36), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n471), .A2(new_n360), .ZN(new_n539));
  INV_X1    g338(.A(G227gat), .ZN(new_n540));
  INV_X1    g339(.A(G233gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n467), .A2(new_n353), .A3(new_n470), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G15gat), .B(G43gat), .Z(new_n547));
  XNOR2_X1  g346(.A(G71gat), .B(G99gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n539), .A2(new_n543), .ZN(new_n551));
  INV_X1    g350(.A(new_n542), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT34), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT34), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n551), .B2(new_n552), .ZN(new_n558));
  AOI211_X1 g357(.A(KEYINPUT34), .B(new_n542), .C1(new_n539), .C2(new_n543), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n546), .B(new_n549), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n544), .A2(KEYINPUT32), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n557), .B2(new_n560), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n537), .B(new_n538), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n557), .A2(new_n560), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n561), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(KEYINPUT73), .A3(new_n536), .A4(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n490), .A2(new_n390), .A3(new_n493), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT39), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n332), .A2(new_n354), .A3(KEYINPUT81), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n363), .B1(new_n359), .B2(new_n362), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n372), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT86), .B1(new_n575), .B2(new_n377), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n371), .B1(new_n355), .B2(new_n364), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n577), .A2(new_n578), .A3(new_n366), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n572), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(KEYINPUT86), .A3(new_n377), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n578), .B1(new_n577), .B2(new_n366), .ZN(new_n582));
  INV_X1    g381(.A(new_n376), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n572), .B1(new_n583), .B2(new_n366), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n385), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT40), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n580), .A2(KEYINPUT40), .A3(new_n385), .A4(new_n585), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n534), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT87), .B1(new_n392), .B2(new_n393), .ZN(new_n593));
  INV_X1    g392(.A(new_n387), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n378), .B1(new_n577), .B2(new_n366), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n385), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n596), .A2(new_n597), .A3(new_n391), .A4(new_n390), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(new_n598), .A3(new_n388), .ZN(new_n599));
  INV_X1    g398(.A(new_n489), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n488), .B1(new_n491), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n479), .A2(new_n480), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n603), .B2(new_n408), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n407), .B(new_n464), .C1(new_n473), .C2(new_n475), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT38), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n600), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n491), .A2(new_n601), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n486), .B1(new_n482), .B2(KEYINPUT37), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT38), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n599), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n535), .B(new_n570), .C1(new_n592), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n567), .A2(new_n568), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n495), .A2(new_n534), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n563), .A2(new_n564), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n532), .B1(new_n530), .B2(new_n528), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n617), .A2(new_n494), .A3(new_n525), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n616), .ZN(new_n620));
  OAI22_X1  g419(.A1(new_n615), .A2(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n295), .B1(new_n613), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G57gat), .B(G64gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT9), .ZN(new_n624));
  NAND2_X1  g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n625), .B(new_n627), .C1(new_n623), .C2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G127gat), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n270), .B1(new_n632), .B2(new_n631), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n309), .ZN(new_n640));
  XOR2_X1   g439(.A(G183gat), .B(G211gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G99gat), .B(G106gat), .Z(new_n647));
  NAND2_X1  g446(.A1(G85gat), .A2(G92gat), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT7), .B1(new_n648), .B2(KEYINPUT96), .ZN(new_n649));
  NAND2_X1  g448(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n650), .A2(new_n651), .A3(G85gat), .A4(G92gat), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G99gat), .ZN(new_n654));
  INV_X1    g453(.A(G106gat), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT8), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT95), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(G85gat), .ZN(new_n659));
  INV_X1    g458(.A(G92gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n647), .B1(new_n653), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n656), .A2(new_n658), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n652), .ZN(new_n666));
  INV_X1    g465(.A(new_n647), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n226), .B2(new_n257), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n255), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(G190gat), .B(G218gat), .Z(new_n673));
  NAND2_X1  g472(.A1(G232gat), .A2(G233gat), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n226), .A2(new_n670), .B1(KEYINPUT41), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n672), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n675), .A2(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g478(.A(G134gat), .B(G162gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n673), .B1(new_n672), .B2(new_n677), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n678), .B2(new_n682), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n663), .A2(new_n668), .A3(new_n629), .A4(new_n630), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT10), .B1(new_n687), .B2(KEYINPUT97), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G230gat), .A2(G233gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n631), .B1(new_n664), .B2(new_n669), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(KEYINPUT97), .A3(KEYINPUT10), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n687), .ZN(new_n694));
  INV_X1    g493(.A(new_n690), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(G120gat), .B(G148gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT98), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n693), .A2(new_n696), .A3(new_n701), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n646), .A2(new_n686), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n622), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n394), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G1gat), .ZN(G1324gat));
  INV_X1    g510(.A(new_n494), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT16), .B(G8gat), .Z(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT99), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(G8gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(G1325gat));
  INV_X1    g519(.A(new_n708), .ZN(new_n721));
  OAI21_X1  g520(.A(G15gat), .B1(new_n721), .B2(new_n570), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n708), .A2(new_n229), .A3(new_n617), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n534), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT43), .B(G22gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  INV_X1    g526(.A(new_n646), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n705), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n686), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n622), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n709), .A2(new_n218), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT100), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n735), .A2(KEYINPUT45), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT45), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n619), .ZN(new_n741));
  INV_X1    g540(.A(new_n388), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n596), .A2(new_n391), .A3(new_n390), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(KEYINPUT87), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT35), .B1(new_n744), .B2(new_n598), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n743), .A2(new_n388), .B1(new_n490), .B2(new_n493), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n746), .A2(new_n617), .A3(new_n525), .A4(new_n618), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n741), .A2(new_n745), .B1(new_n747), .B2(KEYINPUT35), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n565), .A2(new_n569), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n590), .A2(new_n591), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n744), .A2(new_n598), .A3(new_n610), .A4(new_n607), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n535), .A2(KEYINPUT102), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n495), .A2(new_n534), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n748), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n686), .B1(new_n613), .B2(new_n621), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n758), .A2(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT101), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n282), .B2(new_n287), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT101), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n729), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n709), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n218), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n740), .A2(new_n772), .ZN(G1328gat));
  NAND3_X1  g572(.A1(new_n731), .A2(new_n216), .A3(new_n712), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT46), .Z(new_n775));
  NAND3_X1  g574(.A1(new_n763), .A2(new_n712), .A3(new_n768), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n777), .B2(new_n216), .ZN(G1329gat));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n749), .A3(new_n768), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G43gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n731), .A2(new_n206), .A3(new_n617), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1330gat));
  NAND3_X1  g583(.A1(new_n763), .A2(new_n534), .A3(new_n768), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G50gat), .ZN(new_n786));
  NOR2_X1   g585(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n534), .A2(new_n204), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT104), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n731), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(G1331gat));
  NAND3_X1  g592(.A1(new_n751), .A2(new_n591), .A3(new_n590), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n794), .A2(new_n570), .A3(new_n755), .A4(new_n753), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n621), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n765), .A2(new_n766), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n728), .A2(new_n797), .A3(new_n685), .A4(new_n705), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n709), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT107), .B(G57gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(G1332gat));
  AOI21_X1  g603(.A(new_n494), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT108), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT109), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n806), .B(new_n809), .ZN(G1333gat));
  NOR2_X1   g609(.A1(new_n614), .A2(G71gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n801), .A2(new_n749), .ZN(new_n814));
  INV_X1    g613(.A(G71gat), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(new_n812), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n815), .B1(new_n801), .B2(new_n749), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(G1334gat));
  NAND2_X1  g620(.A1(new_n801), .A2(new_n534), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g622(.A1(new_n646), .A2(new_n797), .A3(new_n705), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n613), .A2(new_n621), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n762), .B1(new_n825), .B2(new_n685), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n760), .B1(new_n795), .B2(new_n621), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n709), .B(new_n824), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n763), .A2(KEYINPUT111), .A3(new_n709), .A4(new_n824), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(G85gat), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n646), .A2(new_n797), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n685), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n758), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n837));
  INV_X1    g636(.A(new_n835), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n796), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT51), .B1(new_n796), .B2(new_n838), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n833), .B(new_n835), .C1(new_n795), .C2(new_n621), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT112), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n709), .A2(new_n659), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n840), .A2(new_n843), .A3(new_n704), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n832), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n846), .A3(KEYINPUT113), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1336gat));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n839), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n712), .A2(new_n660), .A3(new_n704), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n763), .A2(new_n712), .A3(new_n824), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(G92gat), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n855), .B(KEYINPUT114), .Z(new_n859));
  AOI22_X1  g658(.A1(new_n857), .A2(G92gat), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n856), .A2(new_n858), .B1(new_n860), .B2(new_n852), .ZN(G1337gat));
  NAND3_X1  g660(.A1(new_n763), .A2(new_n749), .A3(new_n824), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G99gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n843), .A3(new_n704), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n617), .A2(new_n654), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(G1338gat));
  NAND4_X1  g665(.A1(new_n853), .A2(new_n655), .A3(new_n534), .A4(new_n704), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n763), .A2(new_n534), .A3(new_n824), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(G106gat), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n870), .B(new_n872), .ZN(G1339gat));
  NOR2_X1   g672(.A1(new_n706), .A2(new_n797), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n692), .A2(new_n691), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n695), .A3(new_n688), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n701), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n695), .B1(new_n875), .B2(new_n688), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n693), .A3(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(KEYINPUT55), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n703), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(KEYINPUT116), .A3(new_n703), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT55), .B1(new_n878), .B2(new_n880), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n259), .A2(new_n260), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n273), .A2(new_n274), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n280), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n291), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n686), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n291), .A2(new_n891), .A3(new_n704), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n797), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n686), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT117), .B(new_n896), .C1(new_n897), .C2(new_n797), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n894), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n874), .B1(new_n902), .B2(new_n728), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n394), .A3(new_n619), .ZN(new_n904));
  AOI21_X1  g703(.A(G113gat), .B1(new_n904), .B2(new_n797), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT118), .B1(new_n903), .B2(new_n534), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n895), .B1(new_n767), .B2(new_n888), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT117), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n898), .A2(new_n899), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n686), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n646), .B1(new_n911), .B2(new_n894), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n907), .B(new_n591), .C1(new_n912), .C2(new_n874), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n712), .A2(new_n394), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n617), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n295), .A2(new_n343), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n905), .B1(new_n917), .B2(new_n918), .ZN(G1340gat));
  AOI21_X1  g718(.A(G120gat), .B1(new_n904), .B2(new_n704), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n705), .A2(new_n341), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n917), .B2(new_n921), .ZN(G1341gat));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n335), .A3(new_n646), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n914), .A2(new_n728), .A3(new_n916), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n335), .ZN(G1342gat));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n333), .A3(new_n685), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT56), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n926), .A2(KEYINPUT56), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n914), .A2(new_n686), .A3(new_n916), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n333), .ZN(G1343gat));
  NOR2_X1   g729(.A1(new_n903), .A2(new_n394), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n749), .A2(new_n712), .A3(new_n591), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n294), .A2(new_n296), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n570), .A2(new_n915), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n591), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n882), .A2(new_n886), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n288), .A2(new_n292), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n895), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(KEYINPUT119), .A3(new_n895), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n686), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n893), .B1(new_n945), .B2(new_n946), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n646), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n938), .B1(new_n949), .B2(new_n874), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n937), .B1(new_n903), .B2(new_n591), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n936), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n797), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n935), .B1(new_n953), .B2(G141gat), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT58), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n296), .B1(new_n952), .B2(new_n294), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n933), .B2(new_n934), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n954), .A2(new_n955), .B1(new_n956), .B2(new_n957), .ZN(G1344gat));
  NAND2_X1  g757(.A1(new_n944), .A2(new_n686), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT119), .B1(new_n940), .B2(new_n895), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n894), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n728), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n706), .A2(new_n294), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n591), .B1(new_n965), .B2(KEYINPUT121), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT121), .B(new_n963), .C1(new_n961), .C2(new_n728), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT57), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n902), .A2(new_n728), .ZN(new_n970));
  INV_X1    g769(.A(new_n874), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n938), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n570), .A2(new_n704), .A3(new_n915), .ZN(new_n976));
  OAI211_X1 g775(.A(KEYINPUT59), .B(G148gat), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(KEYINPUT59), .B1(new_n933), .B2(new_n705), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n297), .ZN(new_n979));
  INV_X1    g778(.A(new_n952), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n705), .A2(KEYINPUT59), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n977), .B(new_n979), .C1(new_n980), .C2(new_n981), .ZN(G1345gat));
  OAI21_X1  g781(.A(G155gat), .B1(new_n980), .B2(new_n728), .ZN(new_n983));
  INV_X1    g782(.A(new_n933), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(new_n309), .A3(new_n646), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1346gat));
  OAI21_X1  g785(.A(G162gat), .B1(new_n980), .B2(new_n686), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n984), .A2(new_n310), .A3(new_n685), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1347gat));
  NAND2_X1  g788(.A1(new_n712), .A2(new_n394), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n990), .A2(new_n534), .A3(new_n614), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n903), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(G169gat), .B1(new_n993), .B2(new_n797), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n617), .A2(new_n394), .A3(new_n712), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n995), .B1(new_n906), .B2(new_n913), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n294), .A2(G169gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1348gat));
  INV_X1    g797(.A(G176gat), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n999), .B1(new_n996), .B2(new_n704), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT122), .ZN(new_n1001));
  NOR4_X1   g800(.A1(new_n903), .A2(G176gat), .A3(new_n705), .A4(new_n992), .ZN(new_n1002));
  OR3_X1    g801(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1001), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1349gat));
  NOR2_X1   g804(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n423), .B1(new_n996), .B2(new_n646), .ZN(new_n1007));
  NAND2_X1  g806(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n728), .A2(new_n444), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n972), .A2(new_n991), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1010), .A2(KEYINPUT123), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT123), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1012), .B1(new_n993), .B2(new_n1009), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1008), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1006), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1010), .A2(KEYINPUT123), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n993), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1017));
  AOI22_X1  g816(.A1(new_n1016), .A2(new_n1017), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n1018));
  INV_X1    g817(.A(new_n1006), .ZN(new_n1019));
  AOI211_X1 g818(.A(new_n728), .B(new_n995), .C1(new_n906), .C2(new_n913), .ZN(new_n1020));
  OAI211_X1 g819(.A(new_n1018), .B(new_n1019), .C1(new_n423), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g820(.A1(new_n1015), .A2(new_n1021), .ZN(G1350gat));
  AOI21_X1  g821(.A(new_n424), .B1(new_n996), .B2(new_n685), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n1023), .A2(KEYINPUT61), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(KEYINPUT61), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n993), .A2(new_n424), .A3(new_n685), .ZN(new_n1026));
  XOR2_X1   g825(.A(new_n1026), .B(KEYINPUT125), .Z(new_n1027));
  NAND3_X1  g826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(G1351gat));
  NAND3_X1  g827(.A1(new_n570), .A2(new_n712), .A3(new_n534), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n394), .B1(new_n1029), .B2(KEYINPUT126), .ZN(new_n1030));
  AOI211_X1 g829(.A(new_n1030), .B(new_n903), .C1(KEYINPUT126), .C2(new_n1029), .ZN(new_n1031));
  AOI21_X1  g830(.A(G197gat), .B1(new_n1031), .B2(new_n797), .ZN(new_n1032));
  NOR2_X1   g831(.A1(new_n749), .A2(new_n990), .ZN(new_n1033));
  INV_X1    g832(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g833(.A(new_n963), .B1(new_n961), .B2(new_n728), .ZN(new_n1035));
  INV_X1    g834(.A(KEYINPUT121), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n534), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g836(.A(new_n937), .B1(new_n1037), .B2(new_n967), .ZN(new_n1038));
  AOI21_X1  g837(.A(new_n1034), .B1(new_n1038), .B2(new_n973), .ZN(new_n1039));
  AND2_X1   g838(.A1(new_n294), .A2(G197gat), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(G1352gat));
  INV_X1    g840(.A(G204gat), .ZN(new_n1042));
  NAND3_X1  g841(.A1(new_n1031), .A2(new_n1042), .A3(new_n704), .ZN(new_n1043));
  OR2_X1    g842(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1044));
  NAND2_X1  g843(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1045));
  AND2_X1   g844(.A1(new_n1039), .A2(new_n704), .ZN(new_n1046));
  OAI211_X1 g845(.A(new_n1044), .B(new_n1045), .C1(new_n1046), .C2(new_n1042), .ZN(G1353gat));
  INV_X1    g846(.A(G211gat), .ZN(new_n1048));
  NAND3_X1  g847(.A1(new_n1031), .A2(new_n1048), .A3(new_n646), .ZN(new_n1049));
  INV_X1    g848(.A(KEYINPUT63), .ZN(new_n1050));
  AOI211_X1 g849(.A(new_n1050), .B(new_n1048), .C1(new_n1039), .C2(new_n646), .ZN(new_n1051));
  OAI211_X1 g850(.A(new_n646), .B(new_n1033), .C1(new_n969), .C2(new_n974), .ZN(new_n1052));
  AOI21_X1  g851(.A(KEYINPUT63), .B1(new_n1052), .B2(G211gat), .ZN(new_n1053));
  OAI21_X1  g852(.A(new_n1049), .B1(new_n1051), .B2(new_n1053), .ZN(G1354gat));
  INV_X1    g853(.A(G218gat), .ZN(new_n1055));
  AOI21_X1  g854(.A(new_n1055), .B1(new_n1039), .B2(new_n685), .ZN(new_n1056));
  NAND3_X1  g855(.A1(new_n1031), .A2(new_n1055), .A3(new_n685), .ZN(new_n1057));
  INV_X1    g856(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g857(.A(KEYINPUT127), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g858(.A(KEYINPUT127), .ZN(new_n1060));
  AOI211_X1 g859(.A(new_n686), .B(new_n1034), .C1(new_n1038), .C2(new_n973), .ZN(new_n1061));
  OAI211_X1 g860(.A(new_n1060), .B(new_n1057), .C1(new_n1061), .C2(new_n1055), .ZN(new_n1062));
  NAND2_X1  g861(.A1(new_n1059), .A2(new_n1062), .ZN(G1355gat));
endmodule


