//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT68), .B(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n191), .A2(new_n192), .A3(G143), .A4(G214), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT18), .A2(G131), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n197), .B2(new_n198), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n200), .B2(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT72), .B1(new_n207), .B2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G140), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT16), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  AOI21_X1  g027(.A(G146), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n213), .A3(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n208), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n195), .A2(new_n219), .A3(new_n196), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n195), .B2(new_n196), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND4_X1   g038(.A1(KEYINPUT87), .A2(new_n197), .A3(KEYINPUT17), .A4(G131), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT87), .B1(new_n221), .B2(KEYINPUT17), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n204), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n197), .A2(G131), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n195), .A2(new_n219), .A3(new_n196), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n223), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n197), .A2(KEYINPUT17), .A3(G131), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n217), .B1(new_n214), .B2(new_n215), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n207), .A2(KEYINPUT72), .A3(G146), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n221), .A2(KEYINPUT87), .A3(KEYINPUT17), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n235), .A2(new_n238), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n204), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n231), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n231), .A3(new_n244), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT88), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n232), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(G475), .B1(new_n249), .B2(G902), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G122), .ZN(new_n252));
  INV_X1    g066(.A(G122), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G116), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G107), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n194), .A2(KEYINPUT13), .A3(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(G128), .B2(new_n194), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT13), .B1(new_n194), .B2(G128), .ZN(new_n260));
  OAI21_X1  g074(.A(G134), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G128), .B(G143), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(KEYINPUT90), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT90), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n257), .A2(new_n261), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n262), .B(new_n263), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n252), .A2(KEYINPUT14), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n254), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n252), .A2(KEYINPUT14), .ZN(new_n272));
  OAI21_X1  g086(.A(G107), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n255), .A2(new_n256), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n269), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT70), .B(G217), .Z(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT9), .B(G234), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n276), .A2(G953), .A3(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n268), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n268), .B2(new_n275), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT15), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(G478), .ZN(new_n285));
  INV_X1    g099(.A(G478), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n281), .B(new_n282), .C1(KEYINPUT15), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(G234), .A2(G237), .ZN(new_n289));
  INV_X1    g103(.A(G953), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n289), .A2(G952), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n192), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(G902), .A3(new_n289), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n293), .B(KEYINPUT91), .Z(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT21), .B(G898), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT92), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n200), .B(KEYINPUT19), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n201), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n217), .B(new_n302), .C1(new_n220), .C2(new_n221), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n231), .B1(new_n244), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n245), .B1(new_n228), .B2(new_n231), .ZN(new_n306));
  INV_X1    g120(.A(new_n246), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G475), .A2(G902), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT89), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n300), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n304), .B1(new_n248), .B2(new_n246), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n313), .A2(KEYINPUT20), .A3(new_n310), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n250), .B(new_n299), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT93), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n308), .A2(new_n317), .A3(new_n311), .ZN(new_n318));
  INV_X1    g132(.A(new_n300), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n313), .B2(new_n310), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT93), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n250), .A4(new_n299), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n201), .A2(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n194), .A2(G146), .ZN(new_n329));
  AND4_X1   g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(G128), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n331), .A2(G128), .B1(new_n328), .B2(new_n329), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n205), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n335));
  NOR2_X1   g149(.A1(KEYINPUT0), .A2(G128), .ZN(new_n336));
  XNOR2_X1  g150(.A(G143), .B(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(KEYINPUT0), .A2(G128), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n329), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT0), .A3(G128), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n334), .B(new_n335), .C1(new_n205), .C2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT82), .A4(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n290), .A2(G224), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n345), .B(new_n346), .Z(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n230), .B2(G107), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n256), .A2(KEYINPUT3), .A3(G104), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT74), .B1(new_n256), .B2(G104), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n230), .A3(G107), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G101), .ZN(new_n356));
  INV_X1    g170(.A(G101), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n351), .A2(new_n357), .A3(new_n352), .A4(new_n354), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n251), .A2(G119), .ZN(new_n360));
  INV_X1    g174(.A(G119), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT66), .B1(new_n361), .B2(G116), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT66), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n251), .A3(G119), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT2), .B(G113), .Z(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n352), .A2(new_n354), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n357), .B1(new_n368), .B2(new_n351), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n359), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n230), .A2(G107), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n256), .A2(G104), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n358), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n378));
  INV_X1    g192(.A(G113), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n360), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n378), .A2(new_n381), .B1(new_n365), .B2(new_n366), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n358), .A2(new_n383), .A3(new_n375), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n387));
  XNOR2_X1  g201(.A(G110), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n386), .A2(KEYINPUT81), .A3(new_n387), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n387), .B1(new_n386), .B2(new_n389), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n372), .A2(new_n385), .A3(new_n388), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n347), .B(new_n394), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT7), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n346), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n345), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n345), .A2(KEYINPUT84), .A3(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n388), .B(KEYINPUT8), .Z(new_n408));
  INV_X1    g222(.A(new_n382), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n376), .A2(KEYINPUT83), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n376), .A2(KEYINPUT83), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n382), .B1(KEYINPUT83), .B2(new_n376), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n343), .B(new_n344), .C1(new_n401), .C2(new_n346), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n414), .A2(new_n397), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n400), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G210), .B1(G237), .B2(G902), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n419), .B(KEYINPUT85), .Z(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n420), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n400), .A2(new_n417), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n326), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT76), .B1(new_n376), .B2(new_n333), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n331), .A2(G128), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n340), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n337), .A2(G128), .A3(new_n331), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT76), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n358), .A4(new_n375), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n376), .A2(new_n333), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G137), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT64), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT64), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G137), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT11), .A4(G134), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT11), .A2(G134), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT11), .A2(G134), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(G137), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n441), .A2(new_n219), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n219), .B1(new_n441), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n426), .B1(new_n436), .B2(new_n448), .ZN(new_n449));
  AOI211_X1 g263(.A(KEYINPUT12), .B(new_n447), .C1(new_n434), .C2(new_n435), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n192), .A2(G227), .ZN(new_n452));
  XOR2_X1   g266(.A(G110), .B(G140), .Z(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT78), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT10), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n333), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n377), .A2(new_n458), .A3(new_n384), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n369), .A2(new_n370), .B1(new_n341), .B2(new_n339), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n359), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT10), .B1(new_n427), .B2(new_n433), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n456), .B1(new_n464), .B2(new_n447), .ZN(new_n465));
  NOR4_X1   g279(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT78), .A4(new_n448), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n451), .B(new_n455), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n434), .A2(new_n457), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n469), .A2(new_n447), .A3(new_n459), .A4(new_n461), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n464), .A2(new_n456), .A3(new_n447), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n448), .B1(new_n462), .B2(new_n463), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT79), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT79), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n476), .B(new_n448), .C1(new_n462), .C2(new_n463), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n455), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n425), .B(new_n282), .C1(new_n468), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n473), .A2(new_n451), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n454), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n473), .A2(new_n478), .A3(new_n455), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(G469), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n425), .A2(new_n282), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G221), .B1(new_n277), .B2(G902), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n424), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n324), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT73), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT24), .B(G110), .Z(new_n492));
  XNOR2_X1  g306(.A(G119), .B(G128), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n361), .A2(G128), .ZN(new_n496));
  INV_X1    g310(.A(G128), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT23), .A3(G119), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n361), .A2(G128), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n496), .B(new_n498), .C1(new_n499), .C2(KEYINPUT23), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n495), .B1(new_n500), .B2(G110), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n495), .A3(G110), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n218), .B(new_n494), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  OAI22_X1  g318(.A1(new_n500), .A2(G110), .B1(new_n492), .B2(new_n493), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n200), .A2(new_n201), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n217), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G137), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n494), .B1(new_n503), .B2(new_n501), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n507), .B1(new_n241), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n515), .A3(new_n282), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n511), .A2(new_n515), .A3(KEYINPUT25), .A4(new_n282), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n276), .B1(G234), .B2(new_n282), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n515), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n521), .A2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n491), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n521), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n518), .B2(new_n519), .ZN(new_n529));
  INV_X1    g343(.A(new_n526), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT73), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  INV_X1    g347(.A(new_n367), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n438), .A2(new_n440), .A3(new_n263), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n219), .B1(G134), .B2(G137), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT65), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(KEYINPUT65), .A3(new_n536), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n441), .A2(new_n219), .A3(new_n444), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n431), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n342), .B1(new_n445), .B2(new_n446), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n367), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n534), .A2(new_n542), .A3(new_n543), .A4(KEYINPUT28), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n191), .A2(new_n192), .A3(G210), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n551), .A2(KEYINPUT27), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(KEYINPUT27), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT26), .B(G101), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n533), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n542), .A2(new_n543), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n542), .B2(new_n543), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n367), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n557), .B1(new_n563), .B2(new_n544), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n282), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT69), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n548), .A2(new_n566), .A3(new_n544), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n547), .A2(KEYINPUT69), .A3(new_n367), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(KEYINPUT28), .A3(new_n568), .ZN(new_n569));
  AND4_X1   g383(.A1(KEYINPUT29), .A2(new_n569), .A3(new_n557), .A4(new_n546), .ZN(new_n570));
  OAI21_X1  g384(.A(G472), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n563), .A2(new_n557), .A3(new_n544), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n550), .A2(new_n558), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT31), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n563), .A2(new_n575), .A3(new_n557), .A4(new_n544), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n578));
  NOR2_X1   g392(.A1(G472), .A2(G902), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n571), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n532), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n490), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  NAND2_X1  g400(.A1(new_n487), .A2(new_n488), .ZN(new_n587));
  INV_X1    g401(.A(new_n531), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n577), .A2(new_n579), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT73), .B1(new_n529), .B2(new_n530), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n577), .A2(new_n282), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n588), .A2(new_n589), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n281), .A2(new_n286), .A3(new_n282), .ZN(new_n595));
  NAND2_X1  g409(.A1(G478), .A2(G902), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n281), .B(KEYINPUT33), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n286), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n321), .B2(new_n250), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT94), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n421), .A2(new_n600), .A3(new_n423), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n422), .B1(new_n400), .B2(new_n417), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n326), .B1(new_n602), .B2(KEYINPUT94), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n297), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n594), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  NOR3_X1   g422(.A1(new_n313), .A2(new_n319), .A3(new_n310), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(KEYINPUT95), .A3(new_n320), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n612), .B1(new_n312), .B2(new_n609), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n611), .A2(new_n613), .A3(new_n250), .A4(new_n288), .ZN(new_n614));
  NOR4_X1   g428(.A1(new_n614), .A2(new_n604), .A3(new_n587), .A4(new_n593), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G107), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT96), .B(KEYINPUT35), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  XNOR2_X1  g432(.A(new_n513), .B(KEYINPUT97), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n619), .B(new_n620), .Z(new_n621));
  AOI21_X1  g435(.A(new_n529), .B1(new_n621), .B2(new_n525), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n623), .A2(new_n589), .A3(new_n592), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n490), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  AND4_X1   g441(.A1(new_n582), .A2(new_n487), .A3(new_n488), .A4(new_n623), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n601), .A2(new_n603), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G900), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n291), .B1(new_n294), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n614), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  XOR2_X1   g449(.A(new_n632), .B(KEYINPUT39), .Z(new_n636));
  NAND3_X1  g450(.A1(new_n487), .A2(new_n488), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT40), .Z(new_n638));
  INV_X1    g452(.A(new_n423), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n602), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT38), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n563), .A2(new_n544), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n642), .A2(new_n558), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n567), .A2(new_n568), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n643), .B(new_n282), .C1(new_n557), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n581), .B2(new_n580), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n325), .A3(new_n622), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n250), .B1(new_n312), .B2(new_n314), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n288), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n641), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n638), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT98), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G143), .ZN(G45));
  INV_X1    g468(.A(new_n598), .ZN(new_n655));
  INV_X1    g469(.A(new_n632), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT99), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n599), .A2(new_n659), .A3(new_n656), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n630), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G146), .ZN(G48));
  OAI21_X1  g477(.A(new_n282), .B1(new_n468), .B2(new_n479), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G469), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n488), .A3(new_n480), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n583), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n605), .A3(new_n599), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT100), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n667), .A2(new_n605), .A3(new_n670), .A4(new_n599), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NOR4_X1   g488(.A1(new_n614), .A2(new_n604), .A3(new_n666), .A4(new_n583), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n251), .ZN(G18));
  NAND2_X1  g490(.A1(new_n601), .A2(new_n603), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n666), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n582), .A2(new_n623), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n324), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n678), .A2(new_n324), .A3(new_n682), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  AOI22_X1  g499(.A1(new_n472), .A2(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n467), .B1(new_n686), .B2(new_n455), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n687), .A2(new_n425), .A3(new_n282), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n425), .B1(new_n687), .B2(new_n282), .ZN(new_n689));
  INV_X1    g503(.A(new_n488), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT103), .B(G472), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n591), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT104), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n591), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n573), .A2(new_n576), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n557), .B1(new_n569), .B2(new_n546), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n579), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT102), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n701), .B(new_n579), .C1(new_n697), .C2(new_n698), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n694), .A2(new_n696), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n529), .A2(new_n530), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n691), .A2(new_n703), .A3(new_n704), .A4(new_n297), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n601), .A2(new_n649), .A3(new_n603), .A4(new_n288), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT105), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n706), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n700), .A2(new_n702), .ZN(new_n709));
  INV_X1    g523(.A(new_n696), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n695), .B1(new_n591), .B2(new_n692), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n704), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n666), .A2(new_n298), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n708), .A2(new_n714), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n707), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NOR2_X1   g533(.A1(new_n712), .A2(new_n622), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n661), .A2(new_n678), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT106), .B(G125), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G27));
  NOR2_X1   g537(.A1(new_n690), .A2(new_n326), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n639), .A2(new_n602), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n483), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n686), .A2(KEYINPUT107), .A3(new_n455), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(G469), .A3(new_n482), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n480), .A2(new_n486), .ZN(new_n733));
  OAI211_X1 g547(.A(KEYINPUT42), .B(new_n726), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n582), .A2(new_n704), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n421), .A2(new_n423), .A3(new_n724), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n480), .A2(new_n486), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n739), .B1(new_n740), .B2(new_n731), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n658), .A2(new_n660), .A3(new_n741), .A4(new_n584), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n738), .A2(new_n661), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n219), .ZN(G33));
  AND3_X1   g559(.A1(new_n633), .A2(new_n584), .A3(new_n741), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n263), .ZN(G36));
  NAND2_X1  g561(.A1(new_n640), .A2(new_n325), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n321), .A2(new_n250), .A3(new_n655), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT43), .Z(new_n750));
  AOI21_X1  g564(.A(new_n622), .B1(new_n589), .B2(new_n592), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n748), .B1(new_n752), .B2(KEYINPUT44), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(KEYINPUT44), .B2(new_n752), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n730), .A2(KEYINPUT45), .A3(new_n482), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n482), .A2(new_n483), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n425), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n485), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(KEYINPUT46), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n480), .B1(new_n760), .B2(KEYINPUT46), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n488), .A3(new_n636), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n754), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  NAND3_X1  g580(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n488), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n488), .B1(new_n761), .B2(new_n762), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n748), .A2(new_n532), .A3(new_n582), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n661), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n675), .B1(new_n707), .B2(new_n717), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n778), .A2(new_n684), .A3(new_n672), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n611), .A2(new_n613), .A3(new_n250), .ZN(new_n780));
  INV_X1    g594(.A(new_n748), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n285), .A2(KEYINPUT112), .A3(new_n287), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT112), .B1(new_n285), .B2(new_n287), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n783), .A3(new_n632), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n628), .A2(new_n780), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n658), .A2(new_n720), .A3(new_n660), .A4(new_n741), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n744), .A2(new_n746), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n297), .B(new_n325), .C1(new_n639), .C2(new_n602), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n587), .A2(new_n593), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n649), .A2(new_n655), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n321), .B(new_n250), .C1(new_n782), .C2(new_n783), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n599), .A2(KEYINPUT111), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n324), .B(new_n489), .C1(new_n584), .C2(new_n624), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n779), .A2(new_n788), .A3(new_n789), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n630), .B1(new_n661), .B2(new_n633), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n488), .A2(new_n647), .A3(new_n622), .A4(new_n656), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n708), .B(new_n806), .C1(new_n733), .C2(new_n732), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n721), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n805), .A2(new_n721), .A3(KEYINPUT52), .A4(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n798), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT113), .B1(new_n797), .B2(new_n798), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n778), .A2(new_n684), .A3(new_n672), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n789), .B1(new_n818), .B2(new_n788), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT115), .B(new_n777), .C1(new_n813), .C2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n818), .A3(new_n788), .ZN(new_n821));
  XOR2_X1   g635(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n779), .A2(new_n788), .A3(new_n803), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n812), .A3(new_n804), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT115), .B1(new_n827), .B2(new_n777), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT54), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n812), .A2(new_n818), .A3(KEYINPUT53), .A4(new_n788), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n830), .A2(KEYINPUT117), .B1(new_n821), .B2(new_n822), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  INV_X1    g646(.A(new_n825), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT53), .A4(new_n812), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n832), .A4(new_n835), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n750), .A2(new_n291), .A3(new_n714), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n641), .A2(new_n326), .A3(new_n691), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT119), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(KEYINPUT119), .A3(KEYINPUT50), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n532), .A2(new_n291), .ZN(new_n847));
  OR4_X1    g661(.A1(new_n647), .A2(new_n748), .A3(new_n666), .A4(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n649), .A3(new_n655), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n291), .A2(new_n750), .A3(new_n691), .A4(new_n781), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n720), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n845), .A2(KEYINPUT51), .A3(new_n846), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n688), .A2(new_n689), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n690), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n767), .A2(KEYINPUT120), .A3(new_n770), .A4(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n840), .A2(new_n748), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n767), .A2(new_n770), .A3(new_n854), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n852), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n845), .A2(new_n846), .A3(new_n851), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n856), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n736), .A2(new_n737), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n850), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT48), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n840), .A2(new_n677), .A3(new_n666), .ZN(new_n869));
  OAI211_X1 g683(.A(G952), .B(new_n290), .C1(new_n848), .C2(new_n793), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n861), .A2(new_n864), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n829), .A2(new_n838), .A3(new_n839), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT121), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n853), .B(KEYINPUT49), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n749), .A2(new_n647), .A3(new_n713), .A4(new_n725), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n641), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT110), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n877), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n192), .A2(G952), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT123), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n282), .B1(new_n831), .B2(new_n835), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n420), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n347), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n896), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n831), .A2(new_n835), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n836), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n485), .B(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n687), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n890), .A2(new_n759), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n887), .B1(new_n905), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n890), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n908), .A2(new_n313), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n313), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n887), .ZN(G60));
  NAND3_X1  g725(.A1(new_n829), .A2(new_n838), .A3(new_n839), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n596), .B(KEYINPUT59), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n597), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n902), .A2(new_n597), .A3(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n889), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  AND2_X1   g732(.A1(new_n900), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n621), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n888), .C1(new_n524), .C2(new_n919), .ZN(new_n921));
  XOR2_X1   g735(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G66));
  INV_X1    g737(.A(new_n295), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n290), .B1(new_n924), .B2(G224), .ZN(new_n925));
  INV_X1    g739(.A(new_n818), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n192), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n894), .B1(G898), .B2(new_n192), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n927), .B(new_n928), .Z(G69));
  AOI21_X1  g743(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n561), .A2(new_n562), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n301), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n292), .A2(G900), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n773), .B(KEYINPUT109), .ZN(new_n938));
  OR3_X1    g752(.A1(new_n764), .A2(new_n706), .A3(new_n865), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n744), .A2(new_n746), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n805), .A2(new_n721), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n765), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n937), .B1(new_n943), .B2(new_n192), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n653), .A2(new_n941), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT62), .Z(new_n947));
  NOR3_X1   g761(.A1(new_n637), .A2(new_n748), .A3(new_n583), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n795), .B2(new_n796), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n754), .B2(new_n764), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n947), .A2(new_n775), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n192), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n934), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n932), .B1(new_n945), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n935), .B1(new_n953), .B2(new_n192), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n957), .A2(new_n944), .A3(KEYINPUT126), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n931), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n945), .A2(new_n955), .A3(new_n932), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT126), .B1(new_n957), .B2(new_n944), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n930), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(G72));
  NAND2_X1  g777(.A1(new_n642), .A2(new_n558), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n943), .A2(new_n818), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  AOI21_X1  g781(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n887), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n947), .A2(new_n775), .A3(new_n952), .A4(new_n818), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n643), .B1(new_n970), .B2(new_n967), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n824), .A2(new_n828), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n643), .A2(new_n964), .A3(new_n967), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n975), .A2(new_n978), .ZN(G57));
endmodule


