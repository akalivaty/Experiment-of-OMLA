//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT67), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT69), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n465), .A2(new_n467), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(G114), .A2(G2104), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n464), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G102), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n463), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n492), .B(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n491), .A2(new_n494), .ZN(G164));
  AND2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  OAI211_X1 g072(.A(G50), .B(G543), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n503), .A3(G62), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n499), .B1(new_n508), .B2(G651), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n501), .B(new_n503), .C1(new_n496), .C2(new_n497), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n512), .A2(G88), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n509), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  AND2_X1   g093(.A1(new_n514), .A2(G63), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n496), .A2(new_n497), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n500), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(G651), .B1(new_n521), .B2(G51), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n512), .A2(G89), .A3(new_n515), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n524), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n523), .B1(new_n528), .B2(new_n530), .ZN(G168));
  XOR2_X1   g106(.A(KEYINPUT73), .B(G52), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n521), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n512), .A2(new_n515), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n533), .B1(new_n534), .B2(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT74), .Z(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n501), .A2(new_n503), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n543), .A2(G651), .B1(new_n521), .B2(G43), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n512), .A2(G81), .A3(new_n515), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND3_X1  g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT75), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(G188));
  NAND3_X1  g131(.A1(new_n512), .A2(G91), .A3(new_n515), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n541), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n521), .A2(KEYINPUT9), .A3(G53), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n513), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n557), .A2(new_n561), .A3(new_n562), .A4(new_n566), .ZN(G299));
  XNOR2_X1  g142(.A(new_n538), .B(KEYINPUT74), .ZN(G301));
  AND3_X1   g143(.A1(new_n524), .A2(new_n529), .A3(new_n526), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n529), .B1(new_n524), .B2(new_n526), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n522), .B1(new_n569), .B2(new_n570), .ZN(G286));
  NAND3_X1  g146(.A1(new_n512), .A2(G87), .A3(new_n515), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n521), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n512), .A2(G86), .A3(new_n515), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n521), .A2(G48), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n541), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(new_n577), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n541), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n512), .A2(G85), .A3(new_n515), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n521), .A2(G47), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n589), .A2(KEYINPUT78), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n588), .A2(new_n595), .ZN(G290));
  NAND3_X1  g171(.A1(new_n512), .A2(G92), .A3(new_n515), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n541), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n521), .B2(G54), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n512), .A2(new_n515), .A3(new_n603), .A4(G92), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G284));
  OAI21_X1  g183(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G321));
  NAND2_X1  g184(.A1(G299), .A2(new_n606), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G168), .B2(new_n606), .ZN(G280));
  XNOR2_X1  g186(.A(G280), .B(KEYINPUT79), .ZN(G297));
  AND3_X1   g187(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n613));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n468), .A2(new_n489), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(G2100), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n477), .A2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n479), .A2(G135), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT82), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n645), .A2(G14), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2100), .Z(new_n654));
  AND2_X1   g229(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n650), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT83), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n662), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(new_n665), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n667), .C2(new_n669), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(G1986), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT22), .B(G1981), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  MUX2_X1   g255(.A(G6), .B(G305), .S(G16), .Z(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT32), .B(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(G16), .A2(G23), .ZN(new_n685));
  INV_X1    g260(.A(G288), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n684), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT34), .Z(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n587), .B1(new_n593), .B2(new_n594), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G16), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n700));
  OR2_X1    g275(.A1(G16), .A2(G24), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n697), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(G1986), .A3(new_n702), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n477), .A2(G119), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n468), .A2(G131), .A3(new_n463), .ZN(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n709), .B1(new_n714), .B2(new_n708), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n705), .A2(new_n707), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n715), .A2(new_n716), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n696), .A2(new_n718), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n705), .A2(new_n707), .A3(new_n720), .A4(new_n717), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n695), .B(KEYINPUT34), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT36), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n690), .A2(G19), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n547), .B2(new_n690), .ZN(new_n727));
  INV_X1    g302(.A(G1341), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT31), .B(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n477), .A2(G129), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n479), .A2(G141), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n489), .A2(G105), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(G29), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G29), .B2(G32), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G28), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(new_n745), .A3(new_n708), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n729), .A2(new_n730), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n748));
  INV_X1    g323(.A(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT91), .Z(new_n751));
  OR2_X1    g326(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(G29), .B2(G160), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(G2084), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n629), .A2(new_n708), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n747), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n739), .A2(new_n741), .B1(new_n753), .B2(G2084), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n489), .A2(G103), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT25), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n479), .A2(G139), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n760), .A2(KEYINPUT88), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(KEYINPUT88), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(G115), .A2(G2104), .ZN(new_n764));
  INV_X1    g339(.A(G127), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n476), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G2105), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(KEYINPUT89), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(KEYINPUT89), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n762), .A2(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G29), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n708), .A2(G33), .ZN(new_n772));
  AOI21_X1  g347(.A(G2072), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  INV_X1    g349(.A(new_n772), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n774), .B(new_n775), .C1(new_n770), .C2(G29), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n757), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(KEYINPUT93), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(new_n757), .C1(new_n773), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n708), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n708), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT29), .B(G2090), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n690), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n690), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1961), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n756), .A2(new_n781), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G21), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G168), .B2(G16), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G1966), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n787), .A2(G1961), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n690), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n613), .B2(new_n690), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT87), .B(G1348), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n795), .B(new_n796), .Z(new_n797));
  NOR4_X1   g372(.A1(new_n789), .A2(new_n792), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n708), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n708), .ZN(new_n800));
  INV_X1    g375(.A(G2078), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n791), .A2(G1966), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n725), .A2(new_n798), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n805));
  INV_X1    g380(.A(G26), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G29), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(G29), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n477), .A2(G128), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n479), .A2(G140), .ZN(new_n810));
  OR2_X1    g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n808), .B1(new_n813), .B2(G29), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n807), .B1(new_n814), .B2(new_n805), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n690), .A2(KEYINPUT23), .A3(G20), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT23), .ZN(new_n818));
  INV_X1    g393(.A(G20), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G16), .ZN(new_n820));
  INV_X1    g395(.A(G299), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n817), .B(new_n820), .C1(new_n821), .C2(new_n690), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT94), .B(G1956), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n804), .A2(new_n816), .A3(new_n824), .ZN(G311));
  AND3_X1   g400(.A1(new_n725), .A2(new_n798), .A3(new_n803), .ZN(new_n826));
  INV_X1    g401(.A(new_n816), .ZN(new_n827));
  INV_X1    g402(.A(new_n824), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n802), .ZN(G150));
  XOR2_X1   g404(.A(KEYINPUT96), .B(G860), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n541), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n834), .A2(G651), .B1(new_n521), .B2(G55), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n512), .A2(G93), .A3(new_n515), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n605), .A2(new_n614), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n512), .A2(G93), .A3(new_n515), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  INV_X1    g418(.A(G55), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n843), .A2(new_n534), .B1(new_n844), .B2(new_n564), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n545), .B(new_n544), .C1(new_n842), .C2(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n512), .A2(G81), .A3(new_n515), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n513), .A2(G43), .A3(G543), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n534), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n836), .B(new_n835), .C1(new_n847), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n841), .B(new_n852), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT97), .Z(new_n855));
  OAI21_X1  g430(.A(new_n831), .B1(new_n853), .B2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n838), .B1(new_n855), .B2(new_n856), .ZN(G145));
  INV_X1    g432(.A(new_n621), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  OR2_X1    g434(.A1(G106), .A2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(G118), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n464), .B1(new_n861), .B2(G2105), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n477), .A2(G130), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n468), .A2(G142), .A3(new_n463), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n479), .A2(new_n866), .A3(G142), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n863), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n714), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n870), .A2(new_n863), .A3(new_n865), .A4(new_n867), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n859), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n871), .A3(new_n859), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n858), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n876), .A2(new_n872), .A3(new_n621), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT103), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n621), .B1(new_n876), .B2(new_n872), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(new_n858), .A3(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n770), .A2(KEYINPUT100), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n884), .B1(new_n768), .B2(new_n769), .C1(new_n762), .C2(new_n763), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n734), .A2(new_n737), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G164), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n813), .A2(KEYINPUT99), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n809), .A2(new_n810), .A3(new_n890), .A4(new_n812), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n492), .B(KEYINPUT4), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n488), .A3(new_n490), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n734), .A3(new_n737), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n888), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n892), .B1(new_n888), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n886), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n888), .A2(new_n892), .A3(new_n895), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n883), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n878), .A2(new_n882), .A3(new_n898), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n879), .A2(new_n880), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(KEYINPUT103), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(G160), .B(KEYINPUT98), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(new_n483), .ZN(new_n907));
  INV_X1    g482(.A(new_n629), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n483), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n902), .A2(new_n905), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n902), .A2(new_n905), .ZN(new_n915));
  INV_X1    g490(.A(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT105), .B(G37), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n902), .A2(new_n905), .A3(new_n912), .A4(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n914), .A2(new_n917), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g497(.A(new_n606), .B1(new_n842), .B2(new_n845), .ZN(new_n923));
  NAND4_X1  g498(.A1(G303), .A2(new_n577), .A3(new_n576), .A4(new_n581), .ZN(new_n924));
  NAND3_X1  g499(.A1(G305), .A2(new_n516), .A3(new_n509), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(G288), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G288), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n927), .A2(new_n928), .A3(G290), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n686), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n698), .B1(new_n931), .B2(new_n926), .ZN(new_n932));
  NOR4_X1   g507(.A1(new_n929), .A2(new_n932), .A3(KEYINPUT109), .A4(KEYINPUT42), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n929), .B2(new_n932), .ZN(new_n935));
  OAI21_X1  g510(.A(G290), .B1(new_n927), .B2(new_n928), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n698), .A3(new_n926), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n933), .B1(new_n941), .B2(KEYINPUT42), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n605), .A2(G299), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n605), .A2(G299), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT41), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n613), .A2(new_n821), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n605), .A2(G299), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n949), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n616), .B(new_n852), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n954), .A2(KEYINPUT107), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT107), .B1(new_n955), .B2(new_n952), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n942), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n923), .B1(new_n960), .B2(new_n606), .ZN(G295));
  OAI21_X1  g536(.A(new_n923), .B1(new_n960), .B2(new_n606), .ZN(G331));
  AND2_X1   g537(.A1(G168), .A2(new_n852), .ZN(new_n963));
  NOR2_X1   g538(.A1(G168), .A2(new_n852), .ZN(new_n964));
  OAI21_X1  g539(.A(G171), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(G286), .A2(new_n846), .A3(new_n851), .ZN(new_n966));
  NAND2_X1  g541(.A1(G168), .A2(new_n852), .ZN(new_n967));
  NAND3_X1  g542(.A1(G301), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n965), .A2(new_n951), .A3(new_n953), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n952), .ZN(new_n970));
  AND3_X1   g545(.A1(G301), .A2(new_n966), .A3(new_n967), .ZN(new_n971));
  AOI21_X1  g546(.A(G301), .B1(new_n966), .B2(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n939), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n969), .A2(new_n973), .A3(new_n935), .A4(new_n938), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n945), .A2(new_n950), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n965), .A2(new_n980), .A3(new_n968), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n952), .B1(new_n965), .B2(new_n968), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT108), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT108), .B1(new_n936), .B2(new_n937), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n981), .A2(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n918), .A3(new_n977), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n979), .B1(KEYINPUT43), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n985), .A2(new_n977), .A3(new_n991), .A4(new_n918), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(KEYINPUT43), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n975), .A2(new_n994), .A3(new_n976), .A4(new_n977), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(KEYINPUT44), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n993), .A2(KEYINPUT111), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT111), .B1(new_n993), .B2(new_n996), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n989), .B1(new_n997), .B2(new_n998), .ZN(G397));
  INV_X1    g574(.A(new_n471), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n472), .A2(new_n473), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n463), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT112), .B(G40), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n491), .B2(new_n494), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(G1996), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n887), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT113), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n813), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n887), .A2(G1996), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n716), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n714), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n813), .A2(G2067), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1010), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n870), .B(new_n716), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT114), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1010), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n697), .A3(new_n698), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1018), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1011), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT46), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1015), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1025), .B1(new_n1032), .B2(new_n887), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(KEYINPUT46), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1022), .A2(new_n1029), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1005), .B1(new_n1008), .B2(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n1007), .C1(new_n491), .C2(new_n494), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  INV_X1    g618(.A(G2084), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n894), .A2(new_n1045), .A3(new_n1041), .A4(new_n1007), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n894), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1006), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1966), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1039), .B1(new_n1053), .B2(G286), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1047), .A2(new_n1052), .A3(G168), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1039), .B1(new_n1055), .B2(G8), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT62), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(KEYINPUT51), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1060), .B(new_n1061), .C1(new_n1056), .C2(new_n1054), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G303), .A2(G8), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT55), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1065), .A2(new_n1006), .A3(new_n1042), .ZN(new_n1066));
  INV_X1    g641(.A(G2090), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1066), .A2(new_n1067), .B1(new_n1050), .B2(new_n693), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(G305), .B(KEYINPUT49), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n581), .A2(KEYINPUT116), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G1981), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1008), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1069), .B1(new_n1006), .B2(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(G1981), .A3(new_n1072), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n686), .A2(G1976), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(G8), .C1(new_n1008), .C2(new_n1005), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1083));
  INV_X1    g658(.A(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1076), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1080), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1040), .A2(new_n1043), .A3(new_n1067), .A4(new_n1046), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1050), .A2(new_n693), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1064), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(G8), .A3(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1070), .A2(new_n1087), .A3(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1048), .A2(new_n1006), .A3(new_n1049), .A4(new_n801), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1043), .A2(new_n1065), .A3(new_n1006), .A4(new_n1046), .ZN(new_n1098));
  INV_X1    g673(.A(G1961), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1059), .A2(new_n1062), .A3(new_n1093), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1070), .A2(new_n1087), .A3(new_n1092), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1053), .A2(G8), .A3(G168), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1080), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1080), .A2(new_n1086), .A3(KEYINPUT117), .A4(new_n1083), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1069), .B(new_n1064), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1080), .A2(new_n1084), .A3(new_n686), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G305), .A2(G1981), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1116), .B(KEYINPUT118), .Z(new_n1117));
  OAI21_X1  g692(.A(new_n1076), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1108), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1091), .B1(new_n1090), .B2(G8), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1121), .A2(new_n1107), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT63), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1104), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1060), .B1(new_n1056), .B2(new_n1054), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n801), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n471), .A2(new_n474), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1048), .A2(new_n1049), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1048), .A2(KEYINPUT124), .A3(new_n1049), .A4(new_n1128), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1131), .A2(new_n1132), .B1(new_n1095), .B2(new_n1094), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1100), .A2(KEYINPUT123), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1098), .A2(new_n1135), .A3(new_n1099), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(G301), .A4(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1102), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1093), .B(new_n1126), .C1(new_n1138), .C2(KEYINPUT54), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1048), .A2(new_n1006), .A3(new_n1049), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1066), .B2(G1956), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  OAI21_X1  g718(.A(G299), .B1(KEYINPUT119), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(KEYINPUT119), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1146), .B(new_n1141), .C1(new_n1066), .C2(G1956), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1148), .A2(new_n1149), .A3(KEYINPUT122), .A4(KEYINPUT61), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1050), .B2(G1996), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n547), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1162), .A3(new_n547), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1155), .A2(new_n1156), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1006), .A2(new_n1075), .A3(new_n1014), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT120), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1098), .A2(new_n796), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1166), .A2(new_n605), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n605), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT60), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1154), .A2(new_n1164), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1169), .A2(new_n1149), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1174), .A2(new_n1148), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1139), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT125), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1133), .A2(new_n1134), .A3(new_n1179), .A4(new_n1136), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(G171), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1101), .A2(G171), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1181), .A2(KEYINPUT126), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT126), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1125), .B1(new_n1176), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n698), .B(G1986), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1018), .B(new_n1026), .C1(new_n1010), .C2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1038), .B1(new_n1188), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g766(.A(G227), .B1(new_n645), .B2(G14), .ZN(new_n1193));
  AND2_X1   g767(.A1(new_n921), .A2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g768(.A1(new_n1194), .A2(G319), .A3(new_n679), .A4(new_n987), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


