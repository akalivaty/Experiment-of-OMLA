//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n204), .A2(new_n205), .B1(KEYINPUT86), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OR3_X1    g008(.A1(new_n209), .A2(new_n206), .A3(KEYINPUT86), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n203), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n209), .B2(new_n206), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT15), .A3(new_n203), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n202), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g017(.A(KEYINPUT87), .B(KEYINPUT17), .C1(new_n212), .C2(new_n215), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT94), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT8), .ZN(new_n233));
  OR2_X1    g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT95), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT95), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n237), .B1(G99gat), .B2(G106gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n231), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(G99gat), .B(G106gat), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT96), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n233), .A2(KEYINPUT95), .A3(new_n234), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT95), .B1(new_n233), .B2(new_n234), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n242), .B1(new_n247), .B2(new_n231), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n235), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n224), .A2(new_n230), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n243), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n244), .B1(new_n252), .B2(KEYINPUT96), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n216), .A2(new_n217), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n220), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n253), .A2(new_n216), .B1(KEYINPUT41), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G134gat), .B(G162gat), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n261), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n257), .A2(KEYINPUT41), .ZN(new_n265));
  XNOR2_X1  g064(.A(G190gat), .B(G218gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n262), .A2(new_n267), .A3(new_n263), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273));
  INV_X1    g072(.A(G1gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT16), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G1gat), .B2(new_n273), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(G8gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(G8gat), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT88), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n279), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT88), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT92), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G57gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G64gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(G71gat), .A2(G78gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n290));
  NAND2_X1  g089(.A1(G71gat), .A2(G78gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G64gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT9), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(KEYINPUT91), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n289), .B1(new_n297), .B2(new_n291), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n297), .B2(new_n291), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n293), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n285), .B1(KEYINPUT21), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n300), .B(KEYINPUT21), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n285), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n305));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n304), .B(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G231gat), .A2(G233gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT93), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G155gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n312), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n272), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G176gat), .B(G204gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT98), .ZN(new_n318));
  XNOR2_X1  g117(.A(G120gat), .B(G148gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G230gat), .A2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT99), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT97), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n300), .B1(new_n251), .B2(new_n248), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n253), .B2(new_n300), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n327), .B2(KEYINPUT10), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n249), .A2(new_n243), .A3(new_n250), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n243), .B1(new_n249), .B2(new_n250), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT96), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT96), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n251), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n300), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(KEYINPUT97), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n253), .A2(KEYINPUT10), .A3(new_n301), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n324), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n336), .A2(new_n322), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n321), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n321), .ZN(new_n344));
  INV_X1    g143(.A(new_n340), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n328), .B2(new_n338), .ZN(new_n346));
  INV_X1    g145(.A(new_n322), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n316), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT90), .ZN(new_n352));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353));
  INV_X1    g152(.A(G85gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT0), .B(G57gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(KEYINPUT75), .B(KEYINPUT2), .Z(new_n362));
  XNOR2_X1  g161(.A(G141gat), .B(G148gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT76), .ZN(new_n365));
  INV_X1    g164(.A(new_n363), .ZN(new_n366));
  NOR3_X1   g165(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n359), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G113gat), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n372), .A2(G120gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(G120gat), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT1), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G127gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G134gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT68), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n381), .B2(new_n377), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n383), .B2(new_n382), .ZN(new_n385));
  INV_X1    g184(.A(new_n377), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n375), .A2(new_n386), .A3(new_n379), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n368), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n391), .A2(KEYINPUT4), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n389), .A2(new_n388), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(KEYINPUT77), .ZN(new_n395));
  OAI22_X1  g194(.A1(new_n392), .A2(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n394), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n393), .B2(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n391), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n389), .A2(new_n388), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n402), .B(KEYINPUT5), .C1(new_n397), .C2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n358), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G197gat), .B(G204gat), .Z(new_n407));
  AOI21_X1  g206(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT71), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n409), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT71), .B(new_n410), .C1(new_n407), .C2(new_n408), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G169gat), .A2(G176gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT66), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT24), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT67), .B(G190gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(G183gat), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(KEYINPUT25), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n424), .B1(G183gat), .B2(G190gat), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(KEYINPUT25), .ZN(new_n430));
  INV_X1    g229(.A(new_n425), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT27), .B(G183gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT28), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n417), .B(KEYINPUT26), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n421), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n423), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(G226gat), .A3(G233gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT72), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n430), .A2(new_n438), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(KEYINPUT29), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n440), .A2(KEYINPUT72), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n416), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n444), .A2(new_n440), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n415), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT73), .ZN(new_n453));
  XNOR2_X1  g252(.A(G8gat), .B(G36gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n453), .B(new_n454), .Z(new_n455));
  XOR2_X1   g254(.A(new_n455), .B(KEYINPUT74), .Z(new_n456));
  NOR2_X1   g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n455), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT30), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n459), .A2(KEYINPUT30), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n406), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n396), .A2(new_n398), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n404), .A2(new_n397), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(KEYINPUT39), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(new_n358), .C1(KEYINPUT39), .C2(new_n463), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n415), .B1(new_n371), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT3), .B1(new_n411), .B2(new_n471), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n472), .A2(new_n473), .B1(new_n369), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  INV_X1    g275(.A(G228gat), .ZN(new_n477));
  INV_X1    g276(.A(G233gat), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n472), .A2(new_n477), .A3(new_n478), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT3), .B1(new_n415), .B2(new_n471), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n369), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G22gat), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT82), .B1(new_n483), .B2(new_n484), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT80), .B(G50gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n487), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n485), .A2(KEYINPUT82), .A3(new_n486), .A4(new_n493), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n406), .A2(KEYINPUT6), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n399), .A2(new_n358), .A3(new_n405), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n406), .A2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT37), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n451), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n448), .B2(new_n416), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n415), .B1(new_n445), .B2(new_n446), .ZN(new_n505));
  AOI211_X1 g304(.A(KEYINPUT38), .B(new_n456), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n459), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n500), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT38), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n458), .B1(new_n451), .B2(new_n502), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n510), .A2(KEYINPUT83), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n510), .A2(KEYINPUT83), .B1(new_n502), .B2(new_n451), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n470), .B(new_n497), .C1(new_n508), .C2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G43gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(G71gat), .B(G99gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n443), .A2(KEYINPUT70), .A3(new_n385), .A4(new_n387), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n439), .B2(new_n388), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n439), .A2(new_n388), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G227gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT64), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT65), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT33), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n517), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(KEYINPUT32), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR3_X1    g329(.A1(new_n522), .A2(KEYINPUT34), .A3(new_n525), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT34), .B1(new_n522), .B2(new_n524), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n529), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n530), .B2(new_n535), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n540));
  INV_X1    g339(.A(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n536), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n514), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n460), .A2(new_n461), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n399), .A2(new_n405), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n357), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n550), .A2(KEYINPUT78), .A3(new_n551), .A4(new_n499), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n501), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT78), .B1(new_n498), .B2(new_n499), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n497), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n497), .A2(new_n539), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT35), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT35), .B1(new_n500), .B2(new_n501), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(new_n497), .A3(new_n548), .A4(new_n539), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n546), .A2(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n254), .A2(new_n282), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n219), .B2(new_n218), .ZN(new_n564));
  INV_X1    g363(.A(new_n284), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n282), .A2(new_n283), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n216), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n281), .A2(new_n284), .A3(new_n215), .A4(new_n212), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n568), .B(KEYINPUT13), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n569), .A2(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n567), .A2(new_n564), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(KEYINPUT18), .A3(new_n568), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n579));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G169gat), .B(G197gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n575), .A2(new_n577), .A3(new_n585), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT89), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n352), .B1(new_n562), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n559), .A2(new_n561), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n557), .A2(new_n514), .A3(new_n545), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT90), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n351), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n553), .A2(new_n554), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g399(.A1(new_n597), .A2(KEYINPUT100), .A3(new_n547), .ZN(new_n601));
  INV_X1    g400(.A(new_n351), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT90), .B1(new_n594), .B2(new_n595), .ZN(new_n603));
  AOI211_X1 g402(.A(new_n352), .B(new_n590), .C1(new_n592), .C2(new_n593), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n602), .B(new_n547), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT16), .B(G8gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n601), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT42), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n601), .A2(new_n607), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G8gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n608), .A2(new_n611), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n605), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n597), .A2(KEYINPUT101), .A3(new_n547), .A4(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(new_n614), .A3(new_n620), .ZN(G1325gat));
  AOI21_X1  g420(.A(G15gat), .B1(new_n597), .B2(new_n539), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n540), .A2(new_n544), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(G15gat), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n597), .B2(new_n624), .ZN(G1326gat));
  NAND2_X1  g424(.A1(new_n597), .A2(new_n556), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT43), .B(G22gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1327gat));
  AOI211_X1 g427(.A(KEYINPUT44), .B(new_n271), .C1(new_n592), .C2(new_n593), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n594), .A2(new_n272), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT44), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n349), .B(KEYINPUT103), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n588), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n585), .B1(new_n575), .B2(new_n577), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n315), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n313), .A2(KEYINPUT102), .A3(new_n314), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n635), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n598), .ZN(new_n645));
  OAI21_X1  g444(.A(G29gat), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n315), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n647), .A2(new_n271), .A3(new_n349), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n591), .B2(new_n596), .ZN(new_n650));
  INV_X1    g449(.A(G29gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n598), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n646), .B1(new_n653), .B2(new_n654), .ZN(G1328gat));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n548), .A2(G36gat), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n648), .B(new_n657), .C1(new_n603), .C2(new_n604), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G36gat), .B1(new_n644), .B2(new_n548), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(KEYINPUT46), .A3(new_n659), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(G43gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n667), .A3(new_n539), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n271), .B1(new_n592), .B2(new_n593), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n623), .B(new_n643), .C1(new_n671), .C2(new_n629), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G43gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n668), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n668), .B2(new_n673), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(G1330gat));
  OAI211_X1 g476(.A(new_n556), .B(new_n643), .C1(new_n671), .C2(new_n629), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G50gat), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT48), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(G50gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n650), .A2(new_n682), .A3(new_n556), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n679), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n683), .B(new_n679), .C1(new_n680), .C2(KEYINPUT48), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1331gat));
  NOR4_X1   g486(.A1(new_n634), .A2(new_n315), .A3(new_n272), .A4(new_n589), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n594), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n598), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g491(.A1(new_n689), .A2(new_n548), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  AND2_X1   g493(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n539), .A2(KEYINPUT108), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n542), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n689), .B2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n689), .A2(new_n698), .A3(new_n545), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n703), .B(new_n709), .C1(new_n706), .C2(new_n707), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1334gat));
  NAND2_X1  g512(.A1(new_n690), .A2(new_n556), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n647), .A2(new_n589), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n350), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n633), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G85gat), .B1(new_n719), .B2(new_n645), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n631), .B2(new_n717), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n669), .A2(KEYINPUT51), .A3(new_n716), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n724), .A2(new_n354), .A3(new_n598), .A4(new_n349), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n720), .A2(new_n725), .ZN(G1336gat));
  NOR2_X1   g525(.A1(new_n548), .A2(G92gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n635), .A3(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n547), .B(new_n718), .C1(new_n671), .C2(new_n629), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G92gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n730), .A3(KEYINPUT110), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT52), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n728), .A2(new_n730), .A3(KEYINPUT110), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1337gat));
  OAI21_X1  g534(.A(G99gat), .B1(new_n719), .B2(new_n545), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n542), .A2(G99gat), .A3(new_n350), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n724), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1338gat));
  NOR2_X1   g538(.A1(new_n497), .A2(G106gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n635), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(G106gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n718), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n630), .B2(new_n632), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(new_n556), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT53), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G106gat), .B1(new_n719), .B2(new_n497), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n749), .A3(new_n741), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(G1339gat));
  AND2_X1   g550(.A1(new_n640), .A2(new_n641), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT97), .B1(new_n336), .B2(new_n337), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n325), .B(KEYINPUT10), .C1(new_n334), .C2(new_n335), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n324), .B(new_n340), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n756), .B(KEYINPUT54), .C1(new_n346), .C2(new_n347), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n340), .B1(new_n754), .B2(new_n755), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n760), .A3(new_n323), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n321), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n753), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n757), .A2(KEYINPUT55), .A3(new_n321), .A4(new_n761), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(new_n348), .A3(new_n589), .A4(new_n764), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n576), .A2(new_n568), .B1(new_n572), .B2(new_n574), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n583), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n588), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n349), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n272), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n270), .A3(new_n269), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n764), .A2(new_n348), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n320), .B1(new_n341), .B2(new_n760), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT55), .B1(new_n774), .B2(new_n757), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n752), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n316), .A2(new_n350), .A3(new_n638), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(new_n645), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n558), .A2(new_n547), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G113gat), .B1(new_n784), .B2(new_n590), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n589), .A2(new_n372), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1340gat));
  OAI21_X1  g586(.A(G120gat), .B1(new_n784), .B2(new_n634), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n350), .A2(G120gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT112), .ZN(G1341gat));
  NOR3_X1   g590(.A1(new_n784), .A2(new_n376), .A3(new_n752), .ZN(new_n792));
  INV_X1    g591(.A(new_n784), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n647), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n792), .B1(new_n376), .B2(new_n794), .ZN(G1342gat));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n272), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G134gat), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT113), .Z(new_n798));
  NOR2_X1   g597(.A1(new_n796), .A2(G134gat), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT56), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1343gat));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n774), .A2(new_n757), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(KEYINPUT114), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(KEYINPUT114), .B2(new_n803), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n595), .A2(new_n348), .A3(new_n764), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n770), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n271), .ZN(new_n808));
  INV_X1    g607(.A(new_n776), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n647), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n779), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n556), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT57), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n780), .A2(new_n781), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n556), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n623), .A2(new_n645), .A3(new_n547), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G141gat), .B1(new_n818), .B2(new_n590), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n623), .A2(new_n547), .A3(new_n497), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n782), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(G141gat), .A3(new_n590), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(KEYINPUT58), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n818), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n589), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n826), .B2(G141gat), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(G1344gat));
  INV_X1    g628(.A(new_n821), .ZN(new_n830));
  INV_X1    g629(.A(G148gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n349), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n556), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n351), .A2(new_n595), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n815), .B(new_n556), .C1(new_n810), .C2(new_n835), .ZN(new_n836));
  AND4_X1   g635(.A1(new_n349), .A2(new_n834), .A3(new_n836), .A4(new_n817), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(new_n831), .ZN(new_n838));
  XNOR2_X1  g637(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT117), .B(new_n839), .C1(new_n837), .C2(new_n831), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n831), .A2(KEYINPUT59), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n818), .B2(new_n350), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n832), .B1(new_n840), .B2(new_n844), .ZN(G1345gat));
  AOI21_X1  g644(.A(KEYINPUT118), .B1(new_n830), .B2(new_n647), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(G155gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n830), .A2(KEYINPUT118), .A3(new_n647), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n642), .A2(G155gat), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n847), .A2(new_n848), .B1(new_n825), .B2(new_n849), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n818), .B2(new_n271), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n271), .A2(G162gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n821), .B2(new_n852), .ZN(G1347gat));
  NOR3_X1   g652(.A1(new_n780), .A2(new_n781), .A3(new_n598), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n558), .A2(new_n548), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(G169gat), .A3(new_n638), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT119), .Z(new_n858));
  AND4_X1   g657(.A1(new_n547), .A2(new_n497), .A3(new_n699), .A4(new_n701), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n814), .A2(KEYINPUT120), .A3(new_n645), .A4(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n773), .A2(new_n775), .A3(new_n638), .ZN(new_n861));
  INV_X1    g660(.A(new_n770), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n271), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n642), .B1(new_n863), .B2(new_n809), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT111), .B1(new_n864), .B2(new_n811), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(new_n645), .A3(new_n866), .A4(new_n859), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n590), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n858), .A2(new_n871), .ZN(G1348gat));
  NAND4_X1  g671(.A1(new_n860), .A2(new_n869), .A3(G176gat), .A4(new_n635), .ZN(new_n873));
  INV_X1    g672(.A(G176gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n856), .B2(new_n350), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n873), .A2(new_n875), .ZN(G1349gat));
  NAND2_X1  g675(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n647), .A2(new_n432), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n856), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n869), .A3(new_n642), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(G183gat), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n881), .B(new_n882), .ZN(G1350gat));
  NOR3_X1   g682(.A1(new_n856), .A2(new_n271), .A3(new_n425), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT122), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n860), .A2(new_n869), .A3(new_n272), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT123), .B1(new_n886), .B2(G190gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT124), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n886), .A2(G190gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n886), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n894), .A2(KEYINPUT124), .A3(new_n890), .A4(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT61), .B1(new_n887), .B2(new_n888), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n885), .B1(new_n891), .B2(new_n898), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n623), .A2(new_n598), .A3(new_n548), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n834), .A2(new_n836), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(G197gat), .A3(new_n595), .ZN(new_n902));
  INV_X1    g701(.A(G197gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n545), .A2(new_n547), .A3(new_n556), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT125), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n854), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n638), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT126), .ZN(G1352gat));
  INV_X1    g708(.A(G204gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n901), .B2(new_n635), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n350), .A2(G204gat), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OR3_X1    g712(.A1(new_n906), .A2(KEYINPUT62), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT62), .B1(new_n906), .B2(new_n913), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT127), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT127), .B1(new_n911), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1353gat));
  OR3_X1    g718(.A1(new_n906), .A2(G211gat), .A3(new_n315), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n647), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n271), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n272), .A3(new_n854), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n901), .A2(new_n926), .B1(new_n927), .B2(new_n925), .ZN(G1355gat));
endmodule


