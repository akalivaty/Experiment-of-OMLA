

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797;

  NOR2_X1 U368 ( .A1(n459), .A2(n464), .ZN(n578) );
  BUF_X1 U369 ( .A(n606), .Z(n345) );
  NAND2_X1 U370 ( .A1(n394), .A2(n393), .ZN(n682) );
  AND2_X1 U371 ( .A1(n399), .A2(n395), .ZN(n394) );
  NAND2_X1 U372 ( .A1(n469), .A2(n466), .ZN(n582) );
  XNOR2_X1 U373 ( .A(n628), .B(KEYINPUT6), .ZN(n606) );
  XNOR2_X1 U374 ( .A(n502), .B(KEYINPUT64), .ZN(n504) );
  INV_X2 U375 ( .A(G953), .ZN(n787) );
  XNOR2_X1 U376 ( .A(n505), .B(n545), .ZN(n426) );
  AND2_X2 U377 ( .A1(n405), .A2(n402), .ZN(n401) );
  NAND2_X1 U378 ( .A1(KEYINPUT82), .A2(n458), .ZN(n455) );
  AND2_X4 U379 ( .A1(n445), .A2(n443), .ZN(n372) );
  AND2_X2 U380 ( .A1(n452), .A2(n446), .ZN(n445) );
  NAND2_X2 U381 ( .A1(n404), .A2(n403), .ZN(n597) );
  XNOR2_X2 U382 ( .A(n582), .B(n556), .ZN(n575) );
  XNOR2_X2 U383 ( .A(n436), .B(n347), .ZN(n678) );
  XNOR2_X1 U384 ( .A(n578), .B(KEYINPUT35), .ZN(n687) );
  NOR2_X1 U385 ( .A1(n618), .A2(n641), .ZN(n715) );
  XNOR2_X1 U386 ( .A(n646), .B(n645), .ZN(n661) );
  XNOR2_X1 U387 ( .A(n656), .B(n378), .ZN(n746) );
  AND2_X1 U388 ( .A1(n588), .A2(n587), .ZN(n647) );
  AND2_X1 U389 ( .A1(n471), .A2(n470), .ZN(n469) );
  XNOR2_X1 U390 ( .A(KEYINPUT83), .B(KEYINPUT36), .ZN(n609) );
  NAND2_X1 U391 ( .A1(n611), .A2(n610), .ZN(n686) );
  XNOR2_X1 U392 ( .A(n433), .B(n609), .ZN(n611) );
  XNOR2_X2 U393 ( .A(n659), .B(KEYINPUT80), .ZN(n672) );
  INV_X1 U394 ( .A(n596), .ZN(n407) );
  XOR2_X1 U395 ( .A(G146), .B(G125), .Z(n498) );
  XNOR2_X1 U396 ( .A(n498), .B(n487), .ZN(n781) );
  INV_X1 U397 ( .A(n364), .ZN(n764) );
  XNOR2_X1 U398 ( .A(n682), .B(KEYINPUT78), .ZN(n636) );
  OR2_X1 U399 ( .A1(n715), .A2(KEYINPUT47), .ZN(n621) );
  INV_X1 U400 ( .A(KEYINPUT71), .ZN(n391) );
  NOR2_X1 U401 ( .A1(n724), .A2(n472), .ZN(n590) );
  AND2_X1 U402 ( .A1(n595), .A2(KEYINPUT44), .ZN(n453) );
  NOR2_X1 U403 ( .A1(n385), .A2(n384), .ZN(n382) );
  INV_X1 U404 ( .A(KEYINPUT38), .ZN(n378) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n560) );
  NAND2_X1 U406 ( .A1(n746), .A2(n747), .ZN(n752) );
  INV_X1 U407 ( .A(G469), .ZN(n467) );
  NAND2_X1 U408 ( .A1(G902), .A2(G469), .ZN(n470) );
  INV_X1 U409 ( .A(n697), .ZN(n468) );
  XNOR2_X1 U410 ( .A(n543), .B(n542), .ZN(n598) );
  XNOR2_X1 U411 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U412 ( .A(G101), .B(G113), .ZN(n511) );
  XNOR2_X1 U413 ( .A(KEYINPUT3), .B(G119), .ZN(n510) );
  XNOR2_X1 U414 ( .A(G140), .B(KEYINPUT92), .ZN(n532) );
  XNOR2_X1 U415 ( .A(G119), .B(G137), .ZN(n530) );
  XNOR2_X1 U416 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n478) );
  XNOR2_X1 U417 ( .A(n488), .B(KEYINPUT11), .ZN(n423) );
  INV_X1 U418 ( .A(KEYINPUT105), .ZN(n397) );
  NAND2_X1 U419 ( .A1(n398), .A2(n397), .ZN(n396) );
  XNOR2_X1 U420 ( .A(n777), .B(KEYINPUT124), .ZN(n368) );
  NOR2_X1 U421 ( .A1(n764), .A2(n439), .ZN(n438) );
  INV_X1 U422 ( .A(G475), .ZN(n439) );
  NOR2_X1 U423 ( .A1(n764), .A2(n440), .ZN(n371) );
  INV_X1 U424 ( .A(G210), .ZN(n440) );
  XNOR2_X1 U425 ( .A(n570), .B(n361), .ZN(n360) );
  NAND2_X1 U426 ( .A1(n380), .A2(n379), .ZN(n387) );
  NOR2_X1 U427 ( .A1(n412), .A2(n391), .ZN(n380) );
  XNOR2_X1 U428 ( .A(G902), .B(KEYINPUT15), .ZN(n667) );
  INV_X1 U429 ( .A(n665), .ZN(n449) );
  INV_X1 U430 ( .A(n670), .ZN(n451) );
  INV_X1 U431 ( .A(G237), .ZN(n513) );
  NAND2_X1 U432 ( .A1(n407), .A2(n406), .ZN(n400) );
  NOR2_X1 U433 ( .A1(n457), .A2(n595), .ZN(n406) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n488) );
  XNOR2_X1 U435 ( .A(G140), .B(G131), .ZN(n551) );
  NAND2_X1 U436 ( .A1(n450), .A2(n447), .ZN(n446) );
  NAND2_X1 U437 ( .A1(n448), .A2(n670), .ZN(n447) );
  NAND2_X1 U438 ( .A1(n451), .A2(KEYINPUT65), .ZN(n450) );
  NAND2_X1 U439 ( .A1(n449), .A2(KEYINPUT65), .ZN(n448) );
  XNOR2_X1 U440 ( .A(G146), .B(G125), .ZN(n499) );
  NAND2_X1 U441 ( .A1(G234), .A2(G237), .ZN(n520) );
  AND2_X1 U442 ( .A1(n604), .A2(n623), .ZN(n613) );
  XOR2_X1 U443 ( .A(KEYINPUT5), .B(KEYINPUT73), .Z(n562) );
  XOR2_X1 U444 ( .A(G122), .B(KEYINPUT9), .Z(n481) );
  XNOR2_X1 U445 ( .A(G101), .B(G104), .ZN(n547) );
  XNOR2_X1 U446 ( .A(G110), .B(G107), .ZN(n546) );
  NOR2_X1 U447 ( .A1(n752), .A2(n749), .ZN(n640) );
  NAND2_X1 U448 ( .A1(n745), .A2(n463), .ZN(n460) );
  NAND2_X1 U449 ( .A1(n468), .A2(n346), .ZN(n466) );
  INV_X2 U450 ( .A(n598), .ZN(n734) );
  NOR2_X1 U451 ( .A1(n764), .A2(n568), .ZN(n437) );
  XNOR2_X1 U452 ( .A(n414), .B(n537), .ZN(n689) );
  XNOR2_X1 U453 ( .A(n538), .B(n781), .ZN(n414) );
  XNOR2_X1 U454 ( .A(n413), .B(n535), .ZN(n538) );
  AND2_X2 U455 ( .A1(n372), .A2(n364), .ZN(n688) );
  XNOR2_X1 U456 ( .A(n377), .B(KEYINPUT42), .ZN(n797) );
  NOR2_X1 U457 ( .A1(n767), .A2(n641), .ZN(n377) );
  AND2_X1 U458 ( .A1(n661), .A2(n723), .ZN(n683) );
  NAND2_X1 U459 ( .A1(n643), .A2(n397), .ZN(n393) );
  AND2_X1 U460 ( .A1(n396), .A2(n351), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n367), .B(n366), .ZN(G69) );
  XNOR2_X1 U462 ( .A(n780), .B(KEYINPUT125), .ZN(n366) );
  NAND2_X1 U463 ( .A1(n368), .A2(n359), .ZN(n367) );
  INV_X1 U464 ( .A(KEYINPUT60), .ZN(n416) );
  INV_X1 U465 ( .A(KEYINPUT56), .ZN(n408) );
  INV_X1 U466 ( .A(n360), .ZN(n796) );
  AND2_X1 U467 ( .A1(n555), .A2(n467), .ZN(n346) );
  XOR2_X1 U468 ( .A(n567), .B(n566), .Z(n347) );
  XOR2_X1 U469 ( .A(G113), .B(G143), .Z(n348) );
  AND2_X1 U470 ( .A1(G214), .A2(n560), .ZN(n349) );
  XNOR2_X1 U471 ( .A(n529), .B(KEYINPUT22), .ZN(n591) );
  XOR2_X1 U472 ( .A(n650), .B(KEYINPUT46), .Z(n350) );
  AND2_X1 U473 ( .A1(n734), .A2(n733), .ZN(n730) );
  AND2_X1 U474 ( .A1(n588), .A2(n586), .ZN(n351) );
  AND2_X1 U475 ( .A1(n461), .A2(n351), .ZN(n352) );
  INV_X1 U476 ( .A(G902), .ZN(n555) );
  AND2_X1 U477 ( .A1(n656), .A2(KEYINPUT105), .ZN(n353) );
  INV_X1 U478 ( .A(n656), .ZN(n398) );
  INV_X1 U479 ( .A(KEYINPUT34), .ZN(n465) );
  XOR2_X1 U480 ( .A(n704), .B(n703), .Z(n354) );
  XOR2_X1 U481 ( .A(n696), .B(KEYINPUT59), .Z(n355) );
  XOR2_X1 U482 ( .A(n678), .B(n677), .Z(n356) );
  AND2_X1 U483 ( .A1(n670), .A2(KEYINPUT65), .ZN(n357) );
  AND2_X1 U484 ( .A1(n665), .A2(n671), .ZN(n358) );
  INV_X1 U485 ( .A(KEYINPUT44), .ZN(n458) );
  NOR2_X1 U486 ( .A1(n787), .A2(G952), .ZN(n705) );
  INV_X1 U487 ( .A(n705), .ZN(n410) );
  XOR2_X1 U488 ( .A(KEYINPUT123), .B(n776), .Z(n359) );
  OR2_X2 U489 ( .A1(n784), .A2(G146), .ZN(n558) );
  AND2_X1 U490 ( .A1(n585), .A2(n465), .ZN(n463) );
  NAND2_X1 U491 ( .A1(n462), .A2(KEYINPUT34), .ZN(n461) );
  NAND2_X1 U492 ( .A1(n719), .A2(n613), .ZN(n421) );
  XOR2_X1 U493 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n361) );
  NAND2_X1 U494 ( .A1(n432), .A2(n455), .ZN(n431) );
  INV_X1 U495 ( .A(n684), .ZN(n411) );
  NAND2_X1 U496 ( .A1(n369), .A2(n410), .ZN(n409) );
  XNOR2_X1 U497 ( .A(n370), .B(n354), .ZN(n369) );
  NAND2_X1 U498 ( .A1(n365), .A2(n786), .ZN(n362) );
  NOR2_X1 U499 ( .A1(n591), .A2(n734), .ZN(n363) );
  NAND2_X1 U500 ( .A1(n365), .A2(n786), .ZN(n728) );
  NOR2_X1 U501 ( .A1(n591), .A2(n734), .ZN(n572) );
  NAND2_X1 U502 ( .A1(n365), .A2(n787), .ZN(n777) );
  NAND2_X1 U503 ( .A1(n729), .A2(n365), .ZN(n364) );
  XNOR2_X2 U504 ( .A(n597), .B(KEYINPUT45), .ZN(n365) );
  NAND2_X1 U505 ( .A1(n372), .A2(n371), .ZN(n370) );
  NAND2_X1 U506 ( .A1(n372), .A2(n437), .ZN(n679) );
  NAND2_X1 U507 ( .A1(n372), .A2(n438), .ZN(n419) );
  NAND2_X1 U508 ( .A1(n688), .A2(G478), .ZN(n694) );
  NAND2_X1 U509 ( .A1(n444), .A2(n357), .ZN(n443) );
  NAND2_X1 U510 ( .A1(n457), .A2(KEYINPUT82), .ZN(n456) );
  XNOR2_X2 U511 ( .A(n581), .B(KEYINPUT31), .ZN(n724) );
  NAND2_X1 U512 ( .A1(n373), .A2(n658), .ZN(n659) );
  NAND2_X1 U513 ( .A1(n374), .A2(n381), .ZN(n373) );
  NAND2_X1 U514 ( .A1(n375), .A2(n392), .ZN(n374) );
  NAND2_X1 U515 ( .A1(n350), .A2(n383), .ZN(n375) );
  NAND2_X1 U516 ( .A1(n376), .A2(n411), .ZN(n650) );
  INV_X1 U517 ( .A(n797), .ZN(n376) );
  INV_X1 U518 ( .A(n746), .ZN(n642) );
  XNOR2_X2 U519 ( .A(n545), .B(n544), .ZN(n784) );
  XNOR2_X2 U520 ( .A(n504), .B(n503), .ZN(n545) );
  NAND2_X1 U521 ( .A1(n387), .A2(n651), .ZN(n384) );
  INV_X1 U522 ( .A(n638), .ZN(n379) );
  NAND2_X1 U523 ( .A1(n382), .A2(n350), .ZN(n381) );
  INV_X1 U524 ( .A(n386), .ZN(n383) );
  INV_X1 U525 ( .A(n388), .ZN(n385) );
  NAND2_X1 U526 ( .A1(n388), .A2(n387), .ZN(n386) );
  AND2_X2 U527 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U528 ( .A1(n412), .A2(n391), .ZN(n389) );
  NAND2_X1 U529 ( .A1(n638), .A2(n391), .ZN(n390) );
  INV_X1 U530 ( .A(n651), .ZN(n392) );
  NAND2_X1 U531 ( .A1(n634), .A2(n353), .ZN(n399) );
  NAND2_X1 U532 ( .A1(n456), .A2(n454), .ZN(n402) );
  NAND2_X1 U533 ( .A1(n401), .A2(n400), .ZN(n404) );
  NAND2_X1 U534 ( .A1(n407), .A2(n458), .ZN(n403) );
  NAND2_X1 U535 ( .A1(n596), .A2(n453), .ZN(n405) );
  XNOR2_X1 U536 ( .A(n409), .B(n408), .ZN(G51) );
  NOR2_X2 U537 ( .A1(n421), .A2(n607), .ZN(n653) );
  NAND2_X1 U538 ( .A1(n633), .A2(n747), .ZN(n415) );
  NAND2_X1 U539 ( .A1(n574), .A2(n528), .ZN(n529) );
  XNOR2_X2 U540 ( .A(n527), .B(KEYINPUT0), .ZN(n574) );
  NAND2_X1 U541 ( .A1(n622), .A2(n686), .ZN(n412) );
  INV_X1 U542 ( .A(n534), .ZN(n413) );
  XNOR2_X2 U543 ( .A(n608), .B(KEYINPUT19), .ZN(n612) );
  XNOR2_X2 U544 ( .A(n415), .B(n519), .ZN(n608) );
  XNOR2_X2 U545 ( .A(n517), .B(n516), .ZN(n633) );
  XNOR2_X1 U546 ( .A(n417), .B(n416), .ZN(G60) );
  NAND2_X1 U547 ( .A1(n418), .A2(n410), .ZN(n417) );
  XNOR2_X1 U548 ( .A(n419), .B(n355), .ZN(n418) );
  NAND2_X1 U549 ( .A1(n420), .A2(n608), .ZN(n433) );
  XNOR2_X1 U550 ( .A(n653), .B(n434), .ZN(n420) );
  XNOR2_X1 U551 ( .A(n424), .B(n422), .ZN(n696) );
  XNOR2_X1 U552 ( .A(n489), .B(n423), .ZN(n422) );
  XNOR2_X1 U553 ( .A(n781), .B(n425), .ZN(n424) );
  XNOR2_X1 U554 ( .A(n507), .B(n349), .ZN(n425) );
  OR2_X1 U555 ( .A1(n594), .A2(n706), .ZN(n457) );
  XNOR2_X1 U556 ( .A(n426), .B(n779), .ZN(n704) );
  XNOR2_X1 U557 ( .A(n512), .B(n566), .ZN(n779) );
  INV_X1 U558 ( .A(n428), .ZN(n430) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n428) );
  NAND2_X1 U560 ( .A1(n429), .A2(n427), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n428), .A2(n499), .ZN(n427) );
  NAND2_X1 U562 ( .A1(n430), .A2(n498), .ZN(n429) );
  OR2_X1 U563 ( .A1(n431), .A2(n594), .ZN(n454) );
  INV_X1 U564 ( .A(n706), .ZN(n432) );
  INV_X1 U565 ( .A(KEYINPUT109), .ZN(n434) );
  XNOR2_X2 U566 ( .A(n435), .B(G472), .ZN(n628) );
  NOR2_X2 U567 ( .A1(n678), .A2(G902), .ZN(n435) );
  NAND2_X1 U568 ( .A1(n558), .A2(n559), .ZN(n436) );
  INV_X1 U569 ( .A(n575), .ZN(n610) );
  XNOR2_X1 U570 ( .A(n580), .B(KEYINPUT100), .ZN(n576) );
  XNOR2_X2 U571 ( .A(n441), .B(KEYINPUT72), .ZN(n580) );
  NOR2_X2 U572 ( .A1(n575), .A2(n442), .ZN(n441) );
  INV_X1 U573 ( .A(n730), .ZN(n442) );
  INV_X1 U574 ( .A(n362), .ZN(n444) );
  NAND2_X1 U575 ( .A1(n728), .A2(n358), .ZN(n452) );
  NAND2_X1 U576 ( .A1(n352), .A2(n460), .ZN(n459) );
  XNOR2_X2 U577 ( .A(n577), .B(KEYINPUT33), .ZN(n745) );
  INV_X1 U578 ( .A(n585), .ZN(n462) );
  NOR2_X1 U579 ( .A1(n745), .A2(n465), .ZN(n464) );
  NAND2_X1 U580 ( .A1(n468), .A2(n555), .ZN(n624) );
  NAND2_X1 U581 ( .A1(n697), .A2(G469), .ZN(n471) );
  XNOR2_X2 U582 ( .A(n554), .B(n553), .ZN(n697) );
  AND2_X1 U583 ( .A1(n585), .A2(n584), .ZN(n472) );
  XOR2_X1 U584 ( .A(n629), .B(KEYINPUT103), .Z(n473) );
  NOR2_X1 U585 ( .A1(n360), .A2(n795), .ZN(n579) );
  INV_X1 U586 ( .A(KEYINPUT82), .ZN(n595) );
  INV_X1 U587 ( .A(KEYINPUT65), .ZN(n671) );
  INV_X1 U588 ( .A(KEYINPUT84), .ZN(n519) );
  XOR2_X1 U589 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n475) );
  NAND2_X1 U590 ( .A1(G234), .A2(n667), .ZN(n474) );
  XNOR2_X1 U591 ( .A(n475), .B(n474), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n539), .A2(G221), .ZN(n477) );
  INV_X1 U593 ( .A(KEYINPUT21), .ZN(n476) );
  XNOR2_X1 U594 ( .A(n477), .B(n476), .ZN(n733) );
  INV_X1 U595 ( .A(n733), .ZN(n493) );
  NAND2_X1 U596 ( .A1(n787), .A2(G234), .ZN(n479) );
  XNOR2_X1 U597 ( .A(n479), .B(n478), .ZN(n536) );
  NAND2_X1 U598 ( .A1(G217), .A2(n536), .ZN(n480) );
  XNOR2_X1 U599 ( .A(n481), .B(n480), .ZN(n485) );
  XOR2_X2 U600 ( .A(G116), .B(G107), .Z(n506) );
  XOR2_X1 U601 ( .A(KEYINPUT7), .B(n506), .Z(n483) );
  XNOR2_X1 U602 ( .A(G143), .B(G128), .ZN(n503) );
  XNOR2_X1 U603 ( .A(n503), .B(G134), .ZN(n482) );
  XNOR2_X1 U604 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U605 ( .A(n485), .B(n484), .ZN(n692) );
  NAND2_X1 U606 ( .A1(n692), .A2(n555), .ZN(n486) );
  XNOR2_X1 U607 ( .A(n486), .B(G478), .ZN(n586) );
  INV_X1 U608 ( .A(KEYINPUT10), .ZN(n487) );
  XOR2_X1 U609 ( .A(G122), .B(G104), .Z(n507) );
  XNOR2_X1 U610 ( .A(n551), .B(n348), .ZN(n489) );
  NAND2_X1 U611 ( .A1(n696), .A2(n555), .ZN(n491) );
  XOR2_X1 U612 ( .A(KEYINPUT13), .B(G475), .Z(n490) );
  XNOR2_X1 U613 ( .A(n491), .B(n490), .ZN(n588) );
  NOR2_X1 U614 ( .A1(n586), .A2(n588), .ZN(n492) );
  XNOR2_X1 U615 ( .A(n492), .B(KEYINPUT97), .ZN(n749) );
  NOR2_X1 U616 ( .A1(n493), .A2(n749), .ZN(n494) );
  XNOR2_X1 U617 ( .A(KEYINPUT98), .B(n494), .ZN(n528) );
  XNOR2_X2 U618 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n495) );
  INV_X1 U619 ( .A(n495), .ZN(n497) );
  XNOR2_X1 U620 ( .A(KEYINPUT85), .B(KEYINPUT74), .ZN(n496) );
  NAND2_X1 U621 ( .A1(G224), .A2(n787), .ZN(n500) );
  XNOR2_X1 U622 ( .A(n501), .B(n500), .ZN(n505) );
  XNOR2_X2 U623 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n502) );
  XOR2_X1 U624 ( .A(KEYINPUT16), .B(n506), .Z(n509) );
  XNOR2_X1 U625 ( .A(G110), .B(n507), .ZN(n508) );
  XNOR2_X1 U626 ( .A(n509), .B(n508), .ZN(n512) );
  XNOR2_X1 U627 ( .A(n511), .B(n510), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n704), .A2(n667), .ZN(n517) );
  NAND2_X1 U629 ( .A1(n555), .A2(n513), .ZN(n518) );
  NAND2_X1 U630 ( .A1(n518), .A2(G210), .ZN(n515) );
  INV_X1 U631 ( .A(KEYINPUT86), .ZN(n514) );
  XNOR2_X1 U632 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U633 ( .A1(n518), .A2(G214), .ZN(n747) );
  XNOR2_X1 U634 ( .A(n520), .B(KEYINPUT14), .ZN(n522) );
  NAND2_X1 U635 ( .A1(G952), .A2(n522), .ZN(n760) );
  NOR2_X1 U636 ( .A1(n760), .A2(G953), .ZN(n601) );
  NOR2_X1 U637 ( .A1(G898), .A2(n787), .ZN(n521) );
  XNOR2_X1 U638 ( .A(KEYINPUT87), .B(n521), .ZN(n778) );
  NAND2_X1 U639 ( .A1(n522), .A2(G902), .ZN(n523) );
  XNOR2_X1 U640 ( .A(n523), .B(KEYINPUT88), .ZN(n599) );
  NOR2_X1 U641 ( .A1(n778), .A2(n599), .ZN(n524) );
  NOR2_X1 U642 ( .A1(n601), .A2(n524), .ZN(n525) );
  XOR2_X1 U643 ( .A(KEYINPUT89), .B(n525), .Z(n526) );
  NOR2_X2 U644 ( .A1(n612), .A2(n526), .ZN(n527) );
  XOR2_X1 U645 ( .A(G110), .B(G128), .Z(n531) );
  XNOR2_X1 U646 ( .A(n531), .B(n530), .ZN(n535) );
  XOR2_X1 U647 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n533) );
  XNOR2_X1 U648 ( .A(n533), .B(n532), .ZN(n534) );
  AND2_X1 U649 ( .A1(G221), .A2(n536), .ZN(n537) );
  NOR2_X1 U650 ( .A1(n689), .A2(G902), .ZN(n543) );
  NAND2_X1 U651 ( .A1(G217), .A2(n539), .ZN(n541) );
  XOR2_X1 U652 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n540) );
  XNOR2_X1 U653 ( .A(G137), .B(G134), .ZN(n544) );
  NAND2_X1 U654 ( .A1(n784), .A2(G146), .ZN(n559) );
  NAND2_X1 U655 ( .A1(n558), .A2(n559), .ZN(n554) );
  XNOR2_X1 U656 ( .A(n547), .B(n546), .ZN(n550) );
  NAND2_X1 U657 ( .A1(n787), .A2(G227), .ZN(n548) );
  XNOR2_X1 U658 ( .A(n548), .B(KEYINPUT91), .ZN(n549) );
  XNOR2_X1 U659 ( .A(n550), .B(n549), .ZN(n552) );
  XNOR2_X1 U660 ( .A(n551), .B(KEYINPUT90), .ZN(n782) );
  XNOR2_X1 U661 ( .A(n552), .B(n782), .ZN(n553) );
  XNOR2_X1 U662 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n556) );
  BUF_X1 U663 ( .A(n575), .Z(n557) );
  NAND2_X1 U664 ( .A1(n560), .A2(G210), .ZN(n561) );
  XNOR2_X1 U665 ( .A(n562), .B(n561), .ZN(n565) );
  XNOR2_X1 U666 ( .A(G131), .B(KEYINPUT95), .ZN(n563) );
  XNOR2_X1 U667 ( .A(n563), .B(G116), .ZN(n564) );
  XNOR2_X1 U668 ( .A(n565), .B(n564), .ZN(n567) );
  INV_X1 U669 ( .A(G472), .ZN(n568) );
  NOR2_X1 U670 ( .A1(n557), .A2(n345), .ZN(n569) );
  NAND2_X1 U671 ( .A1(n572), .A2(n569), .ZN(n570) );
  AND2_X1 U672 ( .A1(n628), .A2(n557), .ZN(n571) );
  NAND2_X1 U673 ( .A1(n363), .A2(n571), .ZN(n573) );
  XNOR2_X1 U674 ( .A(n573), .B(KEYINPUT99), .ZN(n795) );
  BUF_X2 U675 ( .A(n574), .Z(n585) );
  NAND2_X1 U676 ( .A1(n576), .A2(n345), .ZN(n577) );
  NAND2_X1 U677 ( .A1(n579), .A2(n687), .ZN(n596) );
  INV_X1 U678 ( .A(n628), .ZN(n736) );
  AND2_X1 U679 ( .A1(n580), .A2(n736), .ZN(n741) );
  NAND2_X1 U680 ( .A1(n585), .A2(n741), .ZN(n581) );
  NAND2_X1 U681 ( .A1(n730), .A2(n582), .ZN(n583) );
  NOR2_X1 U682 ( .A1(n583), .A2(n736), .ZN(n584) );
  INV_X1 U683 ( .A(n586), .ZN(n587) );
  INV_X1 U684 ( .A(n647), .ZN(n589) );
  OR2_X1 U685 ( .A1(n588), .A2(n587), .ZN(n660) );
  AND2_X1 U686 ( .A1(n589), .A2(n660), .ZN(n751) );
  NOR2_X1 U687 ( .A1(n590), .A2(n751), .ZN(n594) );
  NAND2_X1 U688 ( .A1(n557), .A2(n734), .ZN(n592) );
  OR2_X1 U689 ( .A1(n592), .A2(n345), .ZN(n593) );
  NOR2_X1 U690 ( .A1(n591), .A2(n593), .ZN(n706) );
  AND2_X1 U691 ( .A1(n598), .A2(n733), .ZN(n604) );
  OR2_X1 U692 ( .A1(n599), .A2(n787), .ZN(n600) );
  OR2_X1 U693 ( .A1(n600), .A2(G900), .ZN(n603) );
  INV_X1 U694 ( .A(n601), .ZN(n602) );
  NAND2_X1 U695 ( .A1(n603), .A2(n602), .ZN(n623) );
  INV_X1 U696 ( .A(KEYINPUT101), .ZN(n605) );
  XNOR2_X2 U697 ( .A(n605), .B(n647), .ZN(n719) );
  INV_X1 U698 ( .A(n606), .ZN(n607) );
  BUF_X1 U699 ( .A(n612), .Z(n618) );
  INV_X1 U700 ( .A(n613), .ZN(n614) );
  OR2_X1 U701 ( .A1(n628), .A2(n614), .ZN(n616) );
  XOR2_X1 U702 ( .A(KEYINPUT106), .B(KEYINPUT28), .Z(n615) );
  XNOR2_X1 U703 ( .A(n616), .B(n615), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n617), .A2(n582), .ZN(n641) );
  OR2_X1 U705 ( .A1(n751), .A2(KEYINPUT47), .ZN(n619) );
  NAND2_X1 U706 ( .A1(n715), .A2(n619), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n730), .A2(n623), .ZN(n626) );
  XOR2_X1 U709 ( .A(n624), .B(G469), .Z(n625) );
  NOR2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n632) );
  INV_X1 U711 ( .A(n747), .ZN(n627) );
  NOR2_X2 U712 ( .A1(n628), .A2(n627), .ZN(n630) );
  XNOR2_X1 U713 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n629) );
  XNOR2_X1 U714 ( .A(n630), .B(n473), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n643) );
  INV_X1 U716 ( .A(n643), .ZN(n634) );
  BUF_X2 U717 ( .A(n633), .Z(n656) );
  NAND2_X1 U718 ( .A1(n751), .A2(KEYINPUT47), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n637), .B(KEYINPUT76), .ZN(n638) );
  XNOR2_X1 U721 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n639) );
  XNOR2_X1 U722 ( .A(n640), .B(n639), .ZN(n767) );
  OR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n646) );
  INV_X1 U724 ( .A(KEYINPUT81), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n644), .B(KEYINPUT39), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n661), .A2(n647), .ZN(n649) );
  XNOR2_X1 U727 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n649), .B(n648), .ZN(n684) );
  XNOR2_X1 U729 ( .A(KEYINPUT70), .B(KEYINPUT48), .ZN(n651) );
  AND2_X1 U730 ( .A1(n557), .A2(n747), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U732 ( .A(KEYINPUT102), .B(KEYINPUT43), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n657) );
  AND2_X1 U734 ( .A1(n657), .A2(n398), .ZN(n727) );
  INV_X1 U735 ( .A(n727), .ZN(n658) );
  INV_X1 U736 ( .A(n660), .ZN(n723) );
  NOR2_X2 U737 ( .A1(n672), .A2(n683), .ZN(n786) );
  INV_X1 U738 ( .A(KEYINPUT79), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n662), .A2(KEYINPUT2), .ZN(n664) );
  AND2_X1 U740 ( .A1(KEYINPUT2), .A2(KEYINPUT79), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n667), .A2(n663), .ZN(n666) );
  AND2_X1 U742 ( .A1(n664), .A2(n666), .ZN(n665) );
  INV_X1 U743 ( .A(n666), .ZN(n669) );
  INV_X1 U744 ( .A(n667), .ZN(n668) );
  OR2_X1 U745 ( .A1(n669), .A2(n668), .ZN(n670) );
  INV_X1 U746 ( .A(n672), .ZN(n676) );
  INV_X1 U747 ( .A(n683), .ZN(n673) );
  NAND2_X1 U748 ( .A1(n673), .A2(KEYINPUT2), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n674), .B(KEYINPUT75), .ZN(n675) );
  AND2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n729) );
  XNOR2_X1 U751 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n677) );
  XNOR2_X1 U752 ( .A(n679), .B(n356), .ZN(n680) );
  NAND2_X1 U753 ( .A1(n680), .A2(n410), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n681), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U755 ( .A(n682), .B(G143), .ZN(G45) );
  XOR2_X1 U756 ( .A(G134), .B(n683), .Z(G36) );
  XOR2_X1 U757 ( .A(G131), .B(n684), .Z(G33) );
  XOR2_X1 U758 ( .A(G125), .B(KEYINPUT37), .Z(n685) );
  XNOR2_X1 U759 ( .A(n686), .B(n685), .ZN(G27) );
  XNOR2_X1 U760 ( .A(n687), .B(G122), .ZN(G24) );
  NAND2_X1 U761 ( .A1(n688), .A2(G217), .ZN(n690) );
  XNOR2_X1 U762 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n691), .A2(n705), .ZN(G66) );
  XOR2_X1 U764 ( .A(n692), .B(KEYINPUT122), .Z(n693) );
  XNOR2_X1 U765 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U766 ( .A1(n695), .A2(n705), .ZN(G63) );
  NAND2_X1 U767 ( .A1(n688), .A2(G469), .ZN(n700) );
  XOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n698) );
  XNOR2_X1 U769 ( .A(n697), .B(n698), .ZN(n699) );
  XNOR2_X1 U770 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U771 ( .A1(n701), .A2(n705), .ZN(G54) );
  XOR2_X1 U772 ( .A(KEYINPUT77), .B(KEYINPUT54), .Z(n702) );
  XNOR2_X1 U773 ( .A(n702), .B(KEYINPUT55), .ZN(n703) );
  XOR2_X1 U774 ( .A(G101), .B(n706), .Z(G3) );
  NAND2_X1 U775 ( .A1(n719), .A2(n472), .ZN(n707) );
  XNOR2_X1 U776 ( .A(n707), .B(G104), .ZN(G6) );
  XOR2_X1 U777 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n709) );
  XNOR2_X1 U778 ( .A(G107), .B(KEYINPUT26), .ZN(n708) );
  XNOR2_X1 U779 ( .A(n709), .B(n708), .ZN(n710) );
  XOR2_X1 U780 ( .A(KEYINPUT111), .B(n710), .Z(n712) );
  NAND2_X1 U781 ( .A1(n472), .A2(n723), .ZN(n711) );
  XNOR2_X1 U782 ( .A(n712), .B(n711), .ZN(G9) );
  XOR2_X1 U783 ( .A(G128), .B(KEYINPUT29), .Z(n714) );
  NAND2_X1 U784 ( .A1(n715), .A2(n723), .ZN(n713) );
  XNOR2_X1 U785 ( .A(n714), .B(n713), .ZN(G30) );
  XOR2_X1 U786 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n717) );
  NAND2_X1 U787 ( .A1(n715), .A2(n719), .ZN(n716) );
  XNOR2_X1 U788 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U789 ( .A(G146), .B(n718), .ZN(G48) );
  XOR2_X1 U790 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n721) );
  NAND2_X1 U791 ( .A1(n719), .A2(n724), .ZN(n720) );
  XNOR2_X1 U792 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U793 ( .A(G113), .B(n722), .ZN(G15) );
  XOR2_X1 U794 ( .A(G116), .B(KEYINPUT117), .Z(n726) );
  NAND2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U796 ( .A(n726), .B(n725), .ZN(G18) );
  XOR2_X1 U797 ( .A(G140), .B(n727), .Z(G42) );
  NOR2_X1 U798 ( .A1(n362), .A2(n729), .ZN(n762) );
  NAND2_X1 U799 ( .A1(n557), .A2(n442), .ZN(n731) );
  XNOR2_X1 U800 ( .A(n731), .B(KEYINPUT119), .ZN(n732) );
  XNOR2_X1 U801 ( .A(KEYINPUT50), .B(n732), .ZN(n740) );
  NOR2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U803 ( .A(KEYINPUT49), .B(n735), .Z(n737) );
  NOR2_X1 U804 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U805 ( .A(n738), .B(KEYINPUT118), .Z(n739) );
  NOR2_X1 U806 ( .A1(n740), .A2(n739), .ZN(n742) );
  NOR2_X1 U807 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U808 ( .A(KEYINPUT51), .B(n743), .Z(n744) );
  NOR2_X1 U809 ( .A1(n767), .A2(n744), .ZN(n757) );
  NOR2_X1 U810 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U811 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U812 ( .A(n750), .B(KEYINPUT120), .ZN(n754) );
  NOR2_X1 U813 ( .A1(n752), .A2(n751), .ZN(n753) );
  OR2_X1 U814 ( .A1(n754), .A2(n753), .ZN(n755) );
  AND2_X1 U815 ( .A1(n745), .A2(n755), .ZN(n756) );
  NOR2_X1 U816 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U817 ( .A(n758), .B(KEYINPUT52), .ZN(n759) );
  NOR2_X1 U818 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U819 ( .A1(n762), .A2(n761), .ZN(n766) );
  INV_X1 U820 ( .A(KEYINPUT2), .ZN(n763) );
  OR2_X1 U821 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U822 ( .A1(n766), .A2(n765), .ZN(n772) );
  INV_X1 U823 ( .A(n767), .ZN(n768) );
  NAND2_X1 U824 ( .A1(n745), .A2(n768), .ZN(n769) );
  XOR2_X1 U825 ( .A(KEYINPUT121), .B(n769), .Z(n770) );
  NAND2_X1 U826 ( .A1(n787), .A2(n770), .ZN(n771) );
  NOR2_X1 U827 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U828 ( .A(n773), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U829 ( .A1(G953), .A2(G224), .ZN(n774) );
  XNOR2_X1 U830 ( .A(KEYINPUT61), .B(n774), .ZN(n775) );
  NAND2_X1 U831 ( .A1(n775), .A2(G898), .ZN(n776) );
  NAND2_X1 U832 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U833 ( .A(KEYINPUT126), .B(n781), .Z(n783) );
  XNOR2_X1 U834 ( .A(n783), .B(n782), .ZN(n785) );
  XOR2_X1 U835 ( .A(n784), .B(n785), .Z(n789) );
  XNOR2_X1 U836 ( .A(n786), .B(n789), .ZN(n788) );
  NAND2_X1 U837 ( .A1(n788), .A2(n787), .ZN(n794) );
  XOR2_X1 U838 ( .A(n789), .B(G227), .Z(n790) );
  NAND2_X1 U839 ( .A1(n790), .A2(G900), .ZN(n791) );
  NAND2_X1 U840 ( .A1(n791), .A2(G953), .ZN(n792) );
  XOR2_X1 U841 ( .A(KEYINPUT127), .B(n792), .Z(n793) );
  NAND2_X1 U842 ( .A1(n794), .A2(n793), .ZN(G72) );
  XOR2_X1 U843 ( .A(n795), .B(G110), .Z(G12) );
  XNOR2_X1 U844 ( .A(n796), .B(G119), .ZN(G21) );
  XOR2_X1 U845 ( .A(G137), .B(n797), .Z(G39) );
endmodule

