//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND3_X1  g0042(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(new_n215), .ZN(new_n244));
  NAND2_X1  g0044(.A1(KEYINPUT65), .A2(G58), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT8), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n207), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g0049(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n244), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G50), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n244), .B1(new_n206), .B2(G20), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G50), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G222), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n264), .B1(new_n265), .B2(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n272), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n273), .B1(G226), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n270), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n270), .A2(new_n279), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n261), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT10), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n260), .B1(new_n280), .B2(G169), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n282), .A2(G179), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n262), .A2(G232), .A3(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n262), .A2(G226), .A3(new_n263), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G97), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n269), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n295));
  INV_X1    g0095(.A(new_n272), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G238), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n277), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(KEYINPUT13), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n293), .B2(new_n269), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT13), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT14), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT66), .B1(new_n303), .B2(new_n304), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT66), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n301), .A2(new_n309), .A3(KEYINPUT13), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(new_n304), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n308), .A2(new_n310), .A3(G179), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n301), .A2(KEYINPUT13), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n311), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n307), .A2(new_n312), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n258), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT12), .ZN(new_n319));
  INV_X1    g0119(.A(new_n256), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n202), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n256), .A2(KEYINPUT12), .A3(G68), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n318), .A2(new_n202), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n265), .B2(new_n248), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n325), .A2(KEYINPUT11), .A3(new_n244), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT11), .B1(new_n325), .B2(new_n244), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n317), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G107), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n266), .A2(new_n298), .B1(new_n331), .B2(new_n262), .ZN(new_n332));
  INV_X1    g0132(.A(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n337), .A2(new_n228), .A3(G1698), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n269), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n273), .B1(G244), .B2(new_n278), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G190), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G87), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT15), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(KEYINPUT15), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n248), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n350), .A2(new_n253), .B1(new_n207), .B2(new_n265), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n244), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n258), .A2(G77), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n352), .B(new_n353), .C1(G77), .C2(new_n256), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  INV_X1    g0156(.A(new_n341), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n354), .B1(new_n357), .B2(G169), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n341), .A2(G179), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n289), .A2(new_n330), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n244), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT7), .B1(new_n337), .B2(new_n207), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  AOI211_X1 g0166(.A(new_n366), .B(G20), .C1(new_n334), .C2(new_n336), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n201), .A2(new_n202), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n252), .A2(G159), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n364), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT68), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n366), .B1(new_n262), .B2(G20), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n373), .B1(new_n381), .B2(G68), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n378), .B1(new_n382), .B2(KEYINPUT16), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n202), .B1(new_n379), .B2(new_n380), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n384), .A2(KEYINPUT68), .A3(new_n376), .A4(new_n373), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n377), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT69), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n297), .B1(new_n277), .B2(new_n228), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n262), .A2(G226), .A3(G1698), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n262), .A2(G223), .A3(new_n263), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n333), .C2(new_n344), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(new_n269), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n342), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(G200), .B2(new_n392), .ZN(new_n394));
  INV_X1    g0194(.A(new_n247), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n320), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n318), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n386), .A2(new_n387), .A3(new_n394), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n368), .A2(KEYINPUT16), .A3(new_n374), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n382), .A2(new_n378), .A3(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n397), .B1(new_n405), .B2(new_n377), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n406), .A2(new_n387), .A3(KEYINPUT17), .A4(new_n394), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G179), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n392), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G169), .B2(new_n392), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT18), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n411), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n244), .B1(new_n382), .B2(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n403), .B2(new_n404), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n413), .B(new_n414), .C1(new_n416), .C2(new_n397), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n328), .B1(new_n314), .B2(G200), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n308), .A2(new_n310), .A3(G190), .A4(new_n311), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT67), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(KEYINPUT67), .A3(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n363), .A2(new_n419), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n334), .A2(new_n336), .A3(G244), .A4(new_n263), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G283), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n276), .B1(new_n435), .B2(KEYINPUT72), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n434), .A2(new_n433), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n432), .A4(new_n431), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n206), .A2(G45), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n295), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n269), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G257), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G200), .ZN(new_n449));
  INV_X1    g0249(.A(G97), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n320), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n206), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n256), .A2(new_n452), .A3(new_n215), .A4(new_n243), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n453), .A2(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(KEYINPUT71), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G97), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT70), .B(G107), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(new_n331), .A3(KEYINPUT6), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(KEYINPUT6), .B2(new_n450), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n458), .B(new_n460), .C1(KEYINPUT6), .C2(new_n450), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n207), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n331), .B1(new_n379), .B2(new_n380), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n253), .A2(new_n265), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n451), .B(new_n457), .C1(new_n467), .C2(new_n364), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n449), .B(new_n469), .C1(new_n342), .C2(new_n448), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n440), .A2(new_n409), .A3(new_n445), .A4(new_n447), .ZN(new_n471));
  INV_X1    g0271(.A(new_n445), .ZN(new_n472));
  INV_X1    g0272(.A(new_n447), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(new_n436), .C2(new_n439), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n471), .B(new_n468), .C1(new_n474), .C2(G169), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n298), .A2(new_n263), .ZN(new_n477));
  INV_X1    g0277(.A(G244), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G1698), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n334), .A2(new_n477), .A3(new_n336), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n333), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n276), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n276), .A2(G274), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G250), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n206), .B2(G45), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n276), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT73), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n295), .A2(new_n486), .B1(new_n276), .B2(new_n489), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT73), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G238), .A2(G1698), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n478), .B2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n482), .B1(new_n496), .B2(new_n262), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n493), .B(new_n494), .C1(new_n497), .C2(new_n276), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G169), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n492), .A2(new_n498), .A3(new_n409), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n207), .B1(new_n292), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n344), .A2(new_n450), .A3(new_n331), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n334), .A2(new_n336), .A3(new_n207), .A4(G68), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n503), .B1(new_n248), .B2(new_n450), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(new_n244), .B1(new_n320), .B2(new_n348), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n454), .A2(new_n455), .A3(new_n347), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT74), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n501), .B(new_n502), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n499), .A2(G200), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n454), .A2(new_n455), .A3(G87), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n492), .A2(new_n498), .A3(G190), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n516), .A2(new_n510), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n515), .A2(KEYINPUT75), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT75), .B1(new_n515), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n433), .B(new_n207), .C1(G33), .C2(new_n450), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n481), .A2(G20), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n244), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT20), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n244), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  MUX2_X1   g0329(.A(new_n256), .B(new_n453), .S(G116), .Z(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n334), .A2(new_n336), .A3(G264), .A4(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n334), .A2(new_n336), .A3(G257), .A4(new_n263), .ZN(new_n534));
  INV_X1    g0334(.A(G303), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n533), .B(new_n534), .C1(new_n535), .C2(new_n262), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n536), .A2(new_n269), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n442), .A2(new_n443), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n276), .B1(new_n538), .B2(new_n441), .ZN(new_n539));
  INV_X1    g0339(.A(G270), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n445), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT76), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n446), .A2(G270), .B1(new_n295), .B2(new_n444), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT76), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n536), .A2(new_n269), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(G200), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n542), .A2(new_n546), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n532), .B(new_n547), .C1(new_n548), .C2(new_n342), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n472), .B1(G264), .B2(new_n446), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n334), .A2(new_n336), .A3(G257), .A4(G1698), .ZN(new_n551));
  AND2_X1   g0351(.A1(KEYINPUT80), .A2(G294), .ZN(new_n552));
  NOR2_X1   g0352(.A1(KEYINPUT80), .A2(G294), .ZN(new_n553));
  OAI21_X1  g0353(.A(G33), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT79), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n262), .A2(new_n556), .A3(G250), .A4(new_n263), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n334), .A2(new_n336), .A3(G250), .A4(new_n263), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT79), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n269), .B1(new_n560), .B2(KEYINPUT81), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n557), .ZN(new_n562));
  INV_X1    g0362(.A(new_n555), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT81), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n550), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n334), .A2(new_n336), .A3(new_n207), .A4(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT22), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT22), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n262), .A2(new_n572), .A3(new_n207), .A4(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT23), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n331), .A3(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(KEYINPUT78), .A2(KEYINPUT24), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT78), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n574), .A2(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n585), .B(new_n580), .C1(new_n571), .C2(new_n573), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n244), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n320), .A2(new_n331), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT25), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n456), .B2(G107), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n587), .B(new_n590), .C1(new_n567), .C2(new_n342), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n549), .B1(new_n569), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n409), .B(new_n550), .C1(new_n561), .C2(new_n566), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(new_n590), .ZN(new_n594));
  INV_X1    g0394(.A(new_n550), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n276), .B1(new_n564), .B2(new_n565), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n560), .A2(KEYINPUT81), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n593), .B(new_n594), .C1(new_n598), .C2(G169), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n500), .B1(new_n529), .B2(new_n530), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT77), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n542), .A2(new_n600), .A3(new_n602), .A4(new_n546), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n543), .A2(G179), .A3(new_n545), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n532), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n542), .A2(new_n546), .A3(new_n600), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(KEYINPUT77), .A3(new_n601), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n599), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n592), .A2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n428), .A2(new_n476), .A3(new_n522), .A4(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n475), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n510), .A2(new_n511), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n500), .B1(new_n484), .B2(new_n491), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n502), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n510), .A2(new_n517), .A3(KEYINPUT82), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT82), .B1(new_n510), .B2(new_n517), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n484), .A2(new_n491), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n518), .B1(new_n356), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT26), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n520), .A2(new_n521), .A3(new_n475), .ZN(new_n624));
  XNOR2_X1  g0424(.A(KEYINPUT83), .B(KEYINPUT26), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n594), .B1(G190), .B2(new_n598), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n621), .B1(new_n628), .B2(new_n568), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(new_n609), .A3(new_n475), .A4(new_n470), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n615), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n428), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n288), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n330), .B1(new_n422), .B2(new_n362), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n412), .B(new_n417), .C1(new_n635), .C2(new_n408), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n634), .B1(new_n636), .B2(new_n285), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(G369));
  NAND2_X1  g0438(.A1(new_n606), .A2(new_n608), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n531), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n640), .B(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n549), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n594), .A2(new_n646), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n569), .B2(new_n591), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n599), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n599), .A2(new_n646), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n646), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n639), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n654), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n210), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n505), .A2(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n213), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  INV_X1    g0469(.A(G330), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n473), .B1(new_n436), .B2(new_n439), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n499), .A2(new_n604), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n598), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n598), .A2(new_n671), .A3(new_n672), .A4(KEYINPUT30), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n619), .A2(G179), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n548), .A2(new_n448), .A3(new_n567), .A4(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n679), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT31), .B1(new_n679), .B2(new_n646), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n610), .A2(new_n476), .A3(new_n522), .A4(new_n658), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n670), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n632), .A2(new_n658), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n475), .A2(new_n621), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n515), .A2(new_n519), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT75), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n515), .A2(new_n519), .A3(KEYINPUT75), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n612), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n689), .B1(new_n694), .B2(new_n625), .ZN(new_n695));
  INV_X1    g0495(.A(new_n615), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT84), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n612), .A2(KEYINPUT26), .A3(new_n622), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n624), .B2(new_n626), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT84), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n615), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(new_n701), .A3(new_n630), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .A3(new_n658), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n684), .B1(new_n687), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n669), .B1(new_n704), .B2(G1), .ZN(G364));
  AND2_X1   g0505(.A1(new_n207), .A2(G13), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n206), .B1(new_n706), .B2(G45), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n664), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n649), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n670), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n649), .A2(KEYINPUT85), .A3(G330), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT85), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n650), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n210), .A2(new_n262), .ZN(new_n716));
  INV_X1    g0516(.A(G355), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(G116), .B2(new_n210), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n210), .A2(new_n337), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT86), .Z(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n485), .B2(new_n214), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n238), .A2(new_n485), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n215), .B1(G20), .B2(new_n500), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n709), .B1(new_n724), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n728), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n207), .A2(new_n409), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n207), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n734), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(G311), .A2(new_n736), .B1(new_n739), .B2(G329), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n342), .A3(G200), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n733), .A2(G190), .A3(new_n356), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT87), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(KEYINPUT87), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n743), .B1(G322), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n337), .B1(new_n751), .B2(new_n535), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT89), .Z(new_n753));
  NAND2_X1  g0553(.A1(new_n733), .A2(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n342), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G326), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n552), .A2(new_n553), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n342), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n207), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n754), .A2(G190), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n757), .A2(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n750), .A2(new_n753), .A3(new_n756), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n749), .A2(G58), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n262), .B1(new_n735), .B2(new_n265), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n344), .A2(new_n751), .B1(new_n742), .B2(new_n331), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n766), .B(new_n767), .C1(G50), .C2(new_n755), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G97), .A2(new_n760), .B1(new_n761), .B2(G68), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n738), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT88), .B(KEYINPUT32), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n765), .A2(new_n768), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n732), .B1(new_n764), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n731), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n727), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n649), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n715), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT90), .ZN(G396));
  NAND2_X1  g0580(.A1(new_n362), .A2(KEYINPUT95), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT95), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n360), .B2(new_n361), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n359), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n658), .B(new_n785), .C1(new_n627), .C2(new_n631), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n632), .A2(new_n658), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n354), .A2(new_n646), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n781), .A2(new_n358), .A3(new_n788), .A4(new_n783), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n362), .A2(new_n646), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT96), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n786), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n684), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT97), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n709), .B1(new_n793), .B2(new_n794), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n728), .A2(new_n725), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n709), .B1(G77), .B2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n755), .A2(G137), .B1(new_n736), .B2(G159), .ZN(new_n802));
  INV_X1    g0602(.A(new_n761), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n251), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G143), .B2(new_n749), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT93), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n262), .B1(new_n738), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  INV_X1    g0610(.A(G50), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n759), .A2(new_n201), .B1(new_n751), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n742), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G68), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n807), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n803), .A2(new_n741), .B1(new_n735), .B2(new_n481), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT91), .ZN(new_n818));
  INV_X1    g0618(.A(new_n755), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n817), .A2(new_n818), .B1(new_n535), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n818), .B2(new_n817), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT92), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n262), .B1(new_n739), .B2(G311), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n450), .B2(new_n759), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n344), .A2(new_n742), .B1(new_n751), .B2(new_n331), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(new_n748), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n815), .A2(new_n816), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n801), .B1(new_n829), .B2(new_n728), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n726), .B2(new_n791), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n798), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  AND2_X1   g0633(.A1(new_n462), .A2(new_n463), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(KEYINPUT35), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(KEYINPUT35), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(G116), .A3(new_n216), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT36), .Z(new_n839));
  OR3_X1    g0639(.A1(new_n213), .A2(new_n265), .A3(new_n369), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n811), .A2(G68), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n206), .B(G13), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n427), .B1(new_n685), .B2(new_n686), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n844), .A2(KEYINPUT102), .A3(new_n703), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT102), .B1(new_n844), .B2(new_n703), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n637), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n784), .A2(new_n658), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n786), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n328), .A2(new_n646), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n329), .A2(new_n422), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n317), .B1(new_n424), .B2(new_n425), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n852), .A2(KEYINPUT98), .A3(new_n850), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT98), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n307), .A2(new_n312), .A3(new_n316), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n420), .A2(KEYINPUT67), .A3(new_n421), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT67), .B1(new_n420), .B2(new_n421), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n850), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n851), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n849), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n644), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n416), .B2(new_n397), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n408), .B2(new_n418), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n386), .A2(new_n398), .A3(new_n394), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n411), .B1(new_n386), .B2(new_n398), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(KEYINPUT99), .A3(new_n868), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n869), .A2(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n865), .A2(new_n868), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n875), .A2(KEYINPUT99), .A3(KEYINPUT37), .A4(new_n870), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n867), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n867), .B(KEYINPUT38), .C1(new_n874), .C2(new_n876), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n863), .A2(new_n881), .B1(new_n418), .B2(new_n644), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT100), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n879), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT101), .Z(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n329), .A2(new_n646), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n879), .A2(new_n880), .A3(new_n884), .A4(new_n887), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n847), .B(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n791), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n682), .B2(new_n683), .ZN(new_n896));
  INV_X1    g0696(.A(new_n880), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n872), .A2(new_n873), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n871), .A2(new_n868), .A3(new_n865), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n869), .A2(new_n873), .A3(new_n872), .A4(new_n871), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n902), .B2(new_n867), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n861), .B(new_n896), .C1(new_n897), .C2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n881), .A2(KEYINPUT40), .A3(new_n861), .A4(new_n896), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n682), .A2(new_n683), .ZN(new_n909));
  OR3_X1    g0709(.A1(new_n908), .A2(new_n427), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n427), .B2(new_n909), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(G330), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n894), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n206), .B2(new_n706), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n894), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n843), .B1(new_n914), .B2(new_n915), .ZN(G367));
  OAI21_X1  g0716(.A(new_n476), .B1(new_n469), .B2(new_n658), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n612), .A2(new_n646), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n917), .A2(KEYINPUT103), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT103), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n655), .A2(new_n659), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT42), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n921), .A2(new_n599), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n646), .B1(new_n926), .B2(new_n475), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n618), .A2(new_n646), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n622), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n696), .A2(new_n618), .A3(new_n646), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n928), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n929), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n936), .B(new_n937), .C1(new_n925), .C2(new_n927), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n657), .B2(new_n921), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n657), .A2(new_n921), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n664), .B(new_n943), .Z(new_n944));
  INV_X1    g0744(.A(KEYINPUT106), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n655), .B2(new_n659), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(new_n923), .Z(new_n947));
  INV_X1    g0747(.A(KEYINPUT107), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(new_n650), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n712), .A2(new_n948), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(new_n714), .C1(new_n947), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n704), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n921), .A2(new_n660), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT44), .ZN(new_n955));
  XOR2_X1   g0755(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n956));
  NAND3_X1  g0756(.A1(new_n922), .A2(new_n661), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n921), .B2(new_n660), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n955), .A2(new_n656), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n656), .B1(new_n955), .B2(new_n960), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n944), .B1(new_n963), .B2(new_n704), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n940), .B(new_n942), .C1(new_n708), .C2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n709), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n720), .A2(new_n234), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n730), .B1(new_n663), .B2(new_n347), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n337), .B1(new_n738), .B2(new_n970), .C1(new_n741), .C2(new_n735), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n749), .B2(G303), .ZN(new_n972));
  INV_X1    g0772(.A(new_n751), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(G116), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n761), .A2(new_n757), .B1(new_n813), .B2(G97), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G107), .A2(new_n760), .B1(new_n755), .B2(G311), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n761), .A2(G159), .B1(new_n736), .B2(G50), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT108), .Z(new_n980));
  INV_X1    g0780(.A(G137), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n751), .A2(new_n201), .B1(new_n738), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n755), .A2(G143), .B1(new_n813), .B2(G77), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n337), .B1(new_n760), .B2(G68), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n748), .C2(new_n251), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n978), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT110), .Z(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n969), .B1(new_n933), .B2(new_n777), .C1(new_n990), .C2(new_n732), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n965), .A2(new_n991), .ZN(G387));
  OAI22_X1  g0792(.A1(new_n716), .A2(new_n666), .B1(G107), .B2(new_n210), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n350), .A2(G50), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT50), .Z(new_n995));
  OAI211_X1 g0795(.A(new_n666), .B(new_n485), .C1(new_n202), .C2(new_n265), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n720), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT111), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n231), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n997), .A2(new_n998), .B1(new_n1000), .B2(G45), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n993), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n709), .B1(new_n1002), .B2(new_n730), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n761), .A2(G311), .B1(new_n736), .B2(G303), .ZN(new_n1004));
  INV_X1    g0804(.A(G322), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1004), .B1(new_n1005), .B2(new_n819), .C1(new_n748), .C2(new_n970), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n760), .A2(G283), .B1(new_n973), .B2(new_n757), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT49), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n742), .A2(new_n481), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n262), .B(new_n1015), .C1(G326), .C2(new_n739), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n348), .A2(new_n759), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n819), .B2(new_n770), .C1(new_n247), .C2(new_n803), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n748), .A2(new_n811), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n262), .B1(new_n738), .B2(new_n251), .C1(new_n202), .C2(new_n735), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n265), .A2(new_n751), .B1(new_n742), .B2(new_n450), .ZN(new_n1023));
  OR4_X1    g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n732), .B1(new_n1017), .B2(new_n1024), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1003), .B(new_n1025), .C1(new_n655), .C2(new_n727), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n951), .B2(new_n708), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n952), .A2(new_n664), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n951), .A2(new_n704), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(G393));
  NAND3_X1  g0830(.A1(new_n961), .A2(new_n708), .A3(new_n962), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n729), .B1(new_n450), .B2(new_n210), .C1(new_n721), .C2(new_n241), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n709), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n748), .A2(new_n770), .B1(new_n251), .B2(new_n819), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT51), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n337), .B1(new_n739), .B2(G143), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n202), .B2(new_n751), .C1(new_n344), .C2(new_n742), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT112), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n735), .A2(new_n350), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n759), .A2(new_n265), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G50), .C2(new_n761), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1035), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n749), .A2(G311), .B1(G317), .B2(new_n755), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n803), .A2(new_n535), .B1(new_n742), .B2(new_n331), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n337), .B1(new_n738), .B2(new_n1005), .C1(new_n827), .C2(new_n735), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n759), .A2(new_n481), .B1(new_n751), .B2(new_n741), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1042), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1033), .B1(new_n1049), .B2(new_n728), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n922), .B2(new_n777), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1031), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(KEYINPUT113), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT113), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1031), .B2(new_n1051), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n961), .A2(new_n962), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n952), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n963), .A2(new_n664), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1053), .A2(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(G390));
  NAND2_X1  g0860(.A1(new_n428), .A2(new_n684), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n637), .B(new_n1061), .C1(new_n845), .C2(new_n846), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n702), .A2(new_n658), .A3(new_n785), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n848), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n861), .A2(new_n684), .A3(new_n791), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n861), .B1(new_n684), .B2(new_n792), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n861), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n794), .B2(new_n895), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1070), .A2(new_n1065), .B1(new_n786), .B2(new_n848), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1062), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n889), .A2(new_n891), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n890), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n862), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1069), .B1(new_n1063), .B2(new_n848), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n881), .A2(new_n1075), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1077), .B(new_n1065), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1064), .B2(new_n861), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n889), .A2(new_n891), .B1(new_n862), .B2(new_n1075), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1066), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n665), .B1(new_n1073), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1084), .B2(new_n1073), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1084), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1074), .A2(new_n725), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n709), .B1(new_n395), .B2(new_n800), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n337), .B1(new_n738), .B2(new_n827), .C1(new_n450), .C2(new_n735), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n202), .A2(new_n742), .B1(new_n751), .B2(new_n344), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n749), .C2(G116), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1040), .B1(G107), .B2(new_n761), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n741), .C2(new_n819), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT114), .Z(new_n1095));
  INV_X1    g0895(.A(G125), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT54), .B(G143), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n262), .B1(new_n738), .B2(new_n1096), .C1(new_n735), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n749), .B2(G132), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G159), .A2(new_n760), .B1(new_n761), .B2(G137), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n755), .A2(G128), .B1(new_n813), .B2(G50), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n751), .A2(new_n251), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT115), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n732), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1095), .A2(KEYINPUT115), .A3(new_n1104), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1089), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1087), .A2(new_n708), .B1(new_n1088), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1086), .A2(new_n1109), .ZN(G378));
  INV_X1    g0910(.A(new_n1062), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1084), .B2(new_n1072), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n906), .A2(G330), .A3(new_n907), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n260), .A2(new_n864), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n289), .B(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n906), .A2(new_n1117), .A3(G330), .A4(new_n907), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n893), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT120), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n892), .A3(new_n882), .A4(new_n1120), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(KEYINPUT120), .A3(new_n893), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1112), .A2(new_n1125), .A3(KEYINPUT57), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT57), .B1(new_n1112), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT121), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1127), .B(new_n664), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(KEYINPUT121), .B(KEYINPUT57), .C1(new_n1112), .C2(new_n1128), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n708), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1118), .A2(new_n725), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n709), .B1(G50), .B2(new_n800), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n819), .A2(new_n481), .B1(new_n202), .B2(new_n759), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT116), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n751), .A2(new_n265), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n742), .A2(new_n201), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(G97), .C2(new_n761), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n262), .A2(G41), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n741), .B2(new_n738), .C1(new_n348), .C2(new_n735), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n749), .B2(G107), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1138), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT58), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1142), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n811), .C1(G33), .C2(G41), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n748), .A2(new_n1151), .B1(new_n751), .B2(new_n1097), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT117), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n755), .A2(G125), .B1(new_n736), .B2(G137), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G150), .A2(new_n760), .B1(new_n761), .B2(G132), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT118), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n813), .A2(G159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G33), .B(G41), .C1(new_n739), .C2(G124), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1150), .B1(new_n1146), .B2(new_n1145), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1136), .B1(new_n1164), .B2(new_n728), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1135), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1134), .A2(KEYINPUT119), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT119), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n707), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1166), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1133), .A2(new_n1172), .ZN(G375));
  INV_X1    g0973(.A(new_n944), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1062), .A2(new_n1072), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1073), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n966), .B1(new_n202), .B2(new_n799), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n749), .A2(G137), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n262), .B1(new_n738), .B2(new_n1151), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G150), .B2(new_n736), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1140), .B1(G50), .B2(new_n760), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n755), .A2(G132), .B1(new_n973), .B2(G159), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n803), .C2(new_n1097), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n761), .A2(G116), .B1(new_n736), .B2(G107), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT122), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n337), .B1(new_n742), .B2(new_n265), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT123), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n755), .A2(G294), .B1(new_n973), .B2(G97), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1019), .B(new_n1189), .C1(new_n535), .C2(new_n738), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G283), .B2(new_n749), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1186), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1184), .A2(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1177), .B1(new_n732), .B2(new_n1193), .C1(new_n861), .C2(new_n726), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1072), .B2(new_n707), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1176), .A2(new_n1196), .ZN(G381));
  NOR2_X1   g0997(.A1(G375), .A2(G378), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR4_X1    g0999(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1200));
  OR4_X1    g1000(.A1(G387), .A2(new_n1199), .A3(G381), .A4(new_n1200), .ZN(G407));
  OAI211_X1 g1001(.A(G407), .B(G213), .C1(G343), .C2(new_n1199), .ZN(G409));
  INV_X1    g1002(.A(KEYINPUT61), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1073), .A2(KEYINPUT60), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1175), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1062), .A2(new_n1072), .A3(KEYINPUT60), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1206), .A2(new_n664), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G384), .B1(new_n1208), .B2(new_n1196), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1195), .B(new_n832), .C1(new_n1205), .C2(new_n1207), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n645), .A2(G213), .A3(G2897), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(G378), .B(new_n1172), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1112), .A2(new_n1174), .A3(new_n1128), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1125), .A2(new_n708), .A3(new_n1126), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1166), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n1086), .A3(new_n1109), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1214), .A2(new_n1218), .B1(G213), .B2(new_n645), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1203), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n645), .A2(G213), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1211), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT63), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G390), .A2(new_n965), .A3(new_n991), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G390), .B1(new_n965), .B2(new_n991), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT124), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(G393), .B(G396), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G390), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G387), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1227), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1231), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(KEYINPUT124), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1225), .A2(KEYINPUT63), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1221), .A2(new_n1226), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1219), .C2(new_n1211), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1224), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1222), .A2(KEYINPUT62), .A3(new_n1223), .A4(new_n1211), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1219), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1211), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1220), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1240), .B1(new_n1251), .B2(new_n1238), .ZN(G405));
  AOI21_X1  g1052(.A(new_n1236), .B1(new_n1235), .B2(KEYINPUT124), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1254), .B(new_n1231), .C1(new_n1234), .C2(new_n1227), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT127), .B(new_n1211), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1211), .A2(KEYINPUT127), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1232), .A2(new_n1237), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G378), .B1(new_n1133), .B2(new_n1172), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1214), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1260), .A2(new_n1261), .B1(KEYINPUT127), .B2(new_n1211), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1259), .B(new_n1262), .ZN(G402));
endmodule


