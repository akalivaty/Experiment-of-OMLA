//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(G41), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(KEYINPUT64), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT64), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G41), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT5), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n205), .A2(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n253), .B1(KEYINPUT5), .B2(new_n243), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n249), .A2(G274), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT5), .B1(new_n244), .B2(new_n246), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(new_n248), .B2(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(G270), .B(new_n252), .C1(new_n256), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n252), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G303), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  OAI211_X1 g0071(.A(G257), .B(new_n271), .C1(new_n264), .C2(new_n265), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT77), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT77), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(G257), .A4(new_n271), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT78), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n263), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI211_X1 g0079(.A(KEYINPUT78), .B(new_n270), .C1(new_n273), .C2(new_n276), .ZN(new_n280));
  OAI211_X1 g0080(.A(G190), .B(new_n262), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G116), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(new_n212), .B1(G20), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(G20), .B1(G33), .B2(G283), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G33), .B2(new_n219), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT20), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT79), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n288), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT79), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n284), .A2(new_n286), .A3(new_n291), .A4(KEYINPUT20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n282), .A2(new_n212), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n205), .A2(G33), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G116), .ZN(new_n299));
  INV_X1    g0099(.A(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(G116), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n266), .A2(new_n269), .ZN(new_n304));
  AOI21_X1  g0104(.A(G1698), .B1(new_n267), .B2(new_n268), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n275), .B1(new_n305), .B2(G257), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n272), .A2(KEYINPUT77), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n252), .B1(new_n308), .B2(KEYINPUT78), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n277), .A2(new_n278), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n261), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n281), .B(new_n303), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(G179), .A3(new_n302), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n262), .B1(new_n279), .B2(new_n280), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT21), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n293), .B2(new_n301), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n315), .B2(new_n318), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n313), .B(new_n314), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n302), .A2(G179), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n302), .A2(G169), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT21), .B1(new_n311), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT80), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n313), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n271), .B1(new_n267), .B2(new_n268), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n264), .A2(new_n265), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n332), .A2(G223), .B1(new_n333), .B2(G77), .ZN(new_n334));
  INV_X1    g0134(.A(G222), .ZN(new_n335));
  INV_X1    g0135(.A(new_n305), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n263), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT64), .B(G41), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n257), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n205), .A2(G274), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n243), .A2(new_n257), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n205), .A2(new_n344), .B1(new_n250), .B2(new_n251), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(G226), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G190), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G150), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n206), .A2(G33), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G50), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n206), .B1(new_n201), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n294), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n300), .A2(new_n294), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n205), .A2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(G50), .A3(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n356), .B(new_n359), .C1(G50), .C2(new_n296), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT9), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n361), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n348), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n347), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(G200), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT10), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT68), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n369), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT65), .B1(new_n347), .B2(G169), .ZN(new_n372));
  INV_X1    g0172(.A(G179), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n347), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT65), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n360), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n370), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n351), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(KEYINPUT66), .B2(new_n349), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(KEYINPUT66), .B2(new_n349), .ZN(new_n382));
  INV_X1    g0182(.A(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT15), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT15), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G87), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G77), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n352), .B1(new_n206), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n294), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n205), .B2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n357), .A2(new_n392), .B1(new_n389), .B2(new_n300), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n332), .A2(G238), .B1(new_n333), .B2(G107), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n218), .B2(new_n336), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n263), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n343), .B1(G244), .B2(new_n345), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n394), .B1(new_n400), .B2(G190), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n312), .B2(new_n400), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n399), .A2(new_n317), .B1(new_n391), .B2(new_n393), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n373), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT67), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G68), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n349), .A2(G50), .B1(G20), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n389), .B2(new_n352), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT11), .B1(new_n411), .B2(new_n294), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT69), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n300), .A2(new_n409), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n357), .A2(G68), .A3(new_n358), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n414), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT69), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n412), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n415), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n218), .A2(G1698), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n274), .B(new_n425), .C1(G226), .C2(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n263), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n345), .A2(G238), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n342), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n252), .B1(new_n426), .B2(new_n427), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n342), .A2(new_n430), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT13), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT14), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(G169), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n433), .A2(G179), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n437), .B2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n424), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n437), .A2(G200), .ZN(new_n444));
  INV_X1    g0244(.A(G190), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n423), .B(new_n444), .C1(new_n445), .C2(new_n437), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n402), .A2(KEYINPUT67), .A3(new_n405), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n408), .A2(new_n443), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n217), .A2(new_n409), .ZN(new_n449));
  OAI21_X1  g0249(.A(G20), .B1(new_n449), .B2(new_n201), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n349), .A2(G159), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT7), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n274), .B2(G20), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n333), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT70), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(G68), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(KEYINPUT16), .B(new_n453), .C1(new_n458), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT16), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n409), .B1(new_n455), .B2(new_n456), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(new_n452), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n294), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n357), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n380), .A2(new_n358), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n467), .A2(new_n468), .B1(new_n296), .B2(new_n380), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n345), .A2(G232), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n342), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G226), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G1698), .ZN(new_n475));
  OAI221_X1 g0275(.A(new_n475), .B1(G223), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G87), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n252), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(G169), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n263), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n340), .A2(new_n341), .B1(new_n345), .B2(G232), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(G179), .A3(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n471), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT18), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n473), .A2(new_n478), .A3(new_n445), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n312), .B1(new_n481), .B2(new_n482), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n466), .A2(new_n490), .A3(new_n470), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT17), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n484), .B1(new_n466), .B2(new_n470), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT18), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n466), .A2(new_n490), .A3(new_n470), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n487), .A2(new_n492), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n379), .A2(new_n448), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT76), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n298), .A2(KEYINPUT72), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT72), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n357), .A2(new_n503), .A3(new_n297), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n504), .A3(G87), .ZN(new_n505));
  NAND3_X1  g0305(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n206), .ZN(new_n507));
  INV_X1    g0307(.A(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n383), .A2(new_n219), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n206), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n352), .B2(new_n219), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n294), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n387), .A2(new_n296), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT75), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT75), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n519), .B(new_n516), .C1(new_n514), .C2(new_n294), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n505), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT74), .ZN(new_n522));
  AND2_X1   g0322(.A1(G33), .A2(G41), .ZN(new_n523));
  OAI21_X1  g0323(.A(G274), .B1(new_n523), .B2(new_n212), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n524), .B2(new_n253), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n252), .A2(KEYINPUT74), .A3(G274), .A4(new_n258), .ZN(new_n526));
  INV_X1    g0326(.A(G250), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n258), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n525), .A2(new_n526), .B1(new_n252), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n530));
  OAI211_X1 g0330(.A(G238), .B(new_n271), .C1(new_n264), .C2(new_n265), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n263), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n312), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n501), .B1(new_n521), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n515), .A2(new_n517), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n519), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n515), .A2(KEYINPUT75), .A3(new_n517), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n535), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(KEYINPUT76), .A3(new_n541), .A4(new_n505), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n529), .A2(new_n534), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(new_n445), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n502), .A2(new_n504), .A3(new_n387), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n543), .A2(G169), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n529), .A2(G179), .A3(new_n534), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n349), .A2(KEYINPUT71), .A3(G77), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT71), .B1(new_n349), .B2(G77), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n557), .A2(new_n219), .A3(G107), .ZN(new_n558));
  XNOR2_X1  g0358(.A(G97), .B(G107), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n556), .B1(new_n560), .B2(new_n206), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n508), .B1(new_n455), .B2(new_n456), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n294), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n502), .A2(new_n504), .A3(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n300), .A2(new_n219), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G257), .B(new_n252), .C1(new_n256), .C2(new_n259), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n255), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n332), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT73), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(new_n271), .C1(new_n264), .C2(new_n265), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n305), .A2(KEYINPUT73), .A3(KEYINPUT4), .A4(G244), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n572), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n568), .B1(new_n576), .B2(new_n263), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G190), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n566), .B(new_n578), .C1(new_n312), .C2(new_n577), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n373), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(G169), .C2(new_n577), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n553), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n527), .A2(new_n271), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n220), .A2(G1698), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n264), .C2(new_n265), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n252), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n263), .B1(new_n249), .B2(new_n254), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(G264), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n317), .B1(new_n591), .B2(new_n255), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(new_n588), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n263), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(new_n252), .C1(new_n256), .C2(new_n259), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n255), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n373), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT82), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n508), .A2(KEYINPUT23), .A3(G20), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT23), .B1(new_n508), .B2(G20), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(new_n600), .B1(G20), .B2(new_n532), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n206), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n274), .A2(new_n604), .A3(new_n206), .A4(G87), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT24), .B(new_n601), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT24), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n605), .ZN(new_n608));
  INV_X1    g0408(.A(new_n601), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n294), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n502), .A2(new_n504), .A3(G107), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n205), .A2(new_n508), .A3(G13), .A4(G20), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT25), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT81), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n615), .B(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n596), .A2(G169), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT82), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n373), .C2(new_n596), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n598), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n591), .A2(G190), .A3(new_n255), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n596), .A2(G200), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n611), .A2(new_n618), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n331), .A2(new_n500), .A3(new_n584), .A4(new_n627), .ZN(G372));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT83), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n521), .B2(new_n535), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n540), .A2(KEYINPUT83), .A3(new_n541), .A4(new_n505), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n632), .A3(new_n545), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n552), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n629), .B1(new_n634), .B2(new_n582), .ZN(new_n635));
  INV_X1    g0435(.A(new_n582), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n546), .A2(new_n636), .A3(KEYINPUT26), .A4(new_n552), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n619), .B1(new_n592), .B2(new_n597), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n328), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n548), .A2(new_n551), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n540), .A2(new_n541), .A3(new_n505), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n544), .B1(new_n642), .B2(new_n630), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n632), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n579), .A2(new_n582), .A3(new_n626), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n552), .B(KEYINPUT84), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n500), .B1(new_n638), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n378), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n370), .A2(new_n371), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n493), .B(KEYINPUT18), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n446), .A2(new_n403), .A3(new_n404), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n443), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n496), .B(KEYINPUT17), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n651), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n650), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n303), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n329), .B1(new_n328), .B2(new_n313), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n328), .A2(new_n670), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n619), .A2(new_n667), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n623), .A2(new_n626), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n623), .B2(new_n668), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n676), .A2(KEYINPUT86), .A3(G330), .A4(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n322), .B2(new_n330), .ZN(new_n681));
  OAI211_X1 g0481(.A(G330), .B(new_n679), .C1(new_n681), .C2(new_n674), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT86), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n627), .A2(new_n686), .A3(new_n668), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n639), .A2(new_n667), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(KEYINPUT87), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n685), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n209), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n247), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n509), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n215), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT88), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n623), .A2(new_n626), .A3(new_n668), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n553), .A2(new_n703), .A3(new_n583), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n671), .B2(new_n672), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n529), .A2(G179), .A3(new_n534), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n577), .A2(new_n707), .A3(new_n591), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n708), .B2(new_n315), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n594), .A2(new_n595), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n550), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n311), .A2(KEYINPUT30), .A3(new_n577), .A4(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n543), .A2(new_n373), .A3(new_n596), .ZN(new_n713));
  INV_X1    g0513(.A(new_n577), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n315), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT31), .B1(new_n716), .B2(new_n667), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n705), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n702), .B1(new_n721), .B2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  AOI211_X1 g0523(.A(KEYINPUT88), .B(new_n723), .C1(new_n705), .C2(new_n720), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n328), .A2(new_n623), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n644), .A3(new_n646), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT26), .B1(new_n634), .B2(new_n582), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n546), .A2(new_n636), .A3(new_n629), .A4(new_n552), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n727), .A2(new_n648), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .A3(new_n668), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n641), .B(KEYINPUT84), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n634), .A2(new_n645), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(new_n640), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n635), .A2(new_n637), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n667), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n731), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n725), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n701), .B1(new_n738), .B2(G1), .ZN(G364));
  INV_X1    g0539(.A(G13), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n205), .B1(new_n741), .B2(G45), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n697), .A2(KEYINPUT89), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT89), .ZN(new_n744));
  INV_X1    g0544(.A(new_n742), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n696), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n676), .B2(G330), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G330), .B2(new_n676), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n212), .B1(G20), .B2(new_n317), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n206), .A2(G179), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G190), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(G20), .A2(G179), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n753), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G329), .A2(new_n755), .B1(new_n759), .B2(G311), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n756), .A2(new_n445), .A3(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n274), .B1(G322), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(new_n445), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G317), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT33), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n765), .A2(KEYINPUT33), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n760), .A2(new_n762), .A3(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT92), .B(G326), .Z(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n756), .A2(new_n445), .A3(new_n312), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n373), .A2(new_n312), .A3(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(new_n772), .B1(G294), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT93), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT94), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n752), .A2(new_n445), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT91), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n769), .B(new_n782), .C1(G283), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n274), .B1(new_n763), .B2(new_n409), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n755), .A2(G159), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(KEYINPUT32), .B2(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G50), .A2(new_n772), .B1(new_n761), .B2(G58), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(new_n389), .C2(new_n758), .ZN(new_n794));
  INV_X1    g0594(.A(new_n774), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n219), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n797), .B1(new_n383), .B2(new_n779), .C1(new_n791), .C2(KEYINPUT32), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n794), .B(new_n798), .C1(G107), .C2(new_n788), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n751), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n695), .A2(new_n333), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT90), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G355), .B1(new_n283), .B2(new_n695), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n241), .A2(new_n257), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n695), .A2(new_n274), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G45), .B2(new_n215), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n751), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n747), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n811), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n800), .B(new_n813), .C1(new_n676), .C2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n750), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  AOI211_X1 g0617(.A(new_n274), .B(new_n796), .C1(G294), .C2(new_n761), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n780), .A2(G107), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n788), .A2(G87), .ZN(new_n820));
  INV_X1    g0620(.A(new_n772), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n778), .B1(new_n754), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT95), .B(G283), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n763), .A2(new_n824), .B1(new_n758), .B2(new_n283), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  INV_X1    g0628(.A(G159), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n763), .A2(new_n828), .B1(new_n758), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n821), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n830), .B(new_n832), .C1(G143), .C2(new_n761), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n333), .B1(new_n755), .B2(G132), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(new_n217), .C2(new_n795), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n788), .A2(G68), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n354), .B2(new_n781), .C1(new_n833), .C2(KEYINPUT34), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n827), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n751), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n751), .A2(new_n809), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n747), .B1(new_n389), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n405), .A2(new_n667), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n394), .A2(new_n667), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n402), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n405), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n840), .B(new_n842), .C1(new_n846), .C2(new_n810), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n736), .B(new_n846), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n848), .A2(new_n725), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT96), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n747), .C1(new_n725), .C2(new_n848), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n849), .A2(KEYINPUT96), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n741), .A2(new_n205), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT100), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n623), .A2(new_n626), .A3(new_n668), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n579), .A2(new_n582), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n552), .A4(new_n546), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n330), .B2(new_n322), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n716), .A2(new_n667), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT31), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n717), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n855), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT7), .B1(new_n333), .B2(new_n206), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n409), .B1(new_n866), .B2(new_n459), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n452), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n295), .B1(new_n869), .B2(KEYINPUT16), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n453), .B1(new_n458), .B2(new_n461), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n463), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n469), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n496), .B1(new_n873), .B2(new_n665), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n484), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n665), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n471), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n486), .A2(new_n878), .A3(new_n879), .A4(new_n496), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n873), .A2(new_n665), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n653), .B2(new_n656), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n865), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n499), .A2(new_n882), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n876), .A2(new_n880), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n846), .ZN(new_n890));
  INV_X1    g0690(.A(new_n442), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n446), .A2(new_n440), .A3(new_n891), .A4(new_n439), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT99), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n423), .A2(new_n668), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n443), .B(new_n446), .C1(new_n423), .C2(new_n668), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n890), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n705), .A2(KEYINPUT100), .A3(new_n720), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n864), .A2(new_n889), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n491), .A2(new_n493), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n879), .B1(new_n905), .B2(new_n878), .ZN(new_n906));
  INV_X1    g0706(.A(new_n880), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n878), .B1(new_n653), .B2(new_n656), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n865), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n903), .B1(new_n910), .B2(new_n888), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(new_n864), .A3(new_n900), .A4(new_n901), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n705), .A2(KEYINPUT100), .A3(new_n720), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT100), .B1(new_n705), .B2(new_n720), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n916), .A2(new_n500), .ZN(new_n917));
  OAI21_X1  g0717(.A(G330), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT101), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n913), .A2(new_n917), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n895), .A2(new_n896), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n898), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n668), .B(new_n846), .C1(new_n638), .C2(new_n649), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n843), .B(KEYINPUT98), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n889), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n665), .B1(new_n466), .B2(new_n470), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n499), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n486), .A2(new_n878), .A3(new_n496), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT37), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n880), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n931), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n443), .A2(new_n667), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n939), .B(new_n941), .C1(new_n931), .C2(new_n889), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n653), .A2(new_n877), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n930), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n500), .B(new_n731), .C1(KEYINPUT29), .C2(new_n736), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n945), .A2(new_n659), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n854), .B1(new_n923), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n923), .ZN(new_n949));
  INV_X1    g0749(.A(new_n560), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n283), .B(new_n214), .C1(new_n950), .C2(KEYINPUT35), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(KEYINPUT35), .B2(new_n950), .ZN(new_n952));
  XOR2_X1   g0752(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n215), .A2(new_n389), .A3(new_n449), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n409), .A2(G50), .ZN(new_n956));
  OAI211_X1 g0756(.A(G1), .B(new_n740), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n954), .A3(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n806), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n812), .B1(new_n209), .B2(new_n388), .C1(new_n959), .C2(new_n234), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n748), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n751), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n788), .A2(G77), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n274), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G159), .A2(new_n764), .B1(new_n755), .B2(G137), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n354), .B2(new_n758), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n779), .A2(new_n217), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n795), .A2(new_n409), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n772), .A2(G143), .ZN(new_n970));
  INV_X1    g0770(.A(new_n761), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n971), .B2(new_n828), .ZN(new_n972));
  NOR4_X1   g0772(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n788), .A2(G97), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT46), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n779), .B2(new_n283), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n274), .B1(new_n755), .B2(G317), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n821), .A2(new_n822), .B1(new_n971), .B2(new_n778), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G294), .B2(new_n764), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n976), .A2(new_n978), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT107), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n795), .A2(new_n508), .B1(new_n758), .B2(new_n824), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT106), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n983), .A2(KEYINPUT107), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n974), .A2(new_n975), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT47), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n667), .A2(new_n521), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n644), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT102), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT102), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n648), .C2(new_n991), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n961), .B1(new_n962), .B2(new_n990), .C1(new_n995), .C2(new_n814), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n857), .B1(new_n566), .B2(new_n668), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n636), .A2(new_n667), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n1000));
  NAND3_X1  g0800(.A1(new_n693), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1000), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n687), .A2(KEYINPUT87), .A3(new_n688), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT87), .B1(new_n687), .B2(new_n688), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n999), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT44), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  NOR4_X1   g0809(.A1(new_n1003), .A2(new_n1004), .A3(new_n1009), .A4(new_n999), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1001), .B(new_n1007), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT105), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n680), .A2(new_n684), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n680), .A2(new_n684), .A3(new_n1012), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1009), .B1(new_n693), .B2(new_n999), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n1006), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1018), .A3(new_n1001), .A4(new_n1007), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n721), .A2(new_n702), .A3(G330), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n328), .A2(new_n667), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n687), .B1(new_n679), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n674), .B1(new_n331), .B2(new_n670), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(new_n723), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1022), .B(G330), .C1(new_n681), .C2(new_n674), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n863), .B1(new_n331), .B2(new_n704), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT88), .B1(new_n1028), .B2(new_n723), .ZN(new_n1029));
  AND4_X1   g0829(.A1(new_n1020), .A2(new_n1027), .A3(new_n737), .A4(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1014), .A2(new_n1019), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n738), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n696), .B(KEYINPUT41), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n745), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n999), .A2(new_n627), .A3(new_n1021), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n582), .B1(new_n997), .B2(new_n623), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(KEYINPUT42), .B1(new_n1037), .B2(new_n668), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(KEYINPUT42), .B2(new_n1036), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n680), .A2(new_n684), .A3(new_n999), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT103), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT103), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n680), .A2(new_n684), .A3(new_n1045), .A4(new_n999), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1044), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1041), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n996), .B1(new_n1035), .B2(new_n1056), .ZN(G387));
  OAI21_X1  g0857(.A(new_n806), .B1(new_n231), .B2(new_n257), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n698), .B2(new_n802), .ZN(new_n1059));
  OR3_X1    g0859(.A1(new_n351), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT50), .B1(new_n351), .B2(G50), .ZN(new_n1061));
  AOI21_X1  g0861(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1060), .A2(new_n698), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1059), .A2(new_n1063), .B1(new_n508), .B2(new_n695), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n812), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n748), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n795), .A2(new_n388), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n333), .B(new_n1067), .C1(G150), .C2(new_n755), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n821), .A2(new_n829), .B1(new_n971), .B2(new_n354), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n763), .A2(new_n351), .B1(new_n758), .B2(new_n409), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n779), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(G77), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n976), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n824), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1072), .A2(G294), .B1(new_n1075), .B2(new_n774), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G322), .A2(new_n772), .B1(new_n761), .B2(G317), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n778), .B2(new_n758), .C1(new_n822), .C2(new_n763), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT109), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(KEYINPUT49), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n274), .B1(new_n771), .B2(new_n755), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n283), .C2(new_n787), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT49), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1074), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1066), .B1(new_n1087), .B2(new_n751), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n679), .B2(new_n814), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1089), .A2(KEYINPUT110), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(KEYINPUT110), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1090), .A2(new_n1091), .B1(new_n745), .B2(new_n1027), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1030), .A2(new_n697), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n738), .A2(new_n1027), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(G393));
  XNOR2_X1  g0895(.A(new_n1011), .B(new_n685), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n696), .B(new_n1031), .C1(new_n1096), .C2(new_n1030), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1006), .A2(new_n811), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n812), .B1(new_n219), .B2(new_n209), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n806), .B2(new_n238), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n333), .B1(new_n755), .B2(G143), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n820), .B(new_n1101), .C1(new_n409), .C2(new_n779), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT112), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n821), .A2(new_n828), .B1(new_n971), .B2(new_n829), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n795), .A2(new_n389), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n763), .A2(new_n354), .B1(new_n758), .B2(new_n351), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G317), .A2(new_n772), .B1(new_n761), .B2(G311), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT52), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n788), .A2(G107), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n274), .B1(new_n759), .B2(G294), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G303), .A2(new_n764), .B1(new_n755), .B2(G322), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1072), .A2(new_n1075), .B1(new_n774), .B2(G116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1103), .A2(new_n1111), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT113), .Z(new_n1120));
  AOI211_X1 g0920(.A(new_n747), .B(new_n1100), .C1(new_n1120), .C2(new_n751), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1096), .A2(new_n745), .B1(new_n1098), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1097), .A2(new_n1122), .ZN(G390));
  NAND4_X1  g0923(.A1(new_n864), .A2(G330), .A3(new_n846), .A4(new_n901), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n925), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n925), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n846), .B(new_n1126), .C1(new_n722), .C2(new_n724), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n730), .A2(new_n668), .A3(new_n846), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n928), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n846), .B1(new_n722), .B2(new_n724), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n914), .A2(new_n915), .A3(new_n723), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1132), .A2(new_n925), .B1(new_n1133), .B2(new_n900), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n926), .A2(new_n928), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1131), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1133), .A2(new_n500), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n659), .A3(new_n945), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n939), .B1(new_n931), .B2(new_n889), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n929), .B2(new_n941), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1129), .A2(new_n1126), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n940), .B(KEYINPUT114), .Z(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n888), .B2(new_n910), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1147), .A3(new_n1127), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n916), .A2(G330), .A3(new_n900), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1141), .A2(new_n1151), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1143), .A2(new_n1147), .A3(new_n1127), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1150), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n1140), .A3(new_n1137), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(new_n1156), .A3(new_n696), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT115), .B1(new_n1151), .B2(new_n742), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT115), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1155), .A2(new_n1159), .A3(new_n745), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1142), .A2(new_n809), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n747), .B1(new_n351), .B2(new_n841), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n758), .A2(new_n219), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n971), .A2(new_n283), .B1(new_n763), .B2(new_n508), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(G283), .C2(new_n772), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n274), .B(new_n1108), .C1(G294), .C2(new_n755), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n780), .A2(G87), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n837), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(G132), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n971), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(G128), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT54), .B(G143), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n821), .A2(new_n1172), .B1(new_n758), .B2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1171), .B(new_n1174), .C1(G125), .C2(new_n755), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n788), .A2(G50), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n274), .B1(new_n763), .B2(new_n831), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G159), .B2(new_n774), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n779), .A2(new_n828), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT53), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .A4(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1169), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1162), .B(new_n1163), .C1(new_n962), .C2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1157), .A2(new_n1161), .A3(new_n1183), .ZN(G378));
  INV_X1    g0984(.A(KEYINPUT117), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n877), .A2(new_n360), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT116), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n379), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n370), .A2(new_n371), .A3(new_n378), .A4(new_n1187), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1189), .A2(new_n1192), .A3(new_n1190), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n902), .A2(new_n903), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n912), .A2(G330), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n846), .B1(new_n924), .B2(new_n898), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n914), .A2(new_n915), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n723), .B1(new_n1201), .B2(new_n911), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n904), .A3(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1199), .A2(new_n944), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n944), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1185), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n944), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1197), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1203), .B1(new_n1202), .B2(new_n904), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1199), .A2(new_n1204), .A3(new_n944), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(KEYINPUT117), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1139), .B1(new_n1155), .B2(new_n1137), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT57), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n696), .B1(new_n1219), .B2(new_n1215), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n333), .A2(new_n339), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n354), .C1(G33), .C2(G41), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n755), .C2(G124), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n764), .A2(G132), .B1(new_n772), .B2(G125), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n1172), .B2(new_n971), .C1(new_n831), .C2(new_n758), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n795), .A2(new_n828), .B1(new_n779), .B2(new_n1173), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT59), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1224), .B1(new_n829), .B2(new_n787), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1228), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1223), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1222), .B(new_n969), .C1(G283), .C2(new_n755), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n788), .A2(G58), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n388), .A2(new_n758), .B1(new_n971), .B2(new_n508), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n821), .A2(new_n283), .B1(new_n219), .B2(new_n763), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n1073), .A3(new_n1235), .A4(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT58), .Z(new_n1240));
  OAI21_X1  g1040(.A(new_n751), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n747), .B1(new_n354), .B2(new_n841), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n1203), .C2(new_n810), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1214), .B2(new_n745), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1221), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(G375));
  OAI211_X1 g1047(.A(new_n1139), .B(new_n1131), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1141), .A2(new_n1034), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n925), .A2(new_n809), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n751), .A2(G68), .A3(new_n809), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n780), .A2(G159), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n821), .A2(new_n1170), .B1(new_n758), .B2(new_n828), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n971), .A2(new_n831), .B1(new_n754), .B2(new_n1172), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n274), .B1(new_n763), .B2(new_n1173), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G50), .B2(new_n774), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1235), .A2(new_n1252), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n274), .B(new_n1067), .C1(G283), .C2(new_n761), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n754), .A2(new_n778), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n763), .A2(new_n283), .B1(new_n758), .B2(new_n508), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(G294), .C2(new_n772), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n963), .A3(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n781), .A2(new_n219), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n747), .B(new_n1251), .C1(new_n1265), .C2(new_n751), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1137), .A2(new_n745), .B1(new_n1250), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1249), .A2(new_n1267), .ZN(G381));
  OR4_X1    g1068(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(new_n1269), .A2(G378), .A3(G387), .A4(G381), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1246), .A2(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT118), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(KEYINPUT118), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1272), .A2(new_n1273), .ZN(G407));
  INV_X1    g1074(.A(G213), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G378), .A2(G343), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1246), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT119), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(G409));
  INV_X1    g1080(.A(KEYINPUT123), .ZN(new_n1281));
  INV_X1    g1081(.A(G390), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(G387), .B2(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(G393), .B(new_n816), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1033), .B1(new_n1031), .B2(new_n738), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1055), .B(new_n1049), .C1(new_n1285), .C2(new_n745), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(G390), .A3(new_n996), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G390), .B1(new_n1286), .B2(new_n996), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1283), .A2(new_n1284), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1284), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G387), .A2(new_n1282), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  XOR2_X1   g1094(.A(new_n1294), .B(KEYINPUT126), .Z(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1245), .C1(new_n1217), .C2(new_n1220), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1157), .A2(new_n1161), .A3(new_n1183), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1033), .B(new_n1215), .C1(new_n1207), .C2(new_n1213), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1218), .A2(new_n745), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1243), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1297), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n890), .B1(new_n1029), .B2(new_n1020), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1150), .B1(new_n1303), .B2(new_n1126), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1129), .B1(new_n1124), .B2(new_n925), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1304), .A2(new_n1135), .B1(new_n1127), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT60), .B1(new_n1306), .B2(new_n1139), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1139), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT120), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1248), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n697), .B1(new_n1311), .B2(KEYINPUT121), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT121), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1248), .B2(new_n1310), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1248), .A2(new_n1310), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT120), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(new_n1316), .A3(new_n1141), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1309), .A2(new_n1312), .A3(new_n1314), .A4(new_n1317), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1318), .A2(G384), .A3(new_n1267), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G384), .B1(new_n1318), .B2(new_n1267), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n666), .A2(G213), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1302), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n1296), .A2(new_n1301), .B1(G213), .B2(new_n666), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n666), .A2(G213), .A3(G2897), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1329));
  INV_X1    g1129(.A(G384), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1306), .A2(KEYINPUT121), .A3(KEYINPUT60), .A4(new_n1139), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1314), .A2(new_n1331), .A3(new_n696), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1315), .A2(new_n1316), .A3(new_n1141), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1316), .B1(new_n1315), .B2(new_n1141), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1332), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1267), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1330), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1318), .A2(G384), .A3(new_n1267), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(new_n1338), .A3(new_n1327), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1329), .A2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1324), .B(new_n1325), .C1(new_n1326), .C2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1323), .A2(KEYINPUT122), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT122), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1326), .A2(new_n1343), .A3(new_n1321), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT62), .B1(new_n1342), .B2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1295), .B1(new_n1341), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT125), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1340), .A2(new_n1326), .ZN(new_n1348));
  AND4_X1   g1148(.A1(KEYINPUT63), .A2(new_n1302), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1342), .A2(new_n1351), .A3(new_n1344), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT124), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1353), .B1(new_n1294), .B2(new_n1325), .ZN(new_n1354));
  AOI211_X1 g1154(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n1290), .C2(new_n1293), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  AND4_X1   g1157(.A1(new_n1347), .A2(new_n1350), .A3(new_n1352), .A4(new_n1357), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1302), .A2(new_n1321), .A3(KEYINPUT63), .A4(new_n1322), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1359), .B1(new_n1326), .B2(new_n1340), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1360), .A2(new_n1356), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1347), .B1(new_n1361), .B2(new_n1352), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1346), .B1(new_n1358), .B2(new_n1362), .ZN(G405));
  INV_X1    g1163(.A(new_n1321), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1364), .A2(KEYINPUT127), .ZN(new_n1365));
  XNOR2_X1  g1165(.A(new_n1365), .B(new_n1294), .ZN(new_n1366));
  XNOR2_X1  g1166(.A(new_n1246), .B(new_n1297), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(new_n1366), .B(new_n1367), .ZN(G402));
endmodule


