//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT64), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G97), .A2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT67), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n218), .B(new_n219), .C1(G77), .C2(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G116), .A2(G270), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(new_n234));
  AOI211_X1 g0034(.A(new_n212), .B(new_n228), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  OR2_X1    g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(new_n230), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n252), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n222), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n222), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n259), .B2(new_n201), .ZN(new_n260));
  INV_X1    g0060(.A(G159), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT74), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT16), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n229), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT16), .ZN(new_n269));
  OAI211_X1 g0069(.A(KEYINPUT74), .B(new_n269), .C1(new_n257), .C2(new_n264), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n230), .A2(G1), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT75), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n267), .A2(new_n229), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(new_n274), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n271), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n251), .A2(new_n252), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n221), .A2(G1698), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(G223), .C2(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G87), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n284), .A2(new_n290), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n293), .A2(G232), .ZN(new_n294));
  OR3_X1    g0094(.A1(new_n289), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(G200), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n282), .A2(KEYINPUT17), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT17), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n271), .A2(new_n299), .A3(new_n276), .A4(new_n281), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n297), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n271), .A2(new_n276), .A3(new_n281), .ZN(new_n304));
  NOR4_X1   g0104(.A1(new_n289), .A2(new_n294), .A3(G179), .A4(new_n292), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n295), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(KEYINPUT18), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT18), .B1(new_n304), .B2(new_n307), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n300), .B(new_n303), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n221), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G232), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G1698), .ZN(new_n317));
  AND2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n315), .B(new_n317), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n292), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n284), .A2(G238), .A3(new_n290), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n313), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n284), .B1(new_n320), .B2(new_n321), .ZN(new_n328));
  NOR4_X1   g0128(.A1(new_n328), .A2(KEYINPUT13), .A3(new_n325), .A4(new_n292), .ZN(new_n329));
  OAI21_X1  g0129(.A(G169), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT14), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n327), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  AND4_X1   g0133(.A1(new_n332), .A2(new_n324), .A3(new_n313), .A4(new_n326), .ZN(new_n334));
  OAI21_X1  g0134(.A(G179), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(KEYINPUT14), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G33), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G77), .B1(new_n262), .B2(G50), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n230), .B2(G68), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n268), .ZN(new_n342));
  XOR2_X1   g0142(.A(new_n342), .B(KEYINPUT11), .Z(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n275), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n274), .A2(G68), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n268), .A2(KEYINPUT72), .A3(new_n277), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n348), .B1(KEYINPUT12), .B2(new_n349), .C1(new_n222), .C2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n337), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT69), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G222), .A2(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G223), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G1698), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n357), .A2(new_n359), .B1(new_n251), .B2(new_n252), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n318), .A2(new_n319), .A3(G77), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n314), .A2(G223), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n363), .A2(new_n356), .B1(new_n318), .B2(new_n319), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(KEYINPUT69), .C1(G77), .C2(new_n285), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n365), .A3(new_n323), .ZN(new_n366));
  INV_X1    g0166(.A(new_n292), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n293), .A2(G226), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n306), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n203), .A2(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n262), .A2(G150), .ZN(new_n372));
  INV_X1    g0172(.A(new_n339), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n372), .C1(new_n272), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n268), .ZN(new_n375));
  OAI21_X1  g0175(.A(G50), .B1(new_n268), .B2(new_n277), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT70), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n274), .A2(new_n202), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n366), .A2(new_n382), .A3(new_n367), .A4(new_n368), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n370), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT9), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n375), .B(KEYINPUT9), .C1(new_n379), .C2(new_n380), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT10), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n369), .A2(G200), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n366), .A2(G190), .A3(new_n367), .A4(new_n368), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n386), .A2(new_n391), .A3(new_n387), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n369), .A2(G200), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT10), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n384), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G190), .B1(new_n333), .B2(new_n334), .ZN(new_n397));
  OAI21_X1  g0197(.A(G200), .B1(new_n327), .B2(new_n329), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n352), .A3(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n354), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT76), .ZN(new_n401));
  XOR2_X1   g0201(.A(KEYINPUT8), .B(G58), .Z(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n403));
  XOR2_X1   g0203(.A(KEYINPUT15), .B(G87), .Z(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n373), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n268), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(KEYINPUT71), .A3(new_n268), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n347), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n350), .A2(new_n412), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n285), .A2(G232), .A3(new_n314), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(new_n285), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n323), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n293), .A2(G244), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n367), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n306), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n422), .A2(G179), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n415), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n409), .A2(new_n410), .B1(new_n412), .B2(new_n347), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n422), .A2(new_n296), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(G200), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n414), .A4(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n312), .A2(new_n400), .A3(new_n401), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n304), .A2(new_n307), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n308), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(new_n430), .A3(new_n303), .A4(new_n300), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n354), .A2(new_n396), .A3(new_n399), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT76), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n230), .B(G87), .C1(new_n318), .C2(new_n319), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT22), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n339), .A2(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n230), .A2(G107), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT23), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT24), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n441), .A2(KEYINPUT24), .A3(new_n442), .A4(new_n444), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n268), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n273), .A2(G33), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n280), .A2(new_n274), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G107), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n274), .A2(G107), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT25), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n449), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(G257), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n456));
  OAI211_X1 g0256(.A(G250), .B(new_n314), .C1(new_n318), .C2(new_n319), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G294), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n323), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  INV_X1    g0262(.A(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(new_n291), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(G264), .A3(new_n284), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n460), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(G190), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(KEYINPUT79), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n467), .A2(new_n474), .A3(G264), .A4(new_n284), .ZN(new_n475));
  AOI221_X4 g0275(.A(KEYINPUT80), .B1(new_n459), .B2(new_n323), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT80), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n475), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n460), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n469), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G200), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n455), .B1(new_n472), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G244), .B(new_n314), .C1(new_n318), .C2(new_n319), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n314), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n323), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n467), .A2(G257), .A3(new_n284), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n469), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n255), .A2(new_n256), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G107), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT77), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G97), .A2(G107), .ZN(new_n501));
  NAND2_X1  g0301(.A1(KEYINPUT6), .A2(G107), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n206), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n501), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n498), .B(new_n499), .C1(new_n504), .C2(new_n205), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n230), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n263), .A2(new_n412), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n497), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n510), .A2(new_n268), .B1(new_n511), .B2(new_n275), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n451), .A2(G97), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n491), .A2(G190), .A3(new_n469), .A4(new_n493), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n495), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n223), .A2(new_n314), .ZN(new_n516));
  INV_X1    g0316(.A(G244), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G1698), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n516), .B(new_n518), .C1(new_n318), .C2(new_n319), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n323), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n462), .A2(G274), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n284), .B(G250), .C1(G1), .C2(new_n461), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n230), .B1(new_n321), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G87), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n205), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n230), .B(G68), .C1(new_n318), .C2(new_n319), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n230), .A2(G33), .A3(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n527), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n268), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n451), .A2(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n347), .A2(new_n405), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n522), .A2(G190), .A3(new_n523), .A4(new_n524), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n526), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n451), .A2(new_n404), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n542), .A3(new_n538), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n522), .A2(new_n382), .A3(new_n523), .A4(new_n524), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n284), .B1(new_n519), .B2(new_n520), .ZN(new_n545));
  INV_X1    g0345(.A(new_n524), .ZN(new_n546));
  INV_X1    g0346(.A(new_n523), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n543), .B(new_n544), .C1(G169), .C2(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n494), .A2(new_n306), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n275), .A2(new_n511), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n418), .B1(new_n255), .B2(new_n256), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n553), .A2(new_n506), .A3(new_n508), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n513), .C1(new_n554), .C2(new_n280), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n491), .A2(new_n382), .A3(new_n469), .A4(new_n493), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n515), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n483), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(new_n314), .C1(new_n318), .C2(new_n319), .ZN(new_n561));
  OAI211_X1 g0361(.A(G264), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n251), .A2(G303), .A3(new_n252), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n323), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n467), .A2(G270), .A3(new_n284), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n469), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G169), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n267), .A2(new_n229), .B1(G20), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(G33), .B2(G283), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n338), .A2(G97), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT78), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT78), .B1(new_n571), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT20), .B(new_n570), .C1(new_n573), .C2(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n347), .A2(G116), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n280), .A2(G116), .A3(new_n450), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n346), .A3(new_n345), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n560), .B1(new_n568), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n581), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n571), .A2(new_n572), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT20), .B1(new_n589), .B2(new_n570), .ZN(new_n590));
  INV_X1    g0390(.A(new_n578), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n584), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(KEYINPUT21), .A3(G169), .A4(new_n567), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n567), .A2(G200), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n565), .A2(new_n566), .A3(G190), .A4(new_n469), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n582), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n567), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n592), .A2(G179), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n583), .A2(new_n593), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(G179), .B(new_n469), .C1(new_n476), .C2(new_n479), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n471), .A2(G169), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n599), .B1(new_n455), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n439), .A2(new_n559), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g0404(.A(new_n604), .B(KEYINPUT81), .Z(G372));
  INV_X1    g0405(.A(new_n384), .ZN(new_n606));
  INV_X1    g0406(.A(new_n399), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n354), .B2(new_n425), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n300), .A2(new_n303), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n432), .A2(KEYINPUT83), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT83), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n304), .A2(new_n612), .A3(new_n307), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n304), .A2(new_n612), .A3(new_n307), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n304), .B2(new_n307), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n433), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n608), .A2(new_n610), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n392), .A2(new_n395), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n606), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n549), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n541), .A2(new_n549), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n557), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n557), .B2(new_n623), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n602), .A2(KEYINPUT82), .A3(new_n455), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT82), .B1(new_n602), .B2(new_n455), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n583), .A2(new_n593), .A3(new_n598), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n482), .A2(new_n472), .ZN(new_n633));
  INV_X1    g0433(.A(new_n455), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n515), .A2(new_n550), .A3(new_n557), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n628), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n621), .B1(new_n439), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT84), .ZN(G369));
  INV_X1    g0440(.A(G13), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(G20), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OR3_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .A3(G1), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT27), .B1(new_n643), .B2(G1), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n582), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n631), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n599), .B2(new_n650), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  INV_X1    g0453(.A(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n602), .A2(new_n455), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n483), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n455), .A2(new_n648), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n659), .A2(new_n660), .B1(new_n658), .B2(new_n648), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n631), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n648), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n649), .B1(new_n629), .B2(new_n630), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n662), .A2(new_n667), .ZN(G399));
  NAND2_X1  g0468(.A1(new_n210), .A2(new_n463), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT87), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n669), .A2(KEYINPUT87), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n530), .A2(G116), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT86), .Z(new_n675));
  OR2_X1    g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n673), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n676), .A2(new_n273), .B1(new_n233), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT28), .Z(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n638), .A2(new_n680), .A3(new_n649), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n631), .B1(new_n602), .B2(new_n455), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n682), .A2(new_n483), .A3(new_n558), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT26), .B1(new_n684), .B2(new_n550), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n549), .B1(new_n685), .B2(new_n625), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n649), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n603), .A2(new_n635), .A3(new_n636), .A4(new_n649), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT31), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n478), .A2(new_n460), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT80), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n478), .A2(new_n477), .A3(new_n460), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n494), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n565), .A2(new_n566), .A3(G179), .A4(new_n469), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n525), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n697), .ZN(new_n698));
  AOI211_X1 g0498(.A(new_n468), .B(new_n492), .C1(new_n490), .C2(new_n323), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n697), .B(new_n699), .C1(new_n476), .C2(new_n479), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n480), .A2(new_n382), .A3(new_n494), .A4(new_n567), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n698), .B(new_n702), .C1(new_n703), .C2(new_n548), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n648), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n691), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n654), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n689), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n679), .B1(new_n710), .B2(new_n273), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT88), .Z(G364));
  AOI21_X1  g0512(.A(new_n229), .B1(G20), .B2(new_n306), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n230), .A2(new_n382), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n481), .A2(G190), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G322), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n296), .A2(new_n481), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT90), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G326), .ZN(new_n726));
  INV_X1    g0526(.A(G294), .ZN(new_n727));
  OAI21_X1  g0527(.A(G20), .B1(new_n716), .B2(G179), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n718), .B1(new_n730), .B2(KEYINPUT92), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n230), .A2(G179), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n481), .A2(G190), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G283), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n714), .A2(new_n734), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT91), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n738), .A2(KEYINPUT91), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(KEYINPUT33), .B(G317), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G190), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n733), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n743), .A2(new_n744), .B1(G329), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n719), .A2(new_n733), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n285), .B1(new_n750), .B2(G303), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n732), .A2(new_n737), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n714), .A2(new_n745), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n731), .B(new_n752), .C1(G311), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n285), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n754), .B2(G77), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n717), .A2(G58), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n736), .A2(G107), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n728), .A2(G97), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n743), .A2(G68), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n750), .A2(G87), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT32), .B1(new_n746), .B2(new_n261), .ZN(new_n764));
  OR3_X1    g0564(.A1(new_n746), .A2(KEYINPUT32), .A3(new_n261), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n725), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n761), .B(new_n766), .C1(G50), .C2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n713), .B1(new_n755), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n273), .B1(new_n642), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n673), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n713), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n210), .A2(G355), .A3(new_n285), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G116), .B2(new_n210), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT89), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n210), .A2(new_n756), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n249), .B2(new_n461), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n461), .B2(new_n234), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n776), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n769), .A2(new_n772), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n653), .B2(new_n775), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n655), .A2(new_n772), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n653), .A2(new_n654), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G396));
  INV_X1    g0590(.A(new_n708), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT82), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n657), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n602), .A2(new_n455), .A3(KEYINPUT82), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n793), .A2(new_n663), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n686), .B1(new_n795), .B2(new_n559), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n648), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n415), .A2(new_n648), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n425), .A2(new_n429), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(KEYINPUT93), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT93), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n425), .A2(new_n429), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n425), .A2(new_n649), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n796), .A2(new_n648), .A3(new_n803), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n791), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n808), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n810), .B(new_n708), .C1(new_n797), .C2(new_n806), .ZN(new_n811));
  INV_X1    g0611(.A(new_n772), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n735), .A2(new_n529), .ZN(new_n814));
  INV_X1    g0614(.A(new_n717), .ZN(new_n815));
  INV_X1    g0615(.A(G303), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n756), .B1(new_n727), .B2(new_n815), .C1(new_n725), .C2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n814), .B(new_n817), .C1(G107), .C2(new_n750), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n747), .A2(G311), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n743), .A2(G283), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n754), .A2(G116), .B1(G97), .B2(new_n728), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G137), .A2(new_n767), .B1(new_n743), .B2(G150), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n261), .B2(new_n753), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G143), .B2(new_n717), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  NAND2_X1  g0626(.A1(new_n728), .A2(G58), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n736), .A2(G68), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n285), .B1(new_n746), .B2(new_n830), .C1(new_n202), .C2(new_n749), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n822), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n713), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n804), .B1(new_n800), .B2(new_n802), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n812), .B1(new_n834), .B2(new_n773), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n713), .A2(new_n773), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n833), .B(new_n835), .C1(G77), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n813), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT94), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n839), .B(new_n840), .ZN(G384));
  NAND2_X1  g0641(.A1(new_n503), .A2(new_n505), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n569), .B1(new_n842), .B2(KEYINPUT35), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n232), .C1(KEYINPUT35), .C2(new_n842), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  OAI21_X1  g0645(.A(G77), .B1(new_n258), .B2(new_n222), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n846), .A2(new_n233), .B1(G50), .B2(new_n222), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(G1), .A3(new_n641), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT95), .Z(new_n850));
  INV_X1    g0650(.A(KEYINPUT100), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n707), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n704), .A2(KEYINPUT100), .A3(KEYINPUT31), .A4(new_n648), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n706), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n439), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n646), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n311), .A2(new_n304), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n302), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(new_n298), .B1(new_n304), .B2(new_n857), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(new_n861), .A3(new_n432), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n282), .A2(new_n646), .B1(new_n302), .B2(new_n297), .ZN(new_n863));
  INV_X1    g0663(.A(new_n432), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n858), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n611), .B2(new_n613), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT99), .B(new_n862), .C1(new_n868), .C2(new_n861), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT99), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n615), .A2(new_n616), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n870), .B(KEYINPUT37), .C1(new_n871), .C2(new_n863), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n304), .A2(new_n857), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n609), .B1(new_n617), .B2(new_n614), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n869), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT101), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n834), .B1(new_n706), .B2(new_n854), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT97), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n354), .B2(new_n649), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n337), .A2(KEYINPUT97), .A3(new_n353), .A4(new_n648), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n354), .B(new_n399), .C1(new_n352), .C2(new_n649), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n878), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT40), .B1(new_n877), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n858), .B2(new_n866), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n858), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n878), .A2(new_n890), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n892), .A2(new_n879), .A3(new_n885), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n856), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n654), .B1(new_n887), .B2(new_n895), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n439), .A2(G330), .A3(new_n855), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n425), .A2(new_n648), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT96), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n885), .B1(new_n808), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n867), .A2(new_n888), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n617), .A2(new_n614), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n903), .A2(new_n904), .B1(new_n905), .B2(new_n857), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT98), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(KEYINPUT39), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n354), .A2(new_n648), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n909), .B(new_n910), .C1(new_n877), .C2(KEYINPUT39), .ZN(new_n911));
  OAI221_X1 g0711(.A(KEYINPUT98), .B1(new_n905), .B2(new_n857), .C1(new_n903), .C2(new_n904), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n900), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n621), .B1(new_n689), .B2(new_n439), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n642), .A2(new_n273), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n850), .B1(new_n916), .B2(new_n917), .ZN(G367));
  OR2_X1    g0718(.A1(new_n649), .A2(new_n539), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n550), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT102), .Z(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n549), .B2(new_n919), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT103), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n684), .A2(new_n648), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n555), .A2(new_n648), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n515), .A2(new_n557), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT105), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT105), .B1(new_n927), .B2(new_n929), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(new_n665), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  INV_X1    g0735(.A(new_n933), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n658), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n648), .B1(new_n937), .B2(new_n557), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n935), .A2(KEYINPUT106), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT106), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n934), .B(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n942), .B2(new_n938), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n926), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n940), .A2(new_n943), .A3(new_n926), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n662), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(new_n933), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n933), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n946), .A2(new_n951), .A3(new_n947), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n673), .B(KEYINPUT41), .Z(new_n953));
  INV_X1    g0753(.A(KEYINPUT107), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n661), .B1(new_n663), .B2(new_n648), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n665), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n656), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n710), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n667), .A2(new_n933), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT44), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n667), .A2(new_n933), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n961), .A2(new_n949), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n949), .B1(new_n961), .B2(new_n963), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n955), .B(new_n959), .C1(new_n967), .C2(new_n954), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n953), .B1(new_n968), .B2(new_n709), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n950), .B(new_n952), .C1(new_n969), .C2(new_n771), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n750), .A2(G116), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT46), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n285), .B1(new_n736), .B2(G97), .ZN(new_n973));
  INV_X1    g0773(.A(G311), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n725), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G303), .B2(new_n717), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n743), .A2(G294), .B1(G317), .B2(new_n747), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n754), .A2(G283), .B1(G107), .B2(new_n728), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT108), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n743), .A2(G159), .B1(G50), .B2(new_n754), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n756), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n750), .A2(G58), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n747), .A2(G137), .B1(new_n728), .B2(G68), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n735), .A2(new_n412), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n767), .B2(G143), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(G150), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n815), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n980), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT110), .Z(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n713), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n923), .A2(new_n775), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n776), .B1(new_n210), .B2(new_n405), .C1(new_n780), .C2(new_n242), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n995), .A2(new_n772), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n970), .A2(new_n998), .ZN(G387));
  AOI22_X1  g0799(.A1(G322), .A2(new_n767), .B1(new_n743), .B2(G311), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n816), .B2(new_n753), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G317), .B2(new_n717), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT48), .Z(new_n1003));
  INV_X1    g0803(.A(G283), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n729), .C1(new_n727), .C2(new_n749), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT49), .Z(new_n1006));
  OAI22_X1  g0806(.A1(new_n735), .A2(new_n569), .B1(new_n746), .B2(new_n726), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1006), .A2(new_n285), .A3(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n767), .A2(G159), .B1(G97), .B2(new_n736), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n272), .B2(new_n742), .C1(new_n405), .C2(new_n729), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n750), .A2(G77), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n222), .B2(new_n753), .C1(new_n990), .C2(new_n746), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n815), .A2(new_n202), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1010), .A2(new_n756), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n713), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n661), .A2(new_n775), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n675), .A2(new_n210), .A3(new_n285), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(G107), .B2(new_n210), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT111), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n272), .A2(G50), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1021));
  AOI21_X1  g0821(.A(G45), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n222), .B2(new_n412), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n781), .B1(new_n1023), .B2(new_n675), .C1(new_n461), .C2(new_n239), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n812), .B1(new_n1025), .B2(new_n776), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT113), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1015), .A2(new_n1016), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n959), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n677), .B1(new_n958), .B2(new_n710), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1028), .B(new_n1031), .C1(new_n770), .C2(new_n958), .ZN(G393));
  INV_X1    g0832(.A(new_n966), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n964), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT114), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(KEYINPUT114), .A3(new_n964), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n771), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n814), .B1(G143), .B2(new_n747), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n285), .C1(new_n222), .C2(new_n749), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT115), .Z(new_n1041));
  NAND2_X1  g0841(.A1(new_n728), .A2(G77), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n725), .A2(new_n990), .B1(new_n261), .B2(new_n815), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT51), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n742), .A2(new_n202), .B1(new_n272), .B2(new_n753), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT116), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n767), .A2(G317), .B1(G311), .B2(new_n717), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT52), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n759), .B1(new_n1004), .B2(new_n749), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n756), .B1(new_n729), .B2(new_n569), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n747), .A2(G322), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n727), .C2(new_n753), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n742), .A2(new_n816), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1047), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n713), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n933), .A2(new_n775), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n776), .B1(new_n511), .B2(new_n210), .C1(new_n780), .C2(new_n246), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n772), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1038), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1034), .A2(new_n1029), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n968), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1063), .B2(new_n673), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  INV_X1    g0865(.A(new_n910), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n903), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n872), .B1(new_n874), .B2(new_n873), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n611), .A2(new_n613), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n861), .B1(new_n1069), .B2(new_n860), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT37), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n870), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n876), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT39), .B1(new_n1073), .B2(new_n891), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT39), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n867), .A2(new_n888), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1067), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n902), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n687), .B2(new_n803), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1073), .A2(new_n891), .B1(new_n1079), .B2(new_n885), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1066), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n690), .A2(KEYINPUT31), .B1(new_n648), .B2(new_n704), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n707), .ZN(new_n1083));
  OAI211_X1 g0883(.A(G330), .B(new_n806), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n885), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n654), .B(new_n834), .C1(new_n706), .C2(new_n854), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1088), .B2(KEYINPUT117), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1077), .A2(new_n1081), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n909), .B1(new_n877), .B2(KEYINPUT39), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1091), .A2(new_n1067), .B1(new_n1066), .B2(new_n1080), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n855), .A2(G330), .A3(new_n806), .A4(new_n885), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(KEYINPUT117), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT119), .B1(new_n1096), .B2(new_n770), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(KEYINPUT117), .A3(new_n1094), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT119), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n771), .A4(new_n1090), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n796), .A2(KEYINPUT29), .A3(new_n648), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n628), .B1(new_n637), .B2(new_n682), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n680), .B1(new_n1104), .B2(new_n649), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n439), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n621), .ZN(new_n1107));
  AND4_X1   g0907(.A1(KEYINPUT118), .A2(new_n1106), .A3(new_n899), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT118), .B1(new_n915), .B2(new_n899), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1093), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n808), .A2(new_n902), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n708), .A2(new_n806), .A3(new_n885), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1079), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n1087), .C2(new_n885), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1099), .A2(new_n1090), .A3(new_n1110), .A4(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1106), .A2(new_n899), .A3(new_n1107), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n915), .A2(KEYINPUT118), .A3(new_n899), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1119), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1096), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1120), .A2(new_n1126), .A3(new_n673), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT120), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n749), .A2(KEYINPUT53), .A3(new_n990), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n285), .B1(new_n729), .B2(new_n261), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(new_n767), .C2(G128), .ZN(new_n1131));
  OAI21_X1  g0931(.A(KEYINPUT53), .B1(new_n749), .B2(new_n990), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n202), .B2(new_n735), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT54), .B(G143), .Z(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n753), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1133), .B(new_n1136), .C1(new_n743), .C2(G137), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n747), .A2(G125), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1131), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G132), .B2(new_n717), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n717), .A2(G116), .B1(G77), .B2(new_n728), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n754), .A2(G97), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1141), .A2(new_n756), .A3(new_n763), .A4(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n828), .B1(new_n742), .B2(new_n418), .C1(new_n1004), .C2(new_n725), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G294), .C2(new_n747), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n713), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n772), .C1(new_n402), .C2(new_n837), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1091), .A2(new_n773), .B1(new_n1128), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1128), .B2(new_n1147), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1102), .A2(new_n1127), .A3(new_n1149), .ZN(G378));
  OAI21_X1  g0950(.A(new_n1110), .B1(new_n1096), .B2(new_n1125), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n913), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n619), .A2(new_n606), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n381), .A2(new_n857), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n396), .A2(new_n1154), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n897), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT121), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT121), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n654), .B(new_n1168), .C1(new_n887), .C2(new_n895), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1152), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1168), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n897), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1172), .B(new_n913), .C1(new_n897), .C2(new_n1163), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1151), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT57), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1151), .A2(new_n1170), .A3(new_n1173), .A4(KEYINPUT57), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n673), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1170), .A2(new_n1173), .A3(new_n771), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n725), .A2(new_n569), .B1(new_n418), .B2(new_n815), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n285), .B(new_n1180), .C1(new_n404), .C2(new_n754), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1011), .B1(new_n258), .B2(new_n735), .C1(new_n1004), .C2(new_n746), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G41), .B(new_n1182), .C1(G68), .C2(new_n728), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(new_n511), .C2(new_n742), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT58), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n202), .B1(new_n318), .B2(G41), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n767), .A2(G125), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n743), .A2(G132), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n750), .A2(new_n1134), .B1(new_n728), .B2(G150), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G128), .A2(new_n717), .B1(new_n754), .B2(G137), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT59), .Z(new_n1192));
  OAI21_X1  g0992(.A(new_n463), .B1(new_n735), .B2(new_n261), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G124), .B2(new_n747), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n338), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1185), .A2(new_n1186), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n812), .B1(new_n1196), .B2(new_n713), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(G50), .B2(new_n837), .C1(new_n1171), .C2(new_n774), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1179), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1178), .A2(new_n1200), .ZN(G375));
  AOI21_X1  g1001(.A(new_n770), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1085), .A2(new_n773), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n836), .A2(new_n222), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n725), .A2(new_n830), .B1(new_n258), .B2(new_n735), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G50), .B2(new_n728), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n285), .B1(new_n742), .B2(new_n1135), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G137), .B2(new_n717), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G159), .A2(new_n750), .B1(new_n747), .B2(G128), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G150), .B2(new_n754), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n987), .B1(new_n767), .B2(G294), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n511), .B2(new_n749), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n746), .A2(new_n816), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n756), .B1(new_n1004), .B2(new_n815), .C1(new_n742), .C2(new_n569), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n405), .A2(new_n729), .B1(new_n418), .B2(new_n753), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n713), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1203), .A2(new_n772), .A3(new_n1204), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT122), .B1(new_n1202), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n885), .B1(new_n879), .B2(G330), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1222), .A2(new_n1086), .A3(new_n1079), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1113), .B1(new_n1093), .B2(new_n1111), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n771), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT122), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1226), .A3(new_n1219), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1222), .A2(new_n1086), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1224), .B1(new_n1230), .B2(new_n1117), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n953), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1125), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(new_n1234), .ZN(G381));
  NOR2_X1   g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1064), .A2(new_n970), .A3(new_n998), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G381), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT123), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1236), .A2(new_n1238), .A3(new_n1240), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n647), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(G213), .A3(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1044(.A(KEYINPUT126), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n647), .A2(G213), .A3(G2897), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1229), .A2(new_n1231), .A3(KEYINPUT60), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n673), .A3(new_n1125), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT60), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1228), .B(G384), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1255), .A2(new_n673), .A3(new_n1125), .A4(new_n1249), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G384), .B1(new_n1256), .B2(new_n1228), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1248), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1228), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(KEYINPUT125), .A3(new_n1252), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1247), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1252), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1247), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1245), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1253), .A2(new_n1257), .A3(new_n1248), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT125), .B1(new_n1261), .B2(new_n1252), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1246), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(KEYINPUT126), .A3(new_n1265), .ZN(new_n1271));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1151), .A2(new_n1170), .A3(new_n1173), .A4(new_n1233), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1200), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n647), .A2(G213), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n677), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1199), .B1(new_n1276), .B2(new_n1177), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1274), .B(new_n1275), .C1(new_n1277), .C2(new_n1272), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1267), .A2(new_n1271), .A3(new_n1278), .ZN(new_n1279));
  XOR2_X1   g1079(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1280));
  NAND3_X1  g1080(.A1(new_n1273), .A2(new_n1179), .A3(new_n1198), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1275), .B1(new_n1281), .B2(G378), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(G375), .B2(G378), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT62), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1272), .B1(new_n1178), .B2(new_n1200), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NOR4_X1   g1088(.A1(new_n1287), .A2(new_n1284), .A3(new_n1288), .A4(new_n1282), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1279), .B(new_n1280), .C1(new_n1286), .C2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(G393), .B(new_n789), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1237), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1064), .B1(new_n970), .B2(new_n998), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(G390), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1291), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1237), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1290), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT63), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(new_n1298), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1283), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1279), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(G405));
  OR3_X1    g1105(.A1(new_n1236), .A2(new_n1287), .A3(new_n1284), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1264), .B1(new_n1236), .B2(new_n1287), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1306), .A2(new_n1298), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1298), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(G402));
endmodule


