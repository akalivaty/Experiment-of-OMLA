//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n196), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n196), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n198), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n200), .A2(new_n202), .A3(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n208), .A2(new_n197), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT65), .A2(G134), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(KEYINPUT11), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT65), .A2(G134), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(G134), .B2(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n220), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G137), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n211), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT64), .B(G143), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n206), .B1(new_n229), .B2(G146), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n208), .A2(new_n197), .A3(new_n231), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n214), .A2(G137), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT65), .A2(G134), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n236), .A2(new_n237), .A3(new_n217), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n213), .A2(new_n215), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n238), .A2(G131), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n222), .B1(new_n216), .B2(new_n221), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n234), .B(new_n235), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n243));
  INV_X1    g057(.A(new_n197), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n229), .B2(G146), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n230), .A2(new_n233), .B1(new_n245), .B2(new_n231), .ZN(new_n246));
  OAI21_X1  g060(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n223), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n228), .B1(new_n243), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(KEYINPUT67), .A2(G119), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT67), .A2(G119), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(G116), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT2), .A2(G113), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT2), .A2(G113), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n254), .A2(new_n262), .A3(new_n263), .A4(new_n256), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n194), .B1(new_n251), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n223), .B(new_n226), .C1(new_n207), .C2(new_n210), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n249), .B1(new_n246), .B2(new_n248), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT30), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n265), .A2(new_n267), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n242), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n271), .A2(KEYINPUT70), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT70), .B1(new_n271), .B2(new_n281), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  XOR2_X1   g099(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n286));
  OAI211_X1 g100(.A(new_n270), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n276), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n268), .A2(new_n269), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n278), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n194), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n271), .A2(new_n281), .A3(new_n284), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(KEYINPUT32), .B(new_n187), .C1(new_n285), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n287), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n243), .A2(new_n250), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n270), .B1(new_n298), .B2(new_n272), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT28), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n292), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n194), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n289), .A2(new_n292), .A3(new_n194), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n275), .A2(new_n280), .B1(new_n251), .B2(new_n270), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n302), .B1(new_n307), .B2(new_n193), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G472), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n296), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n312));
  INV_X1    g126(.A(new_n187), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n293), .A2(new_n294), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n271), .A2(new_n281), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n271), .A2(new_n281), .A3(KEYINPUT70), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(KEYINPUT31), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n313), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n321));
  OAI21_X1  g135(.A(new_n312), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n187), .B1(new_n285), .B2(new_n295), .ZN(new_n323));
  INV_X1    g137(.A(new_n321), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(KEYINPUT73), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n311), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n330), .A3(KEYINPUT16), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n329), .A2(KEYINPUT16), .A3(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G146), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G146), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G110), .ZN(new_n337));
  AND2_X1   g151(.A1(KEYINPUT67), .A2(G119), .ZN(new_n338));
  NOR2_X1   g152(.A1(KEYINPUT67), .A2(G119), .ZN(new_n339));
  OAI21_X1  g153(.A(G128), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(G119), .A2(G128), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(KEYINPUT23), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n195), .B1(new_n338), .B2(new_n339), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n337), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n252), .A2(new_n253), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n341), .B1(new_n348), .B2(G128), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT24), .B(G110), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OR3_X1    g165(.A1(new_n336), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n343), .A2(new_n337), .A3(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n328), .A2(new_n330), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n196), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n333), .A2(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n355), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n352), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G137), .ZN(new_n363));
  INV_X1    g177(.A(G221), .ZN(new_n364));
  INV_X1    g178(.A(G234), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n364), .A2(new_n365), .A3(G953), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n363), .B(new_n366), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n352), .B(new_n367), .C1(new_n360), .C2(new_n361), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n305), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n372), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n369), .A2(new_n305), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G217), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(G234), .B2(new_n305), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(G902), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n369), .A2(new_n370), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT77), .B1(new_n326), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n296), .A2(new_n310), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n320), .A2(new_n312), .A3(new_n321), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT73), .B1(new_n323), .B2(new_n324), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n390));
  INV_X1    g204(.A(new_n384), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT99), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT9), .B(G234), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n395), .A2(new_n378), .A3(G953), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT13), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n203), .A2(KEYINPUT96), .A3(new_n195), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT96), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n229), .B2(G128), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n195), .A2(G143), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT97), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT96), .B1(new_n203), .B2(new_n195), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n229), .A2(new_n400), .A3(G128), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(KEYINPUT13), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n255), .A2(KEYINPUT95), .A3(G122), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT95), .B1(new_n255), .B2(G122), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n255), .A2(G122), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(KEYINPUT80), .A2(G107), .ZN(new_n414));
  AND2_X1   g228(.A1(KEYINPUT80), .A2(G107), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n414), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n417), .A3(new_n412), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n408), .A2(G134), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n225), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n404), .B1(new_n399), .B2(new_n401), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n405), .A2(new_n406), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT98), .B1(new_n424), .B2(new_n404), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n420), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n411), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n412), .B(KEYINPUT14), .ZN(new_n429));
  OAI21_X1  g243(.A(G107), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n418), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n422), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n424), .A2(KEYINPUT98), .A3(new_n404), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n225), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n426), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n397), .B1(new_n427), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n432), .A2(new_n225), .A3(new_n433), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n225), .B1(new_n432), .B2(new_n433), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n418), .B(new_n430), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n419), .A2(new_n426), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n396), .ZN(new_n441));
  AOI21_X1  g255(.A(G902), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI211_X1 g260(.A(G902), .B(new_n444), .C1(new_n436), .C2(new_n441), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n394), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n427), .A2(new_n435), .A3(new_n397), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n396), .B1(new_n439), .B2(new_n440), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n305), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n444), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n442), .A2(new_n445), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT99), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(G104), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n188), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n462));
  INV_X1    g276(.A(G214), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n463), .A2(G237), .A3(G953), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n461), .B(new_n462), .C1(new_n203), .C2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n462), .A2(new_n461), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n465), .A2(G131), .A3(new_n467), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n357), .A2(new_n196), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n468), .A2(KEYINPUT18), .B1(new_n358), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n465), .A2(new_n467), .B1(KEYINPUT18), .B2(G131), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n461), .ZN(new_n476));
  INV_X1    g290(.A(new_n464), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n229), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n222), .B1(new_n478), .B2(new_n466), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n465), .A2(new_n467), .A3(G131), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n468), .A2(KEYINPUT17), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n336), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n460), .B1(new_n475), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n469), .A2(new_n358), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n478), .A2(new_n466), .B1(new_n487), .B2(new_n222), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n471), .A2(new_n472), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G131), .B1(new_n465), .B2(new_n467), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n468), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT19), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n357), .B(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n333), .B1(new_n496), .B2(G146), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n460), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n456), .B1(new_n485), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n336), .B1(new_n481), .B2(new_n480), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n494), .B2(new_n480), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n459), .B1(new_n502), .B2(new_n492), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n479), .A2(new_n481), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n357), .B(KEYINPUT19), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n334), .B1(new_n505), .B2(new_n196), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n459), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n475), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(KEYINPUT91), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT92), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT20), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n485), .A2(new_n499), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT20), .B1(new_n512), .B2(KEYINPUT93), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(new_n516), .C1(KEYINPUT93), .C2(new_n512), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n502), .A2(new_n492), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n459), .A2(KEYINPUT94), .ZN(new_n519));
  AOI21_X1  g333(.A(G902), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n518), .B2(new_n519), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n514), .A2(new_n517), .B1(G475), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(KEYINPUT100), .A2(G952), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT100), .A2(G952), .ZN(new_n525));
  AOI21_X1  g339(.A(G953), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n365), .B2(new_n188), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT21), .B(G898), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n305), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n455), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT101), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n455), .A2(KEYINPUT101), .A3(new_n522), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n395), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n364), .B1(new_n538), .B2(new_n305), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT84), .ZN(new_n540));
  INV_X1    g354(.A(G101), .ZN(new_n541));
  INV_X1    g355(.A(G107), .ZN(new_n542));
  AND2_X1   g356(.A1(KEYINPUT79), .A2(G104), .ZN(new_n543));
  NOR2_X1   g357(.A1(KEYINPUT79), .A2(G104), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n545), .A2(KEYINPUT3), .B1(new_n417), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT79), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n458), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT79), .A2(G104), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(G107), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n541), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g366(.A1(KEYINPUT80), .A2(G107), .ZN(new_n553));
  NAND2_X1  g367(.A1(KEYINPUT80), .A2(G107), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(G107), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT3), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n541), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT4), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n551), .B(new_n555), .C1(new_n556), .C2(new_n557), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT4), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(G101), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n246), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT81), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(G101), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n547), .B2(new_n551), .ZN(new_n568));
  AOI21_X1  g382(.A(G146), .B1(new_n200), .B2(new_n202), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(new_n205), .ZN(new_n570));
  INV_X1    g384(.A(new_n233), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n235), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT81), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n562), .A2(G101), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n551), .A2(new_n541), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n547), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n577), .A3(KEYINPUT4), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n566), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n248), .ZN(new_n581));
  AOI21_X1  g395(.A(G104), .B1(new_n553), .B2(new_n554), .ZN(new_n582));
  OAI21_X1  g396(.A(G101), .B1(new_n582), .B2(new_n556), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT1), .B1(new_n229), .B2(G146), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n245), .B1(G128), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n577), .B(new_n583), .C1(new_n585), .C2(new_n210), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n558), .B2(new_n559), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n198), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n230), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n245), .A2(new_n209), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n586), .A2(new_n587), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n580), .A2(new_n581), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT83), .ZN(new_n597));
  INV_X1    g411(.A(new_n245), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT1), .ZN(new_n599));
  OAI21_X1  g413(.A(G128), .B1(new_n569), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n210), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n587), .B1(new_n601), .B2(new_n588), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n593), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n566), .B2(new_n579), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n597), .B1(new_n605), .B2(new_n581), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n574), .B1(new_n573), .B2(new_n578), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n594), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT83), .A3(new_n248), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n596), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n189), .A2(G227), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT78), .ZN(new_n613));
  XNOR2_X1  g427(.A(G110), .B(G140), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n540), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n597), .B(new_n581), .C1(new_n580), .C2(new_n594), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT83), .B1(new_n609), .B2(new_n248), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n595), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT84), .A3(new_n615), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n596), .A2(new_n615), .ZN(new_n622));
  INV_X1    g436(.A(new_n586), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n591), .A2(new_n592), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n589), .A2(new_n624), .ZN(new_n625));
  OAI221_X1 g439(.A(new_n248), .B1(KEYINPUT82), .B2(KEYINPUT12), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n623), .A2(new_n625), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n581), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n629));
  OAI21_X1  g443(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n617), .A2(new_n621), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G469), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n305), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n616), .B1(new_n630), .B2(new_n595), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n606), .A2(new_n610), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n635), .B1(new_n636), .B2(new_n622), .ZN(new_n637));
  OAI21_X1  g451(.A(G469), .B1(new_n637), .B2(G902), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n539), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT6), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n277), .A2(new_n568), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n254), .A2(KEYINPUT5), .A3(new_n256), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(G113), .C1(KEYINPUT5), .C2(new_n254), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n267), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n641), .A2(new_n578), .B1(new_n645), .B2(new_n589), .ZN(new_n646));
  XNOR2_X1  g460(.A(G110), .B(G122), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n641), .A2(new_n578), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n645), .A2(new_n589), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n647), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n651), .A2(new_n640), .A3(new_n652), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT85), .B1(new_n624), .B2(G125), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT85), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n211), .A2(new_n657), .A3(new_n329), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n656), .B(new_n658), .C1(new_n329), .C2(new_n246), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n189), .A2(G224), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT86), .Z(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n659), .B(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n654), .A2(new_n655), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(KEYINPUT7), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n647), .B(KEYINPUT8), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n644), .A2(new_n588), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n650), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n646), .A2(new_n647), .B1(new_n659), .B2(new_n665), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(G210), .B1(G237), .B2(G902), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT88), .Z(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n673), .B(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(G214), .B1(G237), .B2(G902), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n537), .A2(new_n639), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n393), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n541), .ZN(G3));
  INV_X1    g498(.A(new_n639), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n305), .B1(new_n285), .B2(new_n295), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n391), .A2(new_n687), .A3(new_n323), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n673), .A2(new_n676), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n664), .A2(new_n672), .A3(new_n675), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n690), .A2(new_n532), .A3(new_n679), .A4(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT33), .B1(new_n449), .B2(new_n450), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT33), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n436), .A2(new_n441), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(G478), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n443), .A2(new_n305), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n442), .B2(new_n443), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n692), .A2(new_n522), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n689), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G104), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G6));
  NAND2_X1  g518(.A1(new_n521), .A2(G475), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT20), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n706), .A2(new_n500), .A3(new_n509), .A4(new_n512), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(KEYINPUT103), .B2(new_n514), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n513), .A2(new_n709), .A3(KEYINPUT20), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n705), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n711), .A2(new_n455), .A3(new_n692), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n689), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT35), .B(G107), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G9));
  OR3_X1    g529(.A1(new_n362), .A2(KEYINPUT36), .A3(new_n368), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n362), .B1(KEYINPUT36), .B2(new_n368), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n381), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n380), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n687), .A2(new_n323), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n537), .A2(new_n639), .A3(new_n681), .A4(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT37), .B(G110), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G12));
  INV_X1    g539(.A(G900), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n528), .B1(new_n726), .B2(new_n530), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n711), .A2(new_n455), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n721), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n690), .A2(new_n679), .A3(new_n691), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n639), .A2(new_n728), .A3(new_n389), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G128), .ZN(G30));
  XOR2_X1   g547(.A(new_n678), .B(KEYINPUT38), .Z(new_n734));
  NOR2_X1   g548(.A1(new_n455), .A2(new_n522), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n679), .A2(new_n734), .A3(new_n729), .A4(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n727), .B(KEYINPUT39), .Z(new_n737));
  NAND2_X1  g551(.A1(new_n639), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n740));
  INV_X1    g554(.A(G472), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n298), .A2(new_n272), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n290), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n287), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n194), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n317), .A3(new_n318), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n741), .B1(new_n746), .B2(new_n305), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n320), .B2(KEYINPUT32), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n387), .B2(new_n388), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n736), .A2(new_n739), .A3(new_n740), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n203), .ZN(G45));
  NAND2_X1  g565(.A1(new_n514), .A2(new_n517), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n705), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n696), .A2(new_n698), .ZN(new_n754));
  INV_X1    g568(.A(new_n727), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n639), .A2(new_n389), .A3(new_n731), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G146), .ZN(G48));
  NOR2_X1   g573(.A1(new_n326), .A2(new_n384), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n632), .A2(new_n633), .A3(new_n305), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n633), .B1(new_n632), .B2(new_n305), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n761), .A2(new_n762), .A3(new_n539), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n763), .A3(new_n700), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT104), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT41), .B(G113), .Z(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G15));
  NAND3_X1  g581(.A1(new_n760), .A2(new_n763), .A3(new_n712), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G116), .ZN(G18));
  NOR2_X1   g583(.A1(new_n326), .A2(new_n729), .ZN(new_n770));
  INV_X1    g584(.A(new_n730), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n537), .A2(new_n770), .A3(new_n763), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G119), .ZN(G21));
  AND3_X1   g587(.A1(new_n380), .A2(KEYINPUT105), .A3(new_n383), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT105), .B1(new_n380), .B2(new_n383), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n292), .B1(new_n744), .B2(KEYINPUT28), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n294), .B1(new_n777), .B2(new_n193), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n187), .B1(new_n778), .B2(new_n285), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n687), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT106), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n384), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n380), .A2(KEYINPUT105), .A3(new_n383), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n319), .B(new_n294), .C1(new_n193), .C2(new_n777), .ZN(new_n787));
  AOI22_X1  g601(.A1(G472), .A2(new_n686), .B1(new_n787), .B2(new_n187), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n781), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n692), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n735), .A3(new_n791), .A4(new_n763), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G122), .ZN(G24));
  NOR2_X1   g607(.A1(new_n761), .A2(new_n762), .ZN(new_n794));
  INV_X1    g608(.A(new_n539), .ZN(new_n795));
  AOI21_X1  g609(.A(G902), .B1(new_n314), .B2(new_n319), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n779), .B(new_n721), .C1(new_n741), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n756), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n794), .A2(new_n795), .A3(new_n771), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G125), .ZN(G27));
  NAND2_X1  g614(.A1(new_n634), .A2(new_n638), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n678), .A2(new_n679), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n803), .A3(new_n795), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT107), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT107), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n639), .A2(new_n806), .A3(new_n803), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n805), .A2(new_n760), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n756), .A2(KEYINPUT42), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT32), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n323), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT108), .B1(new_n320), .B2(KEYINPUT32), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n386), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n785), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n756), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n805), .A3(new_n807), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n808), .A2(new_n809), .B1(new_n817), .B2(KEYINPUT42), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G131), .ZN(G33));
  NAND4_X1  g633(.A1(new_n805), .A2(new_n760), .A3(new_n728), .A4(new_n807), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G134), .ZN(G36));
  NOR2_X1   g635(.A1(new_n753), .A2(new_n699), .ZN(new_n822));
  NOR2_X1   g636(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n823));
  AND2_X1   g637(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n822), .B2(new_n824), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n729), .B1(new_n323), .B2(new_n687), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(KEYINPUT44), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n637), .A2(KEYINPUT45), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n637), .A2(KEYINPUT45), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(G469), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(G469), .A2(G902), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT46), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(KEYINPUT46), .A3(new_n834), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n634), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n839), .A2(new_n795), .A3(new_n737), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT44), .B1(new_n826), .B2(new_n827), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n802), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n830), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G137), .ZN(G39));
  NOR4_X1   g658(.A1(new_n389), .A2(new_n391), .A3(new_n756), .A4(new_n802), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n839), .A2(KEYINPUT47), .A3(new_n795), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT47), .B1(new_n839), .B2(new_n795), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G140), .ZN(G42));
  NOR3_X1   g663(.A1(new_n734), .A2(new_n539), .A3(new_n680), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n822), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n749), .A3(new_n776), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n794), .B(KEYINPUT111), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT49), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n853), .A2(KEYINPUT49), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n826), .A2(new_n528), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n790), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n846), .A2(new_n847), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n853), .A2(new_n795), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n803), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n794), .A2(new_n795), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n863), .A2(new_n679), .A3(new_n734), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT50), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n863), .A2(new_n802), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n857), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n797), .ZN(new_n869));
  INV_X1    g683(.A(new_n867), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n870), .A2(new_n384), .A3(new_n527), .A4(new_n749), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n753), .A2(new_n754), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n862), .A2(new_n866), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n862), .A2(new_n866), .A3(KEYINPUT51), .A4(new_n873), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n868), .A2(new_n815), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT48), .Z(new_n879));
  NAND4_X1  g693(.A1(new_n857), .A2(new_n771), .A3(new_n763), .A4(new_n790), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT119), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n526), .B(KEYINPUT118), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n522), .A2(new_n699), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n871), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n879), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n876), .A2(new_n877), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n760), .B(new_n763), .C1(new_n700), .C2(new_n712), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n723), .B(new_n887), .C1(new_n393), .C2(new_n682), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n681), .A2(new_n532), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n883), .A2(KEYINPUT112), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n452), .A2(new_n453), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n522), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n522), .B2(new_n699), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n688), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n890), .A2(new_n896), .A3(new_n639), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n792), .A2(new_n772), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n455), .A2(new_n730), .A3(new_n522), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n727), .B(KEYINPUT114), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n721), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n639), .A2(new_n749), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n758), .A2(new_n904), .A3(KEYINPUT52), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n799), .A2(new_n732), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n799), .A2(new_n732), .A3(new_n758), .A4(new_n904), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n805), .A2(new_n798), .A3(new_n807), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n711), .A2(new_n892), .A3(new_n727), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n639), .A3(new_n770), .A4(new_n803), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n820), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n900), .A2(new_n911), .A3(new_n818), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n910), .A2(KEYINPUT115), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n908), .A2(new_n921), .A3(new_n909), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n799), .A2(new_n732), .A3(KEYINPUT113), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT113), .B1(new_n799), .B2(new_n732), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n905), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n920), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n900), .A2(new_n818), .A3(new_n916), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT116), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n919), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n917), .A2(KEYINPUT116), .A3(new_n918), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n917), .A2(new_n918), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n920), .A2(new_n922), .A3(new_n925), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n820), .A2(new_n912), .A3(new_n915), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n935), .A2(new_n888), .A3(new_n899), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT53), .A4(new_n818), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n937), .A3(KEYINPUT117), .ZN(new_n938));
  INV_X1    g752(.A(new_n927), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT53), .A4(new_n934), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n886), .A2(new_n932), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(G952), .A2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n856), .B1(new_n945), .B2(new_n946), .ZN(G75));
  NAND4_X1  g761(.A1(new_n938), .A2(G902), .A3(new_n675), .A4(new_n941), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n654), .A2(new_n655), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n663), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n948), .B2(new_n949), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n189), .A2(G952), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G51));
  XOR2_X1   g770(.A(new_n834), .B(KEYINPUT57), .Z(new_n957));
  AND3_X1   g771(.A1(new_n938), .A2(KEYINPUT54), .A3(new_n941), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT54), .B1(new_n938), .B2(new_n941), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n632), .ZN(new_n961));
  OR3_X1    g775(.A1(new_n942), .A2(new_n305), .A3(new_n833), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n961), .B2(new_n962), .ZN(G54));
  AND2_X1   g777(.A1(KEYINPUT58), .A2(G475), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n938), .A2(G902), .A3(new_n941), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n500), .A2(new_n509), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT120), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n955), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n965), .A2(KEYINPUT120), .A3(new_n966), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G60));
  NAND2_X1  g785(.A1(new_n693), .A2(new_n695), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n932), .A2(new_n944), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n697), .B(KEYINPUT59), .Z(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n972), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n958), .B2(new_n959), .ZN(new_n977));
  INV_X1    g791(.A(new_n955), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n975), .A2(new_n979), .ZN(G63));
  NAND2_X1  g794(.A1(new_n369), .A2(new_n370), .ZN(new_n981));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT60), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n942), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n938), .A2(new_n719), .A3(new_n941), .A4(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n984), .A2(new_n978), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n984), .A2(KEYINPUT61), .A3(new_n978), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  XOR2_X1   g805(.A(new_n900), .B(KEYINPUT121), .Z(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n189), .ZN(new_n993));
  INV_X1    g807(.A(G224), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n529), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n950), .B1(G898), .B2(new_n189), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT122), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G69));
  NAND2_X1  g813(.A1(new_n278), .A2(new_n279), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n275), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT123), .Z(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(new_n505), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n923), .A2(new_n924), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n750), .A3(new_n758), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1004), .A2(KEYINPUT62), .A3(new_n750), .A4(new_n758), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n843), .A2(new_n848), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n385), .A2(new_n392), .ZN(new_n1011));
  INV_X1    g825(.A(new_n738), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1011), .A2(new_n1012), .A3(new_n803), .A4(new_n896), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT124), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(KEYINPUT125), .B(new_n1003), .C1(new_n1016), .C2(G953), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT125), .ZN(new_n1018));
  AOI21_X1  g832(.A(G953), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1003), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1003), .B1(G900), .B2(G953), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n840), .A2(new_n785), .A3(new_n814), .A4(new_n901), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n820), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1010), .A2(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1004), .A2(new_n758), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1025), .A2(new_n818), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1022), .B1(new_n1027), .B2(G953), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1017), .A2(new_n1021), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(G227), .ZN(new_n1030));
  OAI21_X1  g844(.A(G953), .B1(new_n1030), .B2(new_n726), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT126), .Z(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1017), .A2(new_n1021), .A3(new_n1032), .A4(new_n1028), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(G72));
  INV_X1    g850(.A(new_n307), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1037), .A2(new_n193), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n307), .A2(new_n194), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1041), .B(KEYINPUT63), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n955), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1027), .ZN(new_n1044));
  AOI22_X1  g858(.A1(new_n1044), .A2(new_n1038), .B1(new_n1016), .B2(new_n1039), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1043), .B1(new_n1045), .B2(new_n992), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n930), .A2(new_n931), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n282), .A2(new_n283), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1037), .A2(new_n194), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1050), .B(KEYINPUT127), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n1046), .A2(new_n1052), .ZN(G57));
endmodule


