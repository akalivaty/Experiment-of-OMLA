//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1226, new_n1227,
    new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n469), .A2(new_n472), .A3(new_n464), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n478), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n479), .B2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n471), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n473), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n476), .B1(new_n480), .B2(new_n486), .ZN(G160));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n469), .A2(new_n472), .A3(G2105), .A4(new_n473), .ZN(new_n492));
  OAI221_X1 g067(.A(new_n489), .B1(new_n474), .B2(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  AND2_X1   g069(.A1(KEYINPUT4), .A2(G138), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n469), .A2(new_n472), .A3(G126), .A4(new_n473), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n464), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n464), .A2(G138), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT4), .B1(new_n478), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n498), .A2(new_n501), .A3(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n510), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G88), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n506), .B1(new_n516), .B2(new_n518), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n509), .A2(G62), .ZN(new_n523));
  AND2_X1   g098(.A1(G75), .A2(G543), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n515), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT72), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n519), .A2(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n521), .A2(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n507), .A2(new_n534), .A3(new_n508), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n533), .A2(G63), .A3(G651), .A4(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AND2_X1   g113(.A1(new_n512), .A2(new_n514), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n533), .A2(G64), .A3(new_n535), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT73), .B(G90), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT6), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n512), .B2(new_n514), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n509), .B(new_n543), .C1(new_n545), .C2(new_n517), .ZN(new_n546));
  OAI21_X1  g121(.A(G543), .B1(new_n545), .B2(new_n517), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n542), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n509), .B1(new_n545), .B2(new_n517), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n551), .A2(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n533), .A2(G56), .A3(new_n535), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n539), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n545), .C2(new_n517), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n552), .A2(KEYINPUT75), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n568), .B(new_n509), .C1(new_n545), .C2(new_n517), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(G91), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n509), .A2(G65), .ZN(new_n571));
  AND2_X1   g146(.A1(G78), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n566), .A2(new_n570), .A3(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n533), .A2(new_n535), .ZN(new_n576));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n511), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(G49), .B2(new_n521), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n567), .A2(G87), .A3(new_n569), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n567), .A2(G86), .A3(new_n569), .ZN(new_n582));
  INV_X1    g157(.A(new_n508), .ZN(new_n583));
  NOR2_X1   g158(.A1(KEYINPUT5), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n539), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n521), .B2(G48), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n582), .A2(new_n588), .ZN(G305));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n547), .B1(new_n552), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n533), .A2(G60), .A3(new_n535), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n539), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n599));
  NAND4_X1  g174(.A1(new_n567), .A2(G92), .A3(new_n569), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n510), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n521), .A2(G54), .B1(new_n603), .B2(G651), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n567), .A2(G92), .A3(new_n569), .ZN(new_n606));
  INV_X1    g181(.A(new_n599), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n558), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n617), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT77), .ZN(new_n621));
  MUX2_X1   g196(.A(new_n619), .B(new_n621), .S(G868), .Z(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n478), .A2(new_n466), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT78), .Z(new_n629));
  NOR2_X1   g204(.A1(new_n464), .A2(G111), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n468), .B1(new_n630), .B2(KEYINPUT79), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT79), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n492), .ZN(new_n636));
  INV_X1    g211(.A(new_n474), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(G135), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n629), .B(new_n639), .C1(new_n627), .C2(new_n626), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(G14), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  OR3_X1    g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  INV_X1    g238(.A(new_n657), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n658), .B(KEYINPUT17), .Z(new_n665));
  OAI211_X1 g240(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n657), .A3(new_n658), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n661), .A3(new_n664), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT84), .ZN(new_n674));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n681), .A2(new_n689), .A3(new_n684), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(KEYINPUT82), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n681), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G1981), .ZN(new_n698));
  INV_X1    g273(.A(G1981), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n691), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n698), .A2(G1986), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(G1986), .B1(new_n698), .B2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n674), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(new_n674), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n701), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1991), .B(G1996), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n704), .B2(new_n707), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT33), .B(G1976), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n716), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n713), .B(new_n718), .C1(new_n714), .C2(new_n712), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n712), .A2(G22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT87), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G303), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1971), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n717), .A2(new_n719), .A3(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G6), .B(G305), .S(G16), .Z(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT32), .B(G1981), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT88), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n712), .A2(G24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n596), .B2(new_n712), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1986), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G25), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT85), .Z(new_n737));
  AND2_X1   g312(.A1(new_n637), .A2(G131), .ZN(new_n738));
  INV_X1    g313(.A(G119), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n464), .A2(G107), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n492), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n743), .B2(new_n735), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT35), .B(G1991), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT86), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n744), .B(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n734), .B(new_n747), .C1(new_n728), .C2(new_n729), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n731), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT36), .ZN(new_n750));
  NOR2_X1   g325(.A1(G168), .A2(new_n712), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n712), .B2(G21), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT91), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n735), .A2(G32), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(new_n760), .B1(G105), .B2(new_n466), .ZN(new_n761));
  INV_X1    g336(.A(G129), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n492), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G141), .B2(new_n637), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n756), .B1(new_n764), .B2(new_n735), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT27), .B(G1996), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n752), .A2(new_n753), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n755), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT25), .ZN(new_n772));
  NAND2_X1  g347(.A1(G115), .A2(G2104), .ZN(new_n773));
  INV_X1    g348(.A(G127), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n483), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n772), .B1(G2105), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n637), .A2(G139), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n735), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n735), .B2(G33), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G2072), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(G2072), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G11), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT30), .B(G28), .Z(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n638), .B2(G29), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n783), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n735), .B1(KEYINPUT24), .B2(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(KEYINPUT24), .B2(G34), .ZN(new_n791));
  INV_X1    g366(.A(G160), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2084), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n712), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n712), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n793), .A2(new_n794), .B1(new_n796), .B2(G1961), .ZN(new_n797));
  NOR2_X1   g372(.A1(G27), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n770), .A2(new_n789), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n793), .A2(new_n794), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT93), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n796), .A2(G1961), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT92), .Z(new_n805));
  INV_X1    g380(.A(G2090), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G35), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G162), .B2(G29), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n805), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n803), .B(new_n811), .C1(new_n806), .C2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G16), .A2(G19), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n558), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT89), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1341), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n712), .A2(G20), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT23), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n614), .B2(new_n712), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1956), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n735), .A2(G26), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT28), .Z(new_n823));
  OR2_X1    g398(.A1(G104), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n825));
  INV_X1    g400(.A(G140), .ZN(new_n826));
  INV_X1    g401(.A(G128), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n825), .B1(new_n474), .B2(new_n826), .C1(new_n827), .C2(new_n492), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n637), .A2(G140), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n492), .A2(new_n827), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT90), .A4(new_n825), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n823), .B1(new_n834), .B2(G29), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2067), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n817), .A2(new_n821), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n712), .A2(G4), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n610), .B2(new_n712), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1348), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n813), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n750), .A2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n750), .A2(new_n841), .ZN(G150));
  NAND2_X1  g418(.A1(new_n610), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n519), .A2(G93), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT96), .B(G55), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n521), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n533), .A2(G67), .A3(new_n535), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n539), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n846), .B(new_n848), .C1(new_n851), .C2(KEYINPUT95), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(KEYINPUT95), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n619), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n851), .A2(KEYINPUT95), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n846), .A2(new_n848), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n856), .A2(new_n558), .A3(new_n857), .A4(new_n853), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n845), .B(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n861), .A2(new_n862), .A3(G860), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n856), .A2(new_n857), .A3(new_n853), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n863), .A2(new_n866), .ZN(G145));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n638), .B(new_n493), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n792), .ZN(new_n870));
  INV_X1    g445(.A(new_n764), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n830), .A2(G164), .A3(new_n833), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G164), .B1(new_n830), .B2(new_n833), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(new_n779), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n499), .A2(new_n500), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n503), .B1(new_n876), .B2(G2105), .ZN(new_n877));
  INV_X1    g452(.A(new_n498), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n834), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n778), .B1(new_n880), .B2(new_n872), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n871), .B1(new_n875), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(G106), .A2(G2105), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n884));
  INV_X1    g459(.A(G142), .ZN(new_n885));
  INV_X1    g460(.A(G130), .ZN(new_n886));
  OAI221_X1 g461(.A(new_n884), .B1(new_n474), .B2(new_n885), .C1(new_n886), .C2(new_n492), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n625), .ZN(new_n888));
  INV_X1    g463(.A(new_n743), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n779), .B1(new_n873), .B2(new_n874), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n880), .A2(new_n778), .A3(new_n872), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n764), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n882), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT98), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n882), .A2(new_n896), .A3(new_n893), .A4(new_n890), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n882), .A2(new_n893), .ZN(new_n900));
  INV_X1    g475(.A(new_n890), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g477(.A(KEYINPUT97), .B(new_n890), .C1(new_n882), .C2(new_n893), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n870), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n901), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n870), .A3(new_n894), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n868), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(KEYINPUT97), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n900), .A2(new_n899), .A3(new_n901), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(new_n895), .A3(new_n897), .A4(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n870), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT99), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g494(.A(G868), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n864), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n855), .A2(new_n858), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n621), .B(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n614), .A2(new_n608), .A3(new_n605), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n609), .A2(G299), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n926), .B2(KEYINPUT41), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(KEYINPUT41), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n924), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n934), .B2(new_n929), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n928), .B1(new_n935), .B2(new_n923), .ZN(new_n936));
  XNOR2_X1  g511(.A(G288), .B(G166), .ZN(new_n937));
  XNOR2_X1  g512(.A(G305), .B(new_n596), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n936), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n921), .B1(new_n944), .B2(new_n920), .ZN(G295));
  OAI21_X1  g520(.A(new_n921), .B1(new_n944), .B2(new_n920), .ZN(G331));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n947));
  NAND2_X1  g522(.A1(G171), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT102), .B1(new_n542), .B2(new_n549), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(G168), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(G301), .A2(KEYINPUT102), .A3(G286), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n859), .A3(KEYINPUT105), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n950), .A2(new_n855), .A3(new_n858), .A4(new_n951), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(new_n951), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n922), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT104), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n922), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n957), .A2(new_n927), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(KEYINPUT103), .A3(new_n954), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n952), .A2(new_n859), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n963), .B(new_n941), .C1(new_n935), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n908), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n941), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n939), .A2(KEYINPUT106), .A3(new_n940), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT100), .B1(new_n931), .B2(new_n933), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n966), .B(new_n964), .C1(new_n974), .C2(new_n930), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n975), .B2(new_n963), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n968), .A2(new_n908), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n967), .A2(new_n927), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT107), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n957), .A2(new_n960), .A3(new_n962), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n934), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n967), .A2(new_n984), .A3(new_n927), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n973), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n979), .A2(new_n988), .A3(KEYINPUT43), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT44), .B1(new_n978), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n979), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n969), .B2(new_n976), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(KEYINPUT44), .B2(new_n995), .ZN(G397));
  OR2_X1    g571(.A1(new_n834), .A2(G2067), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n834), .A2(G2067), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G164), .B2(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G160), .A2(G40), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT108), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(KEYINPUT108), .ZN(new_n1006));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n764), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1005), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n743), .B(new_n746), .Z(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1003), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1986), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n596), .B(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n1003), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G40), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n1017), .B(new_n476), .C1(new_n480), .C2(new_n486), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1384), .B1(new_n877), .B2(new_n878), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1022), .B(new_n1024), .C1(new_n1023), .C2(G288), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G288), .A2(new_n1023), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n1026), .B2(new_n1021), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n582), .A2(new_n699), .A3(new_n588), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n582), .A2(new_n588), .A3(KEYINPUT111), .A4(new_n699), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G86), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n588), .B1(new_n1034), .B2(new_n552), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G1981), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1031), .A2(new_n1032), .B1(G1981), .B2(new_n1035), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT112), .B1(new_n1041), .B2(KEYINPUT49), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1021), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1028), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1002), .A2(G2090), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT109), .B1(new_n1019), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n879), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1384), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n879), .A2(KEYINPUT45), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1001), .A2(new_n1018), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1971), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G303), .A2(G8), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT55), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1057), .A2(new_n1062), .A3(KEYINPUT110), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1065), .A2(G8), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1055), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT114), .B1(G164), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n879), .A2(new_n1075), .A3(new_n1055), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1018), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n1078));
  AOI21_X1  g653(.A(G2090), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1019), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1002), .B1(new_n1080), .B2(KEYINPUT50), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT115), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1071), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1067), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1060), .A2(new_n753), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1054), .A2(new_n1052), .A3(new_n1018), .A4(new_n1056), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(G2084), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1088), .A2(G8), .A3(G168), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1049), .A2(new_n1070), .A3(new_n1085), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT63), .B1(new_n1090), .B2(KEYINPUT116), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(new_n1048), .A3(new_n1022), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1028), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1093), .A2(new_n1085), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1070), .A4(new_n1089), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1089), .A2(KEYINPUT63), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1065), .A2(G8), .A3(new_n1069), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1067), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1099), .A2(new_n1049), .A3(new_n1101), .A4(new_n1070), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1049), .A2(new_n1070), .A3(new_n1085), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1086), .B(G168), .C1(new_n1087), .C2(G2084), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1109), .B2(new_n1084), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1088), .A2(G286), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1111), .A2(KEYINPUT51), .A3(G8), .A4(new_n1108), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT62), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1961), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1087), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1060), .B2(G2078), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1117), .A2(G2078), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1060), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(G301), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1105), .A2(new_n1106), .A3(new_n1114), .A4(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1049), .A2(new_n1122), .A3(new_n1070), .A4(new_n1085), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT125), .B1(new_n1124), .B2(new_n1113), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT62), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1093), .A2(new_n1023), .A3(new_n714), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1021), .B1(new_n1129), .B2(new_n1033), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1070), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1049), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1103), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n479), .A2(new_n464), .ZN(new_n1135));
  NOR4_X1   g710(.A1(new_n1135), .A2(new_n476), .A3(new_n1017), .A4(new_n1120), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1001), .A2(new_n1059), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1116), .A2(new_n1118), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(G171), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1122), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1095), .A2(new_n1140), .A3(new_n1126), .A4(new_n1070), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(G171), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1121), .A2(new_n1116), .A3(G301), .A4(new_n1118), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT54), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT124), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1104), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1144), .B(KEYINPUT123), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1140), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT117), .B(G1956), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT118), .B1(new_n1077), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1077), .A2(KEYINPUT118), .A3(new_n1153), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n1158));
  XNOR2_X1  g733(.A(G299), .B(KEYINPUT57), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT56), .B(G2072), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1001), .A2(new_n1059), .A3(new_n1018), .A4(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1077), .A2(KEYINPUT118), .A3(new_n1153), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1160), .B(new_n1162), .C1(new_n1164), .C2(new_n1154), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT119), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1162), .B1(new_n1164), .B2(new_n1154), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1159), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1020), .A2(G2067), .ZN(new_n1170));
  INV_X1    g745(.A(G1348), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1087), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n609), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n1168), .B2(new_n1159), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1165), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1165), .A2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1172), .A2(KEYINPUT60), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n610), .B1(new_n1172), .B2(KEYINPUT60), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n619), .A2(KEYINPUT121), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1001), .A2(new_n1059), .A3(new_n1007), .A4(new_n1018), .ZN(new_n1185));
  XOR2_X1   g760(.A(KEYINPUT58), .B(G1341), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n1020), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1188), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1190));
  OAI211_X1 g765(.A(KEYINPUT59), .B(new_n1184), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1172), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT59), .B1(new_n1197), .B2(new_n1184), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1183), .A2(new_n1193), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1180), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(KEYINPUT61), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1174), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1147), .A2(new_n1152), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1016), .B1(new_n1133), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n997), .A2(new_n764), .A3(new_n998), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT46), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1207));
  AOI22_X1  g782(.A1(new_n1205), .A2(new_n1003), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1208), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT47), .Z(new_n1210));
  OR3_X1    g785(.A1(new_n1010), .A2(new_n746), .A3(new_n889), .ZN(new_n1211));
  AOI211_X1 g786(.A(new_n1002), .B(new_n1001), .C1(new_n1211), .C2(new_n997), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1003), .A2(new_n1014), .A3(new_n596), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT48), .ZN(new_n1214));
  AOI211_X1 g789(.A(new_n1210), .B(new_n1212), .C1(new_n1012), .C2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1204), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g791(.A1(new_n462), .A2(G227), .ZN(new_n1218));
  OR2_X1    g792(.A1(new_n1218), .A2(KEYINPUT126), .ZN(new_n1219));
  AOI21_X1  g793(.A(G401), .B1(KEYINPUT126), .B2(new_n1218), .ZN(new_n1220));
  OAI211_X1 g794(.A(new_n1219), .B(new_n1220), .C1(new_n709), .C2(new_n710), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1221), .B1(new_n910), .B2(new_n917), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n1222), .A2(new_n994), .A3(KEYINPUT127), .ZN(new_n1223));
  AOI21_X1  g797(.A(KEYINPUT127), .B1(new_n1222), .B2(new_n994), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n1223), .A2(new_n1224), .ZN(G308));
  NAND2_X1  g799(.A1(new_n1222), .A2(new_n994), .ZN(new_n1226));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1227));
  NAND2_X1  g801(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n1222), .A2(new_n994), .A3(KEYINPUT127), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1229), .ZN(G225));
endmodule


