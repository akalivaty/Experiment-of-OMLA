//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT64), .Z(G173));
  XOR2_X1   g022(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(G234));
  NAND2_X1  g028(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT68), .B1(new_n476), .B2(new_n463), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  INV_X1    g054(.A(new_n470), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(G2105), .C1(new_n482), .C2(new_n474), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n463), .A2(new_n473), .B1(new_n477), .B2(new_n483), .ZN(G160));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n471), .A2(new_n485), .ZN(new_n486));
  AOI211_X1 g061(.A(KEYINPUT70), .B(new_n470), .C1(new_n468), .C2(KEYINPUT3), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT71), .Z(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G112), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n488), .A2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G136), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  AND2_X1   g073(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n463), .C1(new_n499), .C2(new_n470), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n504));
  NAND2_X1  g079(.A1(G126), .A2(G2105), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT4), .A2(G138), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n502), .B(new_n504), .C1(new_n471), .C2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT73), .B1(new_n513), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(new_n511), .A3(KEYINPUT5), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(new_n524), .B1(new_n522), .B2(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(G88), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n517), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n520), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT75), .Z(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n525), .A2(new_n517), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT76), .B(G89), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n535), .B1(new_n528), .B2(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n533), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n519), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT77), .ZN(new_n543));
  INV_X1    g118(.A(new_n537), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n525), .A2(G543), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT78), .B(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n544), .A2(G90), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n543), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n512), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n515), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n552));
  NOR3_X1   g127(.A1(new_n513), .A2(KEYINPUT73), .A3(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n519), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n558), .B1(new_n557), .B2(new_n556), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT80), .B(G81), .Z(new_n560));
  AOI22_X1  g135(.A1(new_n544), .A2(new_n560), .B1(new_n545), .B2(G43), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n545), .A2(new_n570), .A3(G53), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n528), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT81), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G91), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n576), .A2(new_n519), .B1(new_n537), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  OAI21_X1  g157(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n525), .A2(G49), .A3(G543), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n537), .ZN(G288));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  INV_X1    g162(.A(G73), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n554), .A2(new_n587), .B1(new_n588), .B2(new_n511), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n545), .B2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n544), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n544), .A2(G85), .B1(new_n545), .B2(G47), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n519), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n544), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n554), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n545), .B2(G54), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n596), .B1(new_n603), .B2(G868), .ZN(G321));
  MUX2_X1   g180(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g181(.A(G297), .B(KEYINPUT82), .ZN(G280));
  XNOR2_X1  g182(.A(KEYINPUT83), .B(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n603), .B1(G860), .B2(new_n608), .ZN(G148));
  NAND2_X1  g184(.A1(new_n603), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n489), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n463), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n495), .A2(KEYINPUT84), .A3(G135), .ZN(new_n617));
  AOI21_X1  g192(.A(KEYINPUT84), .B1(new_n495), .B2(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n614), .B1(new_n615), .B2(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2096), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2096), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n468), .A2(new_n475), .A3(new_n463), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2100), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(G156));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT85), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n631), .B(new_n637), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(G14), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n639), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NOR2_X1   g220(.A1(G2072), .A2(G2078), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n644), .B(new_n645), .C1(new_n442), .C2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(KEYINPUT86), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n442), .A2(new_n646), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n644), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(KEYINPUT17), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n651), .B(new_n652), .C1(new_n649), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n649), .A3(new_n644), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT88), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n662), .A2(new_n663), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n659), .B(new_n660), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n673), .B2(new_n664), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n668), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  INV_X1    g259(.A(G29), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n685), .A2(G35), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n497), .B2(G29), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT29), .ZN(new_n688));
  INV_X1    g263(.A(G2090), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G19), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n563), .B2(new_n691), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(G1341), .ZN(new_n694));
  NOR2_X1   g269(.A1(G4), .A2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT97), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n598), .A2(new_n602), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n691), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1348), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(G1341), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n691), .A2(G20), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT23), .Z(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G299), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT105), .B(G1956), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n690), .A2(new_n694), .A3(new_n701), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n685), .A2(G26), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n495), .A2(G140), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n489), .A2(G128), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT98), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT98), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n711), .A2(new_n712), .A3(new_n717), .A4(new_n714), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n710), .B1(new_n719), .B2(G29), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G2067), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n688), .B2(new_n689), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n708), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n685), .A2(G32), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n489), .A2(G129), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n495), .A2(G141), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n468), .A2(G105), .A3(new_n463), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT101), .Z(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT26), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n725), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n724), .B1(new_n733), .B2(new_n685), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT102), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(KEYINPUT102), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n685), .A2(G33), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT25), .Z(new_n741));
  AOI22_X1  g316(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n463), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n495), .B2(G139), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT99), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT100), .B(G2072), .Z(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G160), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n749), .A2(G29), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n746), .B2(new_n747), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n738), .A2(new_n748), .A3(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT103), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(KEYINPUT103), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n754), .A2(new_n755), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G11), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT30), .B(G28), .Z(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(G164), .A2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G27), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n761), .B(new_n768), .C1(new_n767), .C2(new_n766), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n691), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n691), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n769), .B1(G1961), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G1961), .B2(new_n771), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n774));
  NOR2_X1   g349(.A1(G168), .A2(new_n691), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n691), .A2(G21), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n775), .A2(G1966), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(G1966), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n777), .B(new_n778), .C1(new_n685), .C2(new_n619), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n759), .A2(new_n760), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(KEYINPUT104), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT104), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n759), .A2(new_n783), .A3(new_n760), .A4(new_n780), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n723), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G6), .B(G305), .S(G16), .Z(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT93), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n786), .B(KEYINPUT93), .ZN(new_n790));
  INV_X1    g365(.A(new_n788), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G22), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G166), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT94), .B(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G23), .B(G288), .S(G16), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n789), .A2(new_n792), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n685), .A2(G25), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT90), .ZN(new_n803));
  OAI211_X1 g378(.A(G131), .B(new_n463), .C1(new_n486), .C2(new_n487), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n805), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(G107), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n489), .B2(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT92), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT92), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n809), .A2(new_n816), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n803), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n801), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n824));
  MUX2_X1   g399(.A(G24), .B(G290), .S(G16), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1986), .ZN(new_n826));
  INV_X1    g401(.A(new_n800), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT34), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n823), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n824), .B1(new_n823), .B2(new_n829), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n831), .A2(new_n832), .B1(KEYINPUT95), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n801), .A3(new_n822), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT96), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(KEYINPUT95), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n837), .A3(new_n830), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n785), .B1(new_n834), .B2(new_n838), .ZN(G311));
  AND3_X1   g414(.A1(new_n723), .A2(new_n782), .A3(new_n784), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n836), .A2(new_n837), .A3(new_n830), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n836), .B2(new_n830), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G150));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n844), .A2(new_n537), .B1(new_n528), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n519), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n603), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT107), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  INV_X1    g430(.A(new_n849), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n562), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n850), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n852), .B1(new_n859), .B2(new_n860), .ZN(G145));
  INV_X1    g436(.A(KEYINPUT110), .ZN(new_n862));
  INV_X1    g437(.A(new_n817), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n816), .B1(new_n809), .B2(new_n813), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n623), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n815), .A2(KEYINPUT110), .A3(new_n817), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT109), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n733), .B1(new_n745), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n744), .B(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(KEYINPUT109), .A3(new_n732), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n869), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n863), .A2(new_n864), .A3(new_n862), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT110), .B1(new_n815), .B2(new_n817), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n623), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n875), .B1(new_n881), .B2(new_n868), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n495), .A2(G142), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n489), .A2(G130), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n463), .A2(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n883), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n719), .A2(new_n509), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n716), .A2(G164), .A3(new_n718), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n888), .A2(new_n887), .A3(new_n889), .ZN(new_n891));
  OAI22_X1  g466(.A1(new_n878), .A2(new_n882), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n876), .B1(new_n869), .B2(new_n877), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n891), .A2(new_n890), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n881), .A2(new_n875), .A3(new_n868), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n497), .B(new_n619), .ZN(new_n898));
  XNOR2_X1  g473(.A(G160), .B(KEYINPUT108), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n892), .A2(new_n902), .A3(new_n896), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT40), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n894), .B1(new_n893), .B2(new_n895), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  AND4_X1   g483(.A1(KEYINPUT40), .A2(new_n907), .A3(new_n903), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n904), .A2(new_n909), .ZN(G395));
  XNOR2_X1  g485(.A(new_n562), .B(new_n849), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n610), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n603), .B(G299), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(KEYINPUT41), .ZN(new_n915));
  XNOR2_X1  g490(.A(G299), .B(new_n697), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n914), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(G288), .B(KEYINPUT111), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(G305), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(G166), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n920), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G868), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G868), .B2(new_n849), .ZN(G295));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n849), .ZN(G331));
  NOR2_X1   g504(.A1(new_n857), .A2(G168), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n911), .A2(G286), .ZN(new_n931));
  OAI21_X1  g506(.A(G301), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n857), .A2(G168), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n911), .A2(G286), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(G171), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n913), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n915), .A2(new_n932), .A3(new_n918), .A4(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n924), .ZN(new_n940));
  INV_X1    g515(.A(new_n924), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n908), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n940), .A2(new_n945), .A3(new_n908), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(G397));
  NAND2_X1  g526(.A1(G168), .A2(G8), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n477), .A2(new_n483), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n466), .A2(G2104), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT3), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n472), .B1(new_n956), .B2(new_n480), .ZN(new_n957));
  INV_X1    g532(.A(new_n469), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n463), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n959), .A3(G40), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n509), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT120), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n509), .A2(new_n961), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT120), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n966), .A2(new_n967), .A3(G160), .A4(G40), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1966), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT121), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n509), .A2(new_n974), .A3(new_n961), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n509), .B2(new_n961), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n960), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT122), .B(G2084), .Z(new_n979));
  AOI22_X1  g554(.A1(new_n972), .A2(new_n973), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n970), .A2(KEYINPUT121), .A3(new_n971), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n952), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT115), .B(G1981), .Z(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n590), .A2(new_n591), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT116), .B(G86), .Z(new_n987));
  NAND3_X1  g562(.A1(new_n525), .A2(new_n517), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n588), .A2(new_n511), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n517), .B2(G61), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n986), .B(new_n988), .C1(new_n990), .C2(new_n519), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n991), .A2(new_n992), .A3(G1981), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n991), .B2(G1981), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT49), .B(new_n985), .C1(new_n993), .C2(new_n994), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n960), .A2(new_n964), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n544), .A2(G87), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1003), .A2(G1976), .A3(new_n584), .A4(new_n583), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(G8), .C1(new_n960), .C2(new_n964), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  NAND4_X1  g581(.A1(G160), .A2(G40), .A3(new_n961), .A4(new_n509), .ZN(new_n1007));
  INV_X1    g582(.A(G1976), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(G288), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1007), .A2(G8), .A3(new_n1004), .A4(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(G166), .B2(new_n1000), .ZN(new_n1015));
  OAI211_X1 g590(.A(G8), .B(new_n1013), .C1(new_n520), .C2(new_n530), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n953), .A2(new_n959), .A3(G40), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n969), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n509), .A2(KEYINPUT113), .A3(KEYINPUT45), .A4(new_n961), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1018), .A2(new_n1020), .A3(new_n966), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1971), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n960), .A2(new_n977), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(new_n689), .A3(new_n975), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1000), .B(new_n1017), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1012), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n975), .B(KEYINPUT119), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1024), .B1(new_n1031), .B2(G2090), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G8), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1017), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n982), .A2(new_n1028), .A3(new_n1029), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1032), .A2(G8), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1038), .A2(new_n1012), .A3(new_n1027), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1029), .B1(new_n1039), .B2(new_n982), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT124), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1028), .A2(new_n1034), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n972), .A2(new_n973), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n978), .A2(new_n979), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n981), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(G8), .A3(G168), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT123), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1036), .A4(new_n1035), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1041), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1000), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1036), .B1(new_n1052), .B2(new_n1017), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n982), .A2(new_n1053), .A3(new_n1028), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT127), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1043), .A2(G168), .A3(new_n981), .A4(new_n1044), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1045), .A2(G286), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(G8), .A3(new_n1057), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1061), .B2(KEYINPUT51), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1056), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1022), .B2(G2078), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1025), .A2(new_n975), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n970), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(G301), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1039), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1059), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1057), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(G168), .B1(new_n980), .B2(new_n981), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1064), .A2(new_n1075), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1027), .ZN(new_n1083));
  INV_X1    g658(.A(new_n985), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(G1976), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1002), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1001), .B(KEYINPUT118), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1083), .A2(new_n1012), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1067), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G2067), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n999), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(KEYINPUT126), .A3(KEYINPUT60), .A4(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1092), .B(KEYINPUT60), .C1(new_n978), .C2(G1348), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n978), .A2(G1348), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1092), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1093), .A2(new_n1096), .B1(new_n1100), .B2(new_n603), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT58), .B(G1341), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1022), .A2(G1996), .B1(new_n999), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n563), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(KEYINPUT59), .A3(new_n563), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1096), .A2(new_n1100), .A3(new_n1093), .A4(new_n603), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1031), .A2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT56), .B(G2072), .Z(new_n1113));
  OR2_X1    g688(.A1(new_n1022), .A2(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n578), .A2(KEYINPUT57), .ZN(new_n1116));
  AOI22_X1  g691(.A1(G299), .A2(KEYINPUT57), .B1(new_n574), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n697), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1109), .A2(new_n1110), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  NOR2_X1   g696(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1115), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1120), .A2(new_n1125), .B1(new_n1117), .B2(new_n1115), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n476), .A2(new_n463), .ZN(new_n1128));
  INV_X1    g703(.A(G40), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1071), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1130), .A2(new_n959), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1131), .A2(new_n1020), .A3(new_n966), .A4(new_n1021), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1066), .A2(new_n1132), .A3(new_n1069), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(G171), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1127), .B1(new_n1073), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1070), .A2(G301), .A3(new_n1072), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1127), .B1(new_n1133), .B2(G171), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1039), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1079), .B2(new_n1076), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1088), .B1(new_n1126), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1055), .A2(new_n1082), .A3(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n719), .B(new_n1091), .ZN(new_n1143));
  INV_X1    g718(.A(G1996), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n733), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n960), .A2(new_n966), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT112), .B1(new_n1147), .B2(new_n732), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n1147), .A2(new_n732), .A3(KEYINPUT112), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1145), .A2(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n818), .A2(new_n821), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n820), .B1(new_n815), .B2(new_n817), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(G290), .B(G1986), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1142), .A2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1147), .B(KEYINPUT46), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1143), .A2(new_n733), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1159), .B2(new_n1146), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT47), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1146), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1164), .A2(G1986), .A3(G290), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT48), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1162), .A2(new_n1163), .B1(new_n1154), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n716), .A2(new_n1091), .A3(new_n718), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1164), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1157), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g747(.A(G319), .ZN(new_n1174));
  NOR3_X1   g748(.A1(G401), .A2(new_n1174), .A3(G227), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n683), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1176), .B1(new_n944), .B2(new_n946), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n901), .A2(new_n903), .ZN(new_n1178));
  AND2_X1   g752(.A1(new_n1177), .A2(new_n1178), .ZN(G308));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(G225));
endmodule


