//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT65), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G137), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n457), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n461), .A2(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n462), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(KEYINPUT69), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n484), .A2(new_n458), .A3(new_n460), .A4(new_n466), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n465), .A2(new_n487), .A3(new_n466), .A4(new_n484), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n458), .A2(new_n460), .A3(G126), .A4(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT67), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n465), .A2(new_n493), .A3(G126), .A4(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n492), .B2(new_n494), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT68), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n490), .B1(new_n502), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n507), .A2(new_n509), .A3(new_n514), .A4(new_n516), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n513), .A2(new_n522), .ZN(G166));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  INV_X1    g099(.A(G89), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n518), .A2(new_n524), .B1(new_n525), .B2(new_n521), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n518), .A2(new_n534), .B1(new_n535), .B2(new_n521), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n507), .A2(new_n509), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n536), .B1(G651), .B2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n512), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n518), .A2(new_n544), .B1(new_n545), .B2(new_n521), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT70), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n538), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n521), .ZN(new_n560));
  AOI22_X1  g135(.A1(G651), .A2(new_n559), .B1(new_n560), .B2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(G171), .A2(KEYINPUT71), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n540), .A2(G651), .ZN(new_n564));
  OAI221_X1 g139(.A(new_n564), .B1(new_n534), .B2(new_n518), .C1(new_n535), .C2(new_n521), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  OAI21_X1  g146(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n510), .A2(new_n517), .A3(G87), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n512), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n510), .A2(new_n517), .A3(G86), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n514), .A2(new_n516), .A3(G48), .A4(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(KEYINPUT72), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(KEYINPUT72), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n560), .A2(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n587), .B2(new_n518), .C1(new_n588), .C2(new_n512), .ZN(G290));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT74), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n538), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n517), .A2(G543), .ZN(new_n594));
  AOI22_X1  g169(.A1(G651), .A2(new_n593), .B1(new_n594), .B2(G54), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT73), .B(KEYINPUT10), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n521), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n521), .B2(new_n596), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(new_n568), .ZN(G284));
  OAI21_X1  g180(.A(new_n604), .B1(new_n603), .B2(new_n568), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  NOR2_X1   g185(.A1(new_n602), .A2(G559), .ZN(new_n611));
  INV_X1    g186(.A(new_n602), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(G860), .B2(new_n612), .ZN(G148));
  OR2_X1    g188(.A1(new_n543), .A2(new_n546), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n603), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n611), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n462), .A2(G135), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT77), .Z(new_n619));
  OR2_X1    g194(.A1(new_n466), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n476), .A2(G123), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n465), .A2(new_n471), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT76), .B(KEYINPUT13), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n625), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT81), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n636), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT80), .B(KEYINPUT14), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(G2451), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT82), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n655), .ZN(new_n658));
  INV_X1    g233(.A(new_n654), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT17), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n653), .B2(new_n655), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n658), .B2(KEYINPUT17), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(KEYINPUT84), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(KEYINPUT84), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n666), .A2(new_n667), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  MUX2_X1   g253(.A(new_n678), .B(new_n677), .S(new_n672), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1991), .ZN(new_n682));
  INV_X1    g257(.A(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(G1996), .ZN(new_n687));
  INV_X1    g262(.A(new_n685), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n689), .A3(new_n691), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G16), .A2(G24), .ZN(new_n696));
  XOR2_X1   g271(.A(G290), .B(KEYINPUT86), .Z(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1986), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n476), .A2(G119), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n462), .A2(G131), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n466), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT35), .B(G1991), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(G6), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G305), .B2(G16), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT88), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n709), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n709), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n714), .A2(new_n715), .A3(new_n719), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n708), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT36), .B1(new_n729), .B2(KEYINPUT89), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(KEYINPUT89), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(KEYINPUT89), .A3(KEYINPUT36), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT97), .B(KEYINPUT23), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n709), .A2(G20), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n736), .B(new_n737), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G299), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n742), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT29), .Z(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G21), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G168), .B2(G16), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G1966), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  NOR2_X1   g325(.A1(G5), .A2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT95), .Z(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n565), .B2(new_n709), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n749), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n748), .A2(G1966), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT30), .B(G28), .Z(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n624), .B2(G29), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n754), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n742), .A2(G33), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n465), .A2(G127), .ZN(new_n762));
  NAND2_X1  g337(.A1(G115), .A2(G2104), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n466), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n471), .A2(G103), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT25), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT25), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n764), .B(new_n768), .C1(G139), .C2(new_n462), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n761), .B1(new_n769), .B2(new_n742), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2072), .Z(new_n771));
  INV_X1    g346(.A(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n742), .B1(new_n772), .B2(G34), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(new_n772), .B2(G34), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  INV_X1    g351(.A(G160), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n742), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n746), .A2(new_n760), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n742), .A2(G26), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n476), .A2(G128), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n462), .A2(G140), .ZN(new_n785));
  OR2_X1    g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(new_n742), .ZN(new_n790));
  MUX2_X1   g365(.A(new_n783), .B(new_n790), .S(KEYINPUT28), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G2067), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(G2067), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n745), .A2(new_n741), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n782), .A2(new_n792), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  OR3_X1    g370(.A1(KEYINPUT90), .A2(G4), .A3(G16), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n602), .A2(new_n709), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT90), .B1(G4), .B2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT91), .B(G1348), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n742), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n742), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n799), .A2(new_n800), .B1(G2078), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(G2078), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n803), .B(new_n804), .C1(new_n800), .C2(new_n799), .ZN(new_n805));
  NAND3_X1  g380(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT26), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G105), .B2(new_n471), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n476), .A2(G129), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n462), .A2(G141), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(new_n742), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n814), .A2(new_n815), .B1(G29), .B2(G32), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT27), .B(G1996), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n709), .A2(G19), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n547), .B2(new_n709), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT92), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1341), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n753), .A2(new_n750), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT96), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT96), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n778), .A2(new_n779), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n818), .A2(new_n822), .A3(new_n828), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n795), .A2(new_n805), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n734), .A2(new_n830), .ZN(G150));
  INV_X1    g406(.A(G150), .ZN(G311));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT101), .B(G93), .Z(new_n834));
  OAI22_X1  g409(.A1(new_n518), .A2(new_n833), .B1(new_n521), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n510), .A2(G67), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n512), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n612), .A2(G559), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n846));
  XOR2_X1   g421(.A(new_n845), .B(new_n846), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n835), .B2(new_n838), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n614), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n547), .A2(new_n839), .A3(KEYINPUT102), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n840), .B1(new_n847), .B2(new_n853), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n842), .B1(new_n854), .B2(new_n855), .ZN(G145));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n476), .A2(G130), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n462), .A2(G142), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n466), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(new_n627), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n704), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n769), .B(KEYINPUT103), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n789), .B(new_n811), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n489), .A3(new_n503), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n811), .B(new_n788), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n503), .A2(new_n489), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n769), .A2(KEYINPUT103), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n866), .A2(new_n867), .A3(new_n874), .A4(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  INV_X1    g454(.A(new_n874), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n865), .B(new_n864), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n624), .B(G162), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G160), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n857), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n884), .B2(new_n882), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(G395));
  INV_X1    g463(.A(new_n853), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n611), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n891));
  INV_X1    g466(.A(new_n600), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G299), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n600), .A2(KEYINPUT105), .A3(new_n556), .A4(new_n561), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT105), .B1(new_n608), .B2(new_n600), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n892), .B2(G299), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(KEYINPUT106), .A3(new_n893), .A4(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n890), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n895), .B2(new_n896), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n899), .A2(KEYINPUT41), .A3(new_n893), .A4(new_n894), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n902), .B1(new_n890), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n908));
  NOR2_X1   g483(.A1(G305), .A2(G166), .ZN(new_n909));
  XNOR2_X1  g484(.A(G290), .B(new_n721), .ZN(new_n910));
  AOI21_X1  g485(.A(G303), .B1(new_n583), .B2(new_n584), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n908), .A3(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n913), .ZN(new_n917));
  OAI221_X1 g492(.A(new_n902), .B1(KEYINPUT107), .B2(new_n917), .C1(new_n890), .C2(new_n906), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n915), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n603), .B1(new_n835), .B2(new_n838), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n922), .ZN(G331));
  NOR3_X1   g499(.A1(new_n895), .A2(new_n903), .A3(new_n896), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n565), .A2(G168), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n853), .B(new_n928), .C1(new_n568), .C2(G286), .ZN(new_n929));
  AOI21_X1  g504(.A(G286), .B1(new_n563), .B2(new_n567), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n852), .B(new_n851), .C1(new_n930), .C2(new_n927), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n925), .A2(new_n926), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n904), .A2(KEYINPUT109), .A3(new_n905), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n929), .A2(new_n931), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(KEYINPUT110), .A3(new_n897), .A4(new_n900), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n897), .A2(new_n929), .A3(new_n900), .A4(new_n931), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n914), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n895), .A2(new_n896), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n929), .A3(new_n931), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n935), .B2(new_n906), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n945), .B2(new_n917), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n914), .B(new_n944), .C1(new_n935), .C2(new_n906), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n945), .A2(new_n917), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n954), .A2(new_n948), .A3(new_n942), .A4(new_n857), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT44), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n946), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n932), .A2(new_n933), .B1(new_n937), .B2(new_n938), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n917), .B1(new_n959), .B2(new_n936), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT111), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n942), .B1(new_n941), .B2(new_n946), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n963), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n953), .B1(new_n962), .B2(new_n965), .ZN(G397));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n872), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G113), .A2(G2104), .ZN(new_n972));
  INV_X1    g547(.A(G125), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n461), .B2(new_n973), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n974), .A2(G2105), .B1(G101), .B2(new_n471), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(G40), .A3(new_n469), .A4(new_n464), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n683), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n788), .B(G2067), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(new_n811), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n978), .A2(new_n979), .B1(new_n981), .B2(new_n977), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n979), .B2(new_n978), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n980), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(KEYINPUT114), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(KEYINPUT114), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n811), .B(G1996), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n986), .B(new_n987), .C1(new_n977), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n977), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n704), .B(new_n706), .Z(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR3_X1    g567(.A1(new_n990), .A2(G1986), .A3(G290), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT48), .Z(new_n994));
  OAI21_X1  g569(.A(new_n984), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n704), .A2(new_n706), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n989), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n788), .A2(G2067), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n990), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n970), .B1(G164), .B2(G1384), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n503), .B2(new_n489), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n976), .B1(KEYINPUT45), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1971), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT68), .B1(new_n495), .B2(new_n499), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n501), .B(new_n498), .C1(new_n492), .C2(new_n494), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n489), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1008), .B2(new_n967), .ZN(new_n1009));
  INV_X1    g584(.A(new_n976), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1009), .A2(new_n1011), .A3(G2090), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1002), .ZN(new_n1015));
  INV_X1    g590(.A(G1976), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G288), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT117), .B(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1015), .A2(G8), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1022), .B(new_n1017), .C1(new_n1010), .C2(new_n1002), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n579), .A2(new_n1027), .A3(new_n580), .A4(new_n581), .ZN(new_n1028));
  INV_X1    g603(.A(G86), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n581), .B1(new_n521), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(G1981), .B1(new_n1030), .B2(new_n578), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1031), .A3(KEYINPUT49), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1015), .A2(new_n1037), .A3(G8), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1026), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1032), .B(KEYINPUT118), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n968), .A2(new_n976), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n1022), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1040), .A2(new_n1042), .A3(KEYINPUT119), .A4(new_n1037), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1025), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n1045));
  NOR2_X1   g620(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n1046));
  OR4_X1    g621(.A1(new_n1022), .A2(G166), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(G166), .B2(new_n1022), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1014), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n721), .A2(new_n1016), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1028), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1008), .A2(new_n1005), .A3(new_n967), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n976), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1056), .A2(new_n741), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(G8), .B1(new_n1004), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1049), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1008), .A2(new_n967), .A3(new_n969), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT45), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n976), .B1(new_n968), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1966), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n976), .B1(new_n1005), .B2(new_n1002), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT120), .B(G2084), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n502), .A2(new_n504), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1384), .B1(new_n1070), .B2(new_n489), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1068), .B(new_n1069), .C1(new_n1071), .C2(new_n1005), .ZN(new_n1072));
  AOI211_X1 g647(.A(new_n1022), .B(G286), .C1(new_n1067), .C2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1049), .B(G8), .C1(new_n1004), .C2(new_n1012), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1061), .A2(new_n1073), .A3(new_n1074), .A4(new_n1044), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT63), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1069), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1009), .A2(new_n1011), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1966), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1080));
  OAI21_X1  g655(.A(G8), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1081), .A2(new_n1076), .A3(G286), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1013), .A2(new_n1060), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1074), .A4(new_n1044), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1055), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1086), .B(G8), .C1(new_n1087), .C2(G286), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G168), .A2(new_n1022), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1081), .A2(KEYINPUT51), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT62), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n969), .B1(new_n1008), .B2(new_n967), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1010), .B1(new_n968), .B2(new_n1063), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n718), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1056), .A2(new_n741), .A3(new_n1057), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1022), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1044), .B(new_n1074), .C1(new_n1099), .C2(new_n1049), .ZN(new_n1100));
  INV_X1    g675(.A(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1062), .A2(new_n1101), .A3(new_n1064), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1062), .A2(KEYINPUT124), .A3(new_n1101), .A4(new_n1064), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1104), .A2(KEYINPUT53), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1001), .A2(new_n1101), .A3(new_n1003), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1068), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n750), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n568), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1100), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1088), .A2(new_n1091), .A3(new_n1116), .A4(new_n1092), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1094), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1085), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1107), .A2(new_n1108), .B1(new_n1111), .B2(new_n750), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1104), .A2(KEYINPUT53), .A3(new_n1105), .ZN(new_n1122));
  AOI21_X1  g697(.A(G301), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1124));
  NAND2_X1  g699(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1108), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1003), .A2(new_n971), .A3(new_n1126), .ZN(new_n1127));
  AND4_X1   g702(.A1(G301), .A2(new_n1109), .A3(new_n1112), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1120), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1100), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n1093), .ZN(new_n1131));
  AOI21_X1  g706(.A(G1348), .B1(new_n1110), .B2(new_n1068), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1015), .A2(G2067), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT60), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1138), .B2(new_n892), .ZN(new_n1139));
  INV_X1    g714(.A(G1348), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1133), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT60), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1143), .A2(KEYINPUT123), .A3(new_n600), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1135), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1095), .A2(new_n1096), .A3(G1996), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(G1341), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1041), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n547), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(KEYINPUT59), .B(new_n547), .C1(new_n1146), .C2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT121), .B(G1956), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT56), .B(G2072), .Z(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1001), .A2(new_n1003), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G299), .B(KEYINPUT57), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1158), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1095), .A2(new_n1096), .A3(new_n1159), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1162), .B1(new_n1165), .B2(new_n1157), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT61), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1154), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1138), .A2(new_n1136), .A3(new_n892), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT123), .B1(new_n1143), .B2(new_n600), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT60), .A4(new_n1134), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1164), .A2(new_n1166), .A3(KEYINPUT61), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1145), .A2(new_n1168), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1164), .B(new_n892), .C1(new_n1133), .C2(new_n1132), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1174), .A2(new_n1166), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1131), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT126), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n565), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1121), .A2(KEYINPUT126), .A3(new_n1127), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT127), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1178), .A2(new_n1182), .A3(new_n1179), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1120), .B1(new_n1184), .B2(G301), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1181), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1119), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n977), .A2(G1986), .A3(G290), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n993), .A2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT113), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n992), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT115), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1000), .B1(new_n1187), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(new_n951), .ZN(new_n1195));
  INV_X1    g769(.A(G319), .ZN(new_n1196));
  NOR3_X1   g770(.A1(G401), .A2(new_n1196), .A3(G227), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n693), .A2(new_n1197), .A3(new_n694), .ZN(new_n1198));
  NOR3_X1   g772(.A1(new_n1195), .A2(new_n1198), .A3(new_n886), .ZN(G308));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n886), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1200), .A2(new_n951), .ZN(G225));
endmodule


