//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n206), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n205), .B1(new_n210), .B2(new_n206), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(G148gat), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n220), .A2(new_n222), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G155gat), .B(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n217), .A2(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n228), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n215), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n223), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(new_n224), .ZN(new_n241));
  XNOR2_X1  g040(.A(G141gat), .B(G148gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n222), .ZN(new_n245));
  AND2_X1   g044(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(new_n248), .B2(G148gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n240), .B1(new_n225), .B2(new_n224), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(KEYINPUT85), .B(new_n238), .C1(new_n212), .C2(new_n213), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n236), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n206), .A2(new_n210), .ZN(new_n254));
  INV_X1    g053(.A(new_n205), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT29), .B1(new_n256), .B2(new_n211), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(KEYINPUT85), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n251), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n239), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(KEYINPUT86), .B(new_n251), .C1(new_n253), .C2(new_n258), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n204), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n239), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT78), .B1(new_n227), .B2(new_n234), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n244), .B(new_n266), .C1(new_n249), .C2(new_n250), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n265), .B(new_n267), .C1(new_n257), .C2(KEYINPUT3), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n264), .A2(new_n204), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(G22gat), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n204), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT3), .B1(new_n257), .B2(KEYINPUT85), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n214), .B2(KEYINPUT29), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n235), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n264), .B1(new_n275), .B2(KEYINPUT86), .ZN(new_n276));
  INV_X1    g075(.A(new_n262), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G22gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n269), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n270), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n260), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n262), .A3(new_n264), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n269), .B1(new_n284), .B2(new_n271), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT87), .B1(new_n285), .B2(new_n279), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G50gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G78gat), .B(G106gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n282), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n270), .A2(new_n281), .A3(KEYINPUT87), .A4(new_n290), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT73), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  OR2_X1    g099(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT27), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n301), .A2(new_n303), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT28), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  AND2_X1   g108(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT27), .B(G183gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT26), .ZN(new_n316));
  INV_X1    g115(.A(G169gat), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n319), .B(new_n320), .C1(new_n317), .C2(new_n318), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n308), .A2(new_n309), .A3(new_n315), .A4(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT23), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT23), .B1(new_n317), .B2(new_n318), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n317), .A2(new_n318), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n329), .B(new_n330), .C1(G183gat), .C2(G190gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n335), .A2(KEYINPUT24), .ZN(new_n336));
  AND3_X1   g135(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n330), .B(new_n334), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n327), .B1(new_n338), .B2(new_n326), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT71), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n330), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n337), .A2(new_n335), .A3(KEYINPUT24), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n326), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT25), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT71), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n322), .A4(new_n332), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n300), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n333), .A2(new_n339), .ZN(new_n349));
  INV_X1    g148(.A(new_n300), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n349), .A2(KEYINPUT29), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n214), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n340), .A2(new_n238), .A3(new_n346), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n300), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n349), .A2(new_n300), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n299), .B(new_n353), .C1(new_n361), .C2(new_n214), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT30), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n298), .B(KEYINPUT74), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n359), .B1(new_n355), .B2(new_n356), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n215), .B1(new_n366), .B2(new_n358), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n367), .B2(new_n353), .ZN(new_n368));
  INV_X1    g167(.A(new_n353), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n354), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT72), .B1(new_n354), .B2(new_n300), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n370), .A2(new_n371), .A3(new_n359), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n298), .B(new_n369), .C1(new_n372), .C2(new_n215), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(KEYINPUT75), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n364), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT3), .ZN(new_n377));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G113gat), .A2(G120gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT1), .ZN(new_n380));
  NAND2_X1  g179(.A1(G113gat), .A2(G120gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G134gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n383), .A2(G127gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(G127gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(G113gat), .B2(G120gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n381), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n384), .A2(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n235), .B2(new_n236), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n377), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n391), .A3(KEYINPUT79), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n382), .A2(new_n389), .ZN(new_n397));
  OR3_X1    g196(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n235), .A2(new_n390), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n265), .A2(new_n267), .A3(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(new_n403), .A3(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(KEYINPUT39), .A3(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G57gat), .B(G85gat), .Z(new_n409));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  INV_X1    g212(.A(KEYINPUT39), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n402), .A2(new_n414), .A3(new_n404), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT40), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n406), .A2(new_n399), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n404), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT81), .B1(new_n420), .B2(KEYINPUT5), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n403), .B1(new_n406), .B2(new_n399), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n377), .A2(new_n391), .A3(KEYINPUT79), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT79), .B1(new_n377), .B2(new_n391), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n403), .B(new_n401), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT80), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n396), .A2(new_n431), .A3(new_n403), .A4(new_n401), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n429), .A2(KEYINPUT5), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n413), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n408), .A2(KEYINPUT40), .A3(new_n413), .A4(new_n415), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n418), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n294), .B1(new_n376), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT37), .B1(new_n367), .B2(new_n353), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT37), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n441), .B(new_n369), .C1(new_n372), .C2(new_n215), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n442), .A3(new_n299), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n362), .B1(new_n443), .B2(KEYINPUT38), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n433), .A2(new_n434), .ZN(new_n445));
  INV_X1    g244(.A(new_n413), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(KEYINPUT6), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n435), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n413), .A3(new_n434), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n365), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n353), .B1(new_n361), .B2(new_n214), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(new_n441), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n357), .A2(new_n215), .A3(new_n358), .A4(new_n360), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT88), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n366), .A2(new_n461), .A3(new_n215), .A4(new_n358), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n348), .A2(new_n352), .A3(new_n214), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n458), .B1(new_n464), .B2(new_n441), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n451), .A3(new_n454), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n439), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n453), .A2(new_n452), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n449), .A2(new_n450), .B1(new_n468), .B2(new_n436), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n294), .B1(new_n469), .B2(new_n376), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT70), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT36), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n344), .A2(new_n390), .A3(new_n322), .A4(new_n332), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n322), .A2(new_n332), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT66), .A3(new_n390), .A4(new_n344), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n397), .B1(new_n333), .B2(new_n339), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(G227gat), .A2(G233gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G71gat), .B(G99gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT68), .ZN(new_n486));
  INV_X1    g285(.A(G15gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n488), .A2(G43gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(G43gat), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT33), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND4_X1   g290(.A1(new_n475), .A2(new_n484), .A3(KEYINPUT32), .A4(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n482), .B2(new_n483), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n475), .B1(new_n494), .B2(new_n491), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n482), .A2(new_n483), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n494), .A2(KEYINPUT67), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n489), .A2(new_n490), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT33), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n484), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n496), .A2(new_n499), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n499), .B1(new_n496), .B2(new_n507), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n473), .B(new_n474), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n496), .A2(new_n507), .ZN(new_n511));
  INV_X1    g310(.A(new_n499), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n499), .A3(new_n507), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n513), .A2(new_n471), .A3(new_n472), .A4(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n467), .A2(new_n470), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT35), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n364), .A2(new_n368), .A3(new_n375), .ZN(new_n519));
  INV_X1    g318(.A(new_n450), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT83), .B1(new_n435), .B2(KEYINPUT6), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n454), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n294), .A2(new_n508), .A3(new_n509), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n518), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n469), .A2(new_n376), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT35), .A3(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n517), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT13), .ZN(new_n532));
  XOR2_X1   g331(.A(G15gat), .B(G22gat), .Z(new_n533));
  INV_X1    g332(.A(G1gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT16), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(G1gat), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT91), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT91), .A3(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(KEYINPUT91), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n535), .A2(new_n538), .A3(new_n543), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G29gat), .ZN(new_n546));
  INV_X1    g345(.A(G36gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT14), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(G29gat), .B2(G36gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(G29gat), .A2(G36gat), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G43gat), .ZN(new_n553));
  INV_X1    g352(.A(G50gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  NAND2_X1  g355(.A1(G43gat), .A2(G50gat), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(KEYINPUT90), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n560));
  INV_X1    g359(.A(new_n557), .ZN(new_n561));
  NOR2_X1   g360(.A1(G43gat), .A2(G50gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(KEYINPUT89), .A3(new_n557), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT15), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT90), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n545), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n552), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n565), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n542), .A2(new_n574), .A3(new_n575), .A4(new_n544), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n532), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT17), .B1(new_n566), .B2(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n579), .A3(new_n575), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n580), .A3(new_n545), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n531), .A3(new_n576), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n581), .A2(KEYINPUT18), .A3(new_n531), .A4(new_n576), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n585), .A2(KEYINPUT92), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(KEYINPUT92), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT11), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(new_n317), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n591), .A2(G197gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(G197gat), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n592), .A2(KEYINPUT12), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT12), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n596), .B(new_n584), .C1(new_n586), .C2(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n530), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G57gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(G64gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n607));
  INV_X1    g406(.A(G64gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(G57gat), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n606), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT96), .B1(new_n608), .B2(G57gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  INV_X1    g412(.A(G71gat), .ZN(new_n614));
  INV_X1    g413(.A(G78gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT9), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n617), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n609), .B2(new_n606), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(new_n614), .A3(new_n615), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n613), .A2(KEYINPUT93), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(G71gat), .A3(G78gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n622), .A2(new_n624), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n621), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n622), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(KEYINPUT95), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n619), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n636), .A2(KEYINPUT97), .A3(KEYINPUT21), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT97), .B1(new_n636), .B2(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n637), .A2(new_n642), .A3(new_n638), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n604), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n636), .A2(KEYINPUT21), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n545), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(KEYINPUT98), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(KEYINPUT98), .ZN(new_n650));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n650), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n653), .B1(new_n656), .B2(new_n648), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n604), .A3(new_n643), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n645), .A2(new_n655), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n655), .ZN(new_n660));
  INV_X1    g459(.A(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n644), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n566), .A2(new_n571), .ZN(new_n664));
  NAND2_X1  g463(.A1(G85gat), .A2(G92gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT7), .ZN(new_n666));
  XNOR2_X1  g465(.A(G99gat), .B(G106gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(G99gat), .A2(G106gat), .ZN(new_n668));
  INV_X1    g467(.A(G85gat), .ZN(new_n669));
  INV_X1    g468(.A(G92gat), .ZN(new_n670));
  AOI22_X1  g469(.A1(KEYINPUT8), .A2(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n666), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n667), .B1(new_n666), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(G232gat), .A2(G233gat), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n664), .A2(new_n674), .B1(KEYINPUT41), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n578), .A2(new_n580), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT99), .ZN(new_n680));
  XNOR2_X1  g479(.A(G190gat), .B(G218gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n679), .B(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n675), .A2(KEYINPUT41), .ZN(new_n687));
  XNOR2_X1  g486(.A(G134gat), .B(G162gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n682), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n682), .A2(new_n686), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n689), .B(new_n690), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n663), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n682), .A2(new_n686), .A3(new_n691), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n694), .B1(new_n682), .B2(new_n686), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n659), .A2(new_n662), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT101), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(G230gat), .A2(G233gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n677), .A2(new_n635), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT10), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n633), .A2(KEYINPUT95), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n628), .A2(new_n629), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n621), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n674), .A2(new_n709), .A3(new_n619), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n636), .A2(KEYINPUT10), .A3(new_n674), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT102), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT102), .B1(new_n711), .B2(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n704), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n705), .A2(new_n710), .ZN(new_n717));
  INV_X1    g516(.A(new_n704), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(G176gat), .B(G204gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G148gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT103), .B(G120gat), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n721), .B(new_n722), .Z(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n716), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n711), .A2(new_n712), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n719), .B1(new_n727), .B2(new_n718), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n723), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n703), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n602), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n522), .A2(KEYINPUT104), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n522), .A2(KEYINPUT104), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT105), .B(G1gat), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1324gat));
  INV_X1    g538(.A(new_n732), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n376), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT16), .B(G8gat), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(G8gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(G1325gat));
  AND3_X1   g546(.A1(new_n510), .A2(new_n515), .A3(KEYINPUT106), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT106), .B1(new_n510), .B2(new_n515), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G15gat), .B1(new_n732), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n508), .A2(new_n509), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n487), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n732), .B2(new_n753), .ZN(G1326gat));
  INV_X1    g553(.A(new_n294), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n732), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT43), .B(G22gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT107), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n756), .B(new_n758), .ZN(G1327gat));
  INV_X1    g558(.A(new_n730), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n663), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n700), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT108), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n602), .A2(new_n546), .A3(new_n735), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT45), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n517), .B2(new_n529), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n761), .A2(new_n600), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT109), .Z(new_n770));
  AOI21_X1  g569(.A(KEYINPUT35), .B1(new_n527), .B2(new_n524), .ZN(new_n771));
  AND4_X1   g570(.A1(KEYINPUT35), .A2(new_n524), .A3(new_n519), .A4(new_n522), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n467), .B(new_n470), .C1(new_n748), .C2(new_n749), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n695), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n768), .B(new_n770), .C1(new_n775), .C2(KEYINPUT44), .ZN(new_n776));
  OAI21_X1  g575(.A(G29gat), .B1(new_n776), .B2(new_n736), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n766), .A2(new_n777), .ZN(G1328gat));
  NAND4_X1  g577(.A1(new_n602), .A2(new_n547), .A3(new_n376), .A4(new_n764), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT46), .Z(new_n780));
  OAI21_X1  g579(.A(G36gat), .B1(new_n776), .B2(new_n519), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1329gat));
  OAI21_X1  g581(.A(G43gat), .B1(new_n776), .B2(new_n750), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n602), .A2(new_n553), .A3(new_n752), .A4(new_n764), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT47), .B1(new_n784), .B2(KEYINPUT110), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1330gat));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n788));
  OAI21_X1  g587(.A(G50gat), .B1(new_n776), .B2(new_n755), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n294), .A2(new_n554), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT111), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n602), .A2(new_n764), .A3(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n789), .B2(new_n793), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n788), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n789), .A2(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n789), .A2(new_n793), .A3(new_n790), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT48), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n796), .A2(new_n800), .ZN(G1331gat));
  NAND2_X1  g600(.A1(new_n773), .A2(new_n774), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n703), .A2(new_n601), .A3(new_n760), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n736), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT113), .B(G57gat), .Z(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1332gat));
  NOR2_X1   g606(.A1(new_n804), .A2(new_n519), .ZN(new_n808));
  NOR2_X1   g607(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n809));
  AND2_X1   g608(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n808), .B2(new_n809), .ZN(G1333gat));
  OAI21_X1  g611(.A(G71gat), .B1(new_n804), .B2(new_n750), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n752), .A2(new_n614), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g615(.A1(new_n804), .A2(new_n755), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(new_n615), .ZN(G1335gat));
  NOR2_X1   g617(.A1(new_n663), .A2(new_n600), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n775), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n819), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n730), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n669), .A3(new_n735), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n775), .A2(KEYINPUT44), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n663), .A2(new_n600), .A3(new_n730), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n768), .A4(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n768), .B(new_n827), .C1(new_n775), .C2(KEYINPUT44), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n735), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n825), .B1(new_n833), .B2(new_n669), .ZN(G1336gat));
  NOR2_X1   g633(.A1(new_n519), .A2(G92gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n837));
  OAI21_X1  g636(.A(G92gat), .B1(new_n829), .B2(new_n519), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n828), .A2(new_n376), .A3(new_n831), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n840), .A2(G92gat), .B1(new_n824), .B2(new_n835), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n841), .B2(new_n837), .ZN(G1337gat));
  AOI21_X1  g641(.A(G99gat), .B1(new_n824), .B2(new_n752), .ZN(new_n843));
  INV_X1    g642(.A(G99gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n750), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n832), .B2(new_n845), .ZN(G1338gat));
  NOR2_X1   g645(.A1(new_n755), .A2(G106gat), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT53), .B1(new_n824), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G106gat), .B1(new_n829), .B2(new_n755), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT115), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n823), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT51), .B1(new_n775), .B2(new_n819), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n760), .B(new_n847), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n854));
  AND4_X1   g653(.A1(KEYINPUT115), .A2(new_n853), .A3(new_n854), .A4(new_n849), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n828), .A2(new_n294), .A3(new_n831), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n856), .A2(G106gat), .B1(new_n824), .B2(new_n847), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n850), .A2(new_n855), .B1(new_n857), .B2(new_n854), .ZN(G1339gat));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n726), .B2(new_n704), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT102), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n726), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n713), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n704), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n726), .A2(new_n865), .A3(new_n704), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(KEYINPUT55), .A3(new_n723), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n859), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n716), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n867), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT116), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n725), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n725), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n864), .B1(new_n863), .B2(new_n867), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n871), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT117), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n723), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n863), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n875), .A2(new_n880), .A3(new_n600), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n592), .A2(new_n593), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n572), .A2(new_n576), .A3(new_n532), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n531), .B1(new_n581), .B2(new_n576), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n599), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n730), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n700), .B1(new_n884), .B2(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n698), .A2(new_n699), .A3(new_n889), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n875), .A2(new_n880), .A3(new_n883), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n701), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n697), .A2(new_n702), .A3(new_n601), .A4(new_n730), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n525), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n736), .A2(new_n376), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n600), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n760), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g704(.A1(new_n900), .A2(new_n701), .ZN(new_n906));
  XOR2_X1   g705(.A(KEYINPUT118), .B(G127gat), .Z(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(G1342gat));
  NOR2_X1   g707(.A1(new_n900), .A2(new_n695), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n383), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n911), .A3(new_n383), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT119), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(KEYINPUT119), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n909), .B2(new_n383), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT120), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1343gat));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n899), .A2(new_n750), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n755), .B1(new_n896), .B2(new_n897), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(KEYINPUT57), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923));
  AND4_X1   g722(.A1(new_n601), .A2(new_n697), .A3(new_n702), .A4(new_n730), .ZN(new_n924));
  AOI221_X4 g723(.A(new_n876), .B1(new_n598), .B2(new_n599), .C1(new_n877), .C2(new_n878), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n883), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n890), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n894), .B1(new_n928), .B2(new_n700), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n924), .B1(new_n929), .B2(new_n701), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n755), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n923), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n883), .B(KEYINPUT121), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n879), .A2(new_n600), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n891), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n695), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n663), .B1(new_n938), .B2(new_n894), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT122), .B(new_n932), .C1(new_n939), .C2(new_n924), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n600), .B(new_n920), .C1(new_n922), .C2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n248), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n919), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n899), .A2(new_n750), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n896), .A2(new_n897), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n294), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n600), .A2(new_n217), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n949), .B1(new_n942), .B2(new_n943), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n944), .A2(new_n950), .A3(KEYINPUT58), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT58), .ZN(new_n952));
  AOI221_X4 g751(.A(new_n949), .B1(new_n919), .B2(new_n952), .C1(new_n942), .C2(new_n943), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n953), .ZN(G1344gat));
  NAND4_X1  g753(.A1(new_n920), .A2(new_n221), .A3(new_n760), .A4(new_n921), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n947), .A2(KEYINPUT57), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n897), .B(KEYINPUT124), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n931), .B(new_n294), .C1(new_n958), .C2(new_n939), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n957), .A2(new_n760), .A3(new_n920), .A4(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n221), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n922), .A2(new_n941), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n945), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT59), .B(new_n221), .C1(new_n966), .C2(new_n760), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n955), .B1(new_n964), .B2(new_n967), .ZN(G1345gat));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n663), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G155gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n920), .A2(new_n921), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n701), .A2(G155gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(G1346gat));
  INV_X1    g772(.A(G162gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n966), .B2(new_n700), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n971), .A2(G162gat), .A3(new_n695), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n975), .A2(new_n976), .ZN(G1347gat));
  NOR2_X1   g776(.A1(new_n735), .A2(new_n519), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n898), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n979), .A2(new_n601), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(new_n317), .ZN(G1348gat));
  NOR2_X1   g780(.A1(new_n979), .A2(new_n730), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(new_n318), .ZN(G1349gat));
  NOR2_X1   g782(.A1(new_n979), .A2(new_n701), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n302), .A2(KEYINPUT126), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n313), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(KEYINPUT126), .A2(G183gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g788(.A1(new_n898), .A2(new_n700), .A3(new_n978), .ZN(new_n990));
  INV_X1    g789(.A(new_n312), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n990), .A2(G190gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n993), .B2(new_n994), .ZN(G1351gat));
  AND2_X1   g795(.A1(new_n978), .A2(new_n750), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n957), .A2(new_n959), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n600), .A2(G197gat), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n997), .A2(new_n921), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n1000), .A2(new_n601), .ZN(new_n1001));
  OAI22_X1  g800(.A1(new_n998), .A2(new_n999), .B1(new_n1001), .B2(G197gat), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(G1352gat));
  NAND3_X1  g802(.A1(new_n957), .A2(new_n760), .A3(new_n959), .ZN(new_n1004));
  INV_X1    g803(.A(new_n997), .ZN(new_n1005));
  OAI21_X1  g804(.A(G204gat), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n730), .A2(G204gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n997), .A2(new_n921), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1009));
  OR2_X1    g808(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n1006), .A2(KEYINPUT127), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1353gat));
  OR2_X1    g814(.A1(new_n998), .A2(new_n701), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT63), .B1(new_n1016), .B2(G211gat), .ZN(new_n1017));
  OAI211_X1 g816(.A(KEYINPUT63), .B(G211gat), .C1(new_n998), .C2(new_n701), .ZN(new_n1018));
  INV_X1    g817(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n663), .A2(new_n208), .ZN(new_n1020));
  OAI22_X1  g819(.A1(new_n1017), .A2(new_n1019), .B1(new_n1000), .B2(new_n1020), .ZN(G1354gat));
  OAI21_X1  g820(.A(new_n209), .B1(new_n1000), .B2(new_n695), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n700), .A2(G218gat), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1022), .B1(new_n998), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g823(.A(new_n1024), .ZN(G1355gat));
endmodule


