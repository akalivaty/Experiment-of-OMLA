

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U554 ( .A(n711), .ZN(n695) );
  NOR2_X1 U555 ( .A1(G2104), .A2(n623), .ZN(n746) );
  NOR2_X1 U556 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n528) );
  INV_X1 U557 ( .A(G2105), .ZN(n623) );
  NOR2_X1 U558 ( .A1(n624), .A2(n623), .ZN(n749) );
  NOR2_X2 U559 ( .A1(n809), .A2(G1384), .ZN(n630) );
  AND2_X1 U560 ( .A1(n552), .A2(n521), .ZN(n548) );
  AND2_X1 U561 ( .A1(n538), .A2(n537), .ZN(n536) );
  OR2_X1 U562 ( .A1(n689), .A2(n534), .ZN(n537) );
  AND2_X2 U563 ( .A1(n618), .A2(G2104), .ZN(n919) );
  NAND2_X1 U564 ( .A1(G8), .A2(n711), .ZN(n740) );
  INV_X1 U565 ( .A(n688), .ZN(n542) );
  INV_X1 U566 ( .A(KEYINPUT32), .ZN(n551) );
  INV_X1 U567 ( .A(G2105), .ZN(n531) );
  INV_X1 U568 ( .A(G2104), .ZN(n532) );
  AND2_X1 U569 ( .A1(n526), .A2(n554), .ZN(n553) );
  OR2_X1 U570 ( .A1(n558), .A2(KEYINPUT33), .ZN(n554) );
  OR2_X1 U571 ( .A1(n863), .A2(n640), .ZN(n765) );
  NAND2_X1 U572 ( .A1(n831), .A2(G51), .ZN(n567) );
  NAND2_X1 U573 ( .A1(G102), .A2(n919), .ZN(n619) );
  NAND2_X1 U574 ( .A1(n542), .A2(KEYINPUT29), .ZN(n541) );
  NAND2_X1 U575 ( .A1(n536), .A2(n535), .ZN(n700) );
  INV_X1 U576 ( .A(KEYINPUT101), .ZN(n709) );
  NAND2_X1 U577 ( .A1(n551), .A2(n550), .ZN(n549) );
  INV_X1 U578 ( .A(G8), .ZN(n550) );
  INV_X1 U579 ( .A(n740), .ZN(n558) );
  XNOR2_X1 U580 ( .A(n729), .B(KEYINPUT102), .ZN(n730) );
  INV_X1 U581 ( .A(n1011), .ZN(n732) );
  XNOR2_X1 U582 ( .A(n630), .B(KEYINPUT64), .ZN(n764) );
  NOR2_X1 U583 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n530) );
  INV_X1 U585 ( .A(KEYINPUT104), .ZN(n744) );
  AND2_X1 U586 ( .A1(n556), .A2(n522), .ZN(n745) );
  XNOR2_X1 U587 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U588 ( .A(n574), .B(KEYINPUT76), .ZN(n575) );
  NOR2_X2 U589 ( .A1(G651), .A2(G543), .ZN(n827) );
  INV_X1 U590 ( .A(KEYINPUT23), .ZN(n633) );
  XOR2_X1 U591 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U592 ( .A(n698), .ZN(n544) );
  AND2_X1 U593 ( .A1(n725), .A2(n549), .ZN(n521) );
  AND2_X1 U594 ( .A1(n743), .A2(n742), .ZN(n522) );
  AND2_X1 U595 ( .A1(n688), .A2(n545), .ZN(n523) );
  NOR2_X1 U596 ( .A1(n698), .A2(n545), .ZN(n524) );
  AND2_X1 U597 ( .A1(n523), .A2(n544), .ZN(n525) );
  NOR2_X1 U598 ( .A1(n733), .A2(n732), .ZN(n526) );
  INV_X1 U599 ( .A(KEYINPUT29), .ZN(n545) );
  AND2_X1 U600 ( .A1(KEYINPUT32), .A2(G8), .ZN(n527) );
  INV_X1 U601 ( .A(KEYINPUT33), .ZN(n557) );
  NAND2_X1 U602 ( .A1(n528), .A2(n623), .ZN(n533) );
  NAND2_X1 U603 ( .A1(n533), .A2(n529), .ZN(n631) );
  NAND2_X1 U604 ( .A1(n530), .A2(KEYINPUT17), .ZN(n529) );
  NAND2_X1 U605 ( .A1(n524), .A2(n693), .ZN(n534) );
  NAND2_X1 U606 ( .A1(n689), .A2(n525), .ZN(n535) );
  NAND2_X1 U607 ( .A1(n539), .A2(n544), .ZN(n538) );
  AND2_X1 U608 ( .A1(n543), .A2(n540), .ZN(n539) );
  NAND2_X1 U609 ( .A1(n693), .A2(n541), .ZN(n540) );
  OR2_X1 U610 ( .A1(n693), .A2(n545), .ZN(n543) );
  NAND2_X1 U611 ( .A1(n548), .A2(n546), .ZN(n738) );
  NAND2_X1 U612 ( .A1(n547), .A2(n551), .ZN(n546) );
  INV_X1 U613 ( .A(n717), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n717), .A2(n527), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n738), .A2(n727), .ZN(n728) );
  NAND2_X1 U616 ( .A1(n555), .A2(n553), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n730), .A2(n557), .ZN(n555) );
  INV_X1 U618 ( .A(G2104), .ZN(n624) );
  AND2_X1 U619 ( .A1(n779), .A2(n789), .ZN(n559) );
  NOR2_X1 U620 ( .A1(n643), .A2(n781), .ZN(n642) );
  INV_X1 U621 ( .A(KEYINPUT100), .ZN(n699) );
  XNOR2_X1 U622 ( .A(KEYINPUT93), .B(n765), .ZN(n641) );
  OR2_X1 U623 ( .A1(n862), .A2(n639), .ZN(n640) );
  INV_X1 U624 ( .A(KEYINPUT13), .ZN(n647) );
  INV_X1 U625 ( .A(KEYINPUT6), .ZN(n574) );
  INV_X1 U626 ( .A(G2105), .ZN(n618) );
  BUF_X1 U627 ( .A(n746), .Z(n926) );
  INV_X1 U628 ( .A(KEYINPUT65), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n655), .A2(n654), .ZN(n812) );
  BUF_X1 U630 ( .A(n812), .Z(n1018) );
  NAND2_X1 U631 ( .A1(n827), .A2(G89), .ZN(n560) );
  XNOR2_X1 U632 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  XOR2_X1 U633 ( .A(KEYINPUT0), .B(G543), .Z(n564) );
  INV_X1 U634 ( .A(G651), .ZN(n568) );
  NOR2_X2 U635 ( .A1(n564), .A2(n568), .ZN(n826) );
  NAND2_X1 U636 ( .A1(G76), .A2(n826), .ZN(n561) );
  NAND2_X1 U637 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U638 ( .A(KEYINPUT5), .B(n563), .Z(n578) );
  NOR2_X1 U639 ( .A1(G651), .A2(n564), .ZN(n566) );
  XNOR2_X2 U640 ( .A(n566), .B(n565), .ZN(n831) );
  XNOR2_X1 U641 ( .A(KEYINPUT75), .B(n567), .ZN(n573) );
  NOR2_X1 U642 ( .A1(G543), .A2(n568), .ZN(n569) );
  XOR2_X1 U643 ( .A(KEYINPUT1), .B(n569), .Z(n649) );
  INV_X1 U644 ( .A(n649), .ZN(n570) );
  INV_X1 U645 ( .A(n570), .ZN(n830) );
  NAND2_X1 U646 ( .A1(n830), .A2(G63), .ZN(n571) );
  XOR2_X1 U647 ( .A(n571), .B(KEYINPUT74), .Z(n572) );
  NOR2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n576) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U650 ( .A(n579), .B(KEYINPUT7), .ZN(n580) );
  XNOR2_X1 U651 ( .A(n580), .B(KEYINPUT77), .ZN(G168) );
  NAND2_X1 U652 ( .A1(n827), .A2(G90), .ZN(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT67), .B(n581), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n826), .A2(G77), .ZN(n582) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n582), .Z(n583) );
  NOR2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U657 ( .A(KEYINPUT69), .B(n585), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT9), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G64), .A2(n830), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G52), .A2(n831), .ZN(n587) );
  AND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(G301) );
  NAND2_X1 U663 ( .A1(G75), .A2(n826), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G88), .A2(n827), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G62), .A2(n830), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G50), .A2(n831), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(G166) );
  INV_X1 U670 ( .A(G166), .ZN(G303) );
  NAND2_X1 U671 ( .A1(G49), .A2(n831), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G74), .A2(G651), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n830), .A2(n599), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n600), .B(KEYINPUT82), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G87), .A2(n564), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U678 ( .A(KEYINPUT83), .B(n603), .Z(G288) );
  NAND2_X1 U679 ( .A1(G86), .A2(n827), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G61), .A2(n830), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n826), .A2(G73), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT2), .B(n606), .Z(n607) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n831), .A2(G48), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(G305) );
  NAND2_X1 U687 ( .A1(G72), .A2(n826), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G85), .A2(n827), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G47), .A2(n831), .ZN(n613) );
  XOR2_X1 U691 ( .A(KEYINPUT66), .B(n613), .Z(n614) );
  NOR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n830), .A2(G60), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(G290) );
  NAND2_X1 U695 ( .A1(n631), .A2(G138), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n622) );
  INV_X1 U697 ( .A(KEYINPUT89), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G126), .A2(n746), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n749), .A2(G114), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT88), .ZN(n628) );
  NOR2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n809) );
  INV_X1 U704 ( .A(n631), .ZN(n632) );
  INV_X2 U705 ( .A(n632), .ZN(n921) );
  NAND2_X1 U706 ( .A1(n921), .A2(G137), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n919), .A2(G101), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n863) );
  NAND2_X1 U710 ( .A1(G125), .A2(n746), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G113), .A2(n749), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n862) );
  INV_X1 U713 ( .A(G40), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n764), .A2(n641), .ZN(n643) );
  INV_X1 U715 ( .A(G1996), .ZN(n781) );
  XNOR2_X1 U716 ( .A(n642), .B(KEYINPUT26), .ZN(n659) );
  NAND2_X1 U717 ( .A1(n643), .A2(G1341), .ZN(n657) );
  NAND2_X1 U718 ( .A1(G68), .A2(n826), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n827), .A2(G81), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n644), .B(KEYINPUT12), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n653) );
  NAND2_X1 U723 ( .A1(G56), .A2(n649), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n650), .B(KEYINPUT14), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT71), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n831), .A2(G43), .ZN(n654) );
  INV_X1 U727 ( .A(n812), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n674) );
  NAND2_X1 U730 ( .A1(G54), .A2(n831), .ZN(n666) );
  NAND2_X1 U731 ( .A1(G79), .A2(n826), .ZN(n661) );
  NAND2_X1 U732 ( .A1(G66), .A2(n830), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U734 ( .A1(G92), .A2(n827), .ZN(n662) );
  XNOR2_X1 U735 ( .A(KEYINPUT73), .B(n662), .ZN(n663) );
  NOR2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X2 U738 ( .A(n667), .B(KEYINPUT15), .ZN(n1014) );
  NAND2_X1 U739 ( .A1(n674), .A2(n1014), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(KEYINPUT96), .ZN(n672) );
  BUF_X2 U741 ( .A(n643), .Z(n711) );
  NOR2_X1 U742 ( .A1(n695), .A2(G1348), .ZN(n670) );
  NOR2_X1 U743 ( .A1(G2067), .A2(n711), .ZN(n669) );
  NOR2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n673), .B(KEYINPUT97), .ZN(n677) );
  NOR2_X1 U747 ( .A1(n1014), .A2(n674), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(KEYINPUT98), .ZN(n676) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U750 ( .A(n678), .B(KEYINPUT99), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n695), .A2(G2072), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n679), .B(KEYINPUT27), .ZN(n681) );
  INV_X1 U753 ( .A(G1956), .ZN(n1043) );
  NOR2_X1 U754 ( .A1(n1043), .A2(n695), .ZN(n680) );
  NOR2_X1 U755 ( .A1(n681), .A2(n680), .ZN(n690) );
  NAND2_X1 U756 ( .A1(G65), .A2(n830), .ZN(n683) );
  NAND2_X1 U757 ( .A1(G53), .A2(n831), .ZN(n682) );
  NAND2_X1 U758 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U759 ( .A1(G78), .A2(n826), .ZN(n685) );
  NAND2_X1 U760 ( .A1(G91), .A2(n827), .ZN(n684) );
  NAND2_X1 U761 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U762 ( .A1(n687), .A2(n686), .ZN(n1021) );
  NAND2_X1 U763 ( .A1(n690), .A2(n1021), .ZN(n688) );
  NOR2_X1 U764 ( .A1(n690), .A2(n1021), .ZN(n692) );
  XNOR2_X1 U765 ( .A(KEYINPUT28), .B(KEYINPUT95), .ZN(n691) );
  XNOR2_X1 U766 ( .A(n692), .B(n691), .ZN(n693) );
  XOR2_X1 U767 ( .A(G2078), .B(KEYINPUT25), .Z(n694) );
  XNOR2_X1 U768 ( .A(KEYINPUT94), .B(n694), .ZN(n990) );
  NOR2_X1 U769 ( .A1(n711), .A2(n990), .ZN(n697) );
  NOR2_X1 U770 ( .A1(n695), .A2(G1961), .ZN(n696) );
  NOR2_X1 U771 ( .A1(n697), .A2(n696), .ZN(n704) );
  NOR2_X1 U772 ( .A1(G301), .A2(n704), .ZN(n698) );
  XNOR2_X1 U773 ( .A(n700), .B(n699), .ZN(n720) );
  NOR2_X1 U774 ( .A1(G1966), .A2(n740), .ZN(n722) );
  NOR2_X1 U775 ( .A1(G2084), .A2(n711), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n722), .A2(n718), .ZN(n701) );
  NAND2_X1 U777 ( .A1(G8), .A2(n701), .ZN(n702) );
  XNOR2_X1 U778 ( .A(KEYINPUT30), .B(n702), .ZN(n703) );
  NOR2_X1 U779 ( .A1(G168), .A2(n703), .ZN(n706) );
  AND2_X1 U780 ( .A1(G301), .A2(n704), .ZN(n705) );
  NOR2_X1 U781 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U782 ( .A(KEYINPUT31), .B(n707), .Z(n719) );
  NAND2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n708) );
  NAND2_X1 U784 ( .A1(n708), .A2(G286), .ZN(n710) );
  XNOR2_X1 U785 ( .A(n710), .B(n709), .ZN(n716) );
  NOR2_X1 U786 ( .A1(G1971), .A2(n740), .ZN(n713) );
  NOR2_X1 U787 ( .A1(G2090), .A2(n711), .ZN(n712) );
  NOR2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U789 ( .A1(G303), .A2(n714), .ZN(n715) );
  NAND2_X1 U790 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U791 ( .A1(G8), .A2(n718), .ZN(n724) );
  AND2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U795 ( .A1(G1976), .A2(G288), .ZN(n1028) );
  NOR2_X1 U796 ( .A1(G1971), .A2(G303), .ZN(n726) );
  NOR2_X1 U797 ( .A1(n1028), .A2(n726), .ZN(n727) );
  NAND2_X1 U798 ( .A1(G1976), .A2(G288), .ZN(n1029) );
  NAND2_X1 U799 ( .A1(n728), .A2(n1029), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n1028), .A2(KEYINPUT33), .ZN(n731) );
  NOR2_X1 U801 ( .A1(n731), .A2(n740), .ZN(n733) );
  XOR2_X1 U802 ( .A(G1981), .B(G305), .Z(n1011) );
  NOR2_X1 U803 ( .A1(G1981), .A2(G305), .ZN(n734) );
  XOR2_X1 U804 ( .A(n734), .B(KEYINPUT24), .Z(n735) );
  OR2_X1 U805 ( .A1(n740), .A2(n735), .ZN(n743) );
  NOR2_X1 U806 ( .A1(G2090), .A2(G303), .ZN(n736) );
  XOR2_X1 U807 ( .A(KEYINPUT103), .B(n736), .Z(n737) );
  NAND2_X1 U808 ( .A1(G8), .A2(n737), .ZN(n739) );
  NAND2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U810 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U811 ( .A(n745), .B(n744), .ZN(n780) );
  NAND2_X1 U812 ( .A1(G131), .A2(n921), .ZN(n748) );
  NAND2_X1 U813 ( .A1(G119), .A2(n926), .ZN(n747) );
  NAND2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n753) );
  NAND2_X1 U815 ( .A1(G95), .A2(n919), .ZN(n751) );
  BUF_X1 U816 ( .A(n749), .Z(n927) );
  NAND2_X1 U817 ( .A1(G107), .A2(n927), .ZN(n750) );
  NAND2_X1 U818 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X1 U819 ( .A1(n753), .A2(n752), .ZN(n937) );
  AND2_X1 U820 ( .A1(n937), .A2(G1991), .ZN(n763) );
  NAND2_X1 U821 ( .A1(G117), .A2(n927), .ZN(n754) );
  XNOR2_X1 U822 ( .A(n754), .B(KEYINPUT92), .ZN(n757) );
  NAND2_X1 U823 ( .A1(G105), .A2(n919), .ZN(n755) );
  XNOR2_X1 U824 ( .A(n755), .B(KEYINPUT38), .ZN(n756) );
  NAND2_X1 U825 ( .A1(n757), .A2(n756), .ZN(n761) );
  NAND2_X1 U826 ( .A1(G141), .A2(n921), .ZN(n759) );
  NAND2_X1 U827 ( .A1(G129), .A2(n926), .ZN(n758) );
  NAND2_X1 U828 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U829 ( .A1(n761), .A2(n760), .ZN(n940) );
  NOR2_X1 U830 ( .A1(n940), .A2(n781), .ZN(n762) );
  NOR2_X1 U831 ( .A1(n763), .A2(n762), .ZN(n972) );
  XOR2_X1 U832 ( .A(G1986), .B(G290), .Z(n1022) );
  NAND2_X1 U833 ( .A1(n972), .A2(n1022), .ZN(n768) );
  BUF_X1 U834 ( .A(n764), .Z(n766) );
  NOR2_X1 U835 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U836 ( .A(KEYINPUT90), .B(n767), .ZN(n794) );
  NAND2_X1 U837 ( .A1(n768), .A2(n794), .ZN(n779) );
  XNOR2_X1 U838 ( .A(G2067), .B(KEYINPUT37), .ZN(n791) );
  NAND2_X1 U839 ( .A1(G140), .A2(n921), .ZN(n770) );
  NAND2_X1 U840 ( .A1(G104), .A2(n919), .ZN(n769) );
  NAND2_X1 U841 ( .A1(n770), .A2(n769), .ZN(n772) );
  XOR2_X1 U842 ( .A(KEYINPUT91), .B(KEYINPUT34), .Z(n771) );
  XNOR2_X1 U843 ( .A(n772), .B(n771), .ZN(n777) );
  NAND2_X1 U844 ( .A1(G128), .A2(n926), .ZN(n774) );
  NAND2_X1 U845 ( .A1(G116), .A2(n927), .ZN(n773) );
  NAND2_X1 U846 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U847 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  NOR2_X1 U848 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U849 ( .A(KEYINPUT36), .B(n778), .ZN(n941) );
  NOR2_X1 U850 ( .A1(n791), .A2(n941), .ZN(n974) );
  NAND2_X1 U851 ( .A1(n974), .A2(n794), .ZN(n789) );
  NAND2_X1 U852 ( .A1(n780), .A2(n559), .ZN(n797) );
  AND2_X1 U853 ( .A1(n781), .A2(n940), .ZN(n782) );
  XOR2_X1 U854 ( .A(KEYINPUT105), .B(n782), .Z(n964) );
  INV_X1 U855 ( .A(n972), .ZN(n786) );
  NOR2_X1 U856 ( .A1(G1991), .A2(n937), .ZN(n783) );
  XNOR2_X1 U857 ( .A(KEYINPUT106), .B(n783), .ZN(n970) );
  NOR2_X1 U858 ( .A1(G1986), .A2(G290), .ZN(n784) );
  NOR2_X1 U859 ( .A1(n970), .A2(n784), .ZN(n785) );
  NOR2_X1 U860 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U861 ( .A1(n964), .A2(n787), .ZN(n788) );
  XNOR2_X1 U862 ( .A(n788), .B(KEYINPUT39), .ZN(n790) );
  NAND2_X1 U863 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U864 ( .A1(n791), .A2(n941), .ZN(n981) );
  NAND2_X1 U865 ( .A1(n792), .A2(n981), .ZN(n793) );
  XOR2_X1 U866 ( .A(KEYINPUT107), .B(n793), .Z(n795) );
  NAND2_X1 U867 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U868 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U869 ( .A(n798), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U870 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U871 ( .A1(G123), .A2(n926), .ZN(n799) );
  XNOR2_X1 U872 ( .A(n799), .B(KEYINPUT18), .ZN(n806) );
  NAND2_X1 U873 ( .A1(G135), .A2(n921), .ZN(n801) );
  NAND2_X1 U874 ( .A1(G111), .A2(n927), .ZN(n800) );
  NAND2_X1 U875 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U876 ( .A1(G99), .A2(n919), .ZN(n802) );
  XNOR2_X1 U877 ( .A(KEYINPUT79), .B(n802), .ZN(n803) );
  NOR2_X1 U878 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U879 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U880 ( .A(KEYINPUT80), .B(n807), .ZN(n967) );
  XNOR2_X1 U881 ( .A(n967), .B(G2096), .ZN(n808) );
  OR2_X1 U882 ( .A1(G2100), .A2(n808), .ZN(G156) );
  BUF_X1 U883 ( .A(n809), .Z(G164) );
  INV_X1 U884 ( .A(G57), .ZN(G237) );
  NAND2_X1 U885 ( .A1(G7), .A2(G661), .ZN(n810) );
  XNOR2_X1 U886 ( .A(n810), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U887 ( .A(G223), .ZN(n864) );
  NAND2_X1 U888 ( .A1(n864), .A2(G567), .ZN(n811) );
  XOR2_X1 U889 ( .A(KEYINPUT11), .B(n811), .Z(G234) );
  INV_X1 U890 ( .A(G860), .ZN(n819) );
  NOR2_X1 U891 ( .A1(n1018), .A2(n819), .ZN(n813) );
  XOR2_X1 U892 ( .A(KEYINPUT72), .B(n813), .Z(G153) );
  NAND2_X1 U893 ( .A1(G868), .A2(G301), .ZN(n815) );
  OR2_X1 U894 ( .A1(n1014), .A2(G868), .ZN(n814) );
  NAND2_X1 U895 ( .A1(n815), .A2(n814), .ZN(G284) );
  XOR2_X1 U896 ( .A(n1021), .B(KEYINPUT70), .Z(G299) );
  INV_X1 U897 ( .A(G868), .ZN(n816) );
  NOR2_X1 U898 ( .A1(G286), .A2(n816), .ZN(n818) );
  NOR2_X1 U899 ( .A1(G868), .A2(G299), .ZN(n817) );
  NOR2_X1 U900 ( .A1(n818), .A2(n817), .ZN(G297) );
  NAND2_X1 U901 ( .A1(n819), .A2(G559), .ZN(n820) );
  NAND2_X1 U902 ( .A1(n820), .A2(n1014), .ZN(n821) );
  XNOR2_X1 U903 ( .A(n821), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U904 ( .A1(G868), .A2(n1018), .ZN(n822) );
  XNOR2_X1 U905 ( .A(KEYINPUT78), .B(n822), .ZN(n825) );
  NAND2_X1 U906 ( .A1(G868), .A2(n1014), .ZN(n823) );
  NOR2_X1 U907 ( .A1(G559), .A2(n823), .ZN(n824) );
  NOR2_X1 U908 ( .A1(n825), .A2(n824), .ZN(G282) );
  NAND2_X1 U909 ( .A1(G80), .A2(n826), .ZN(n829) );
  NAND2_X1 U910 ( .A1(G93), .A2(n827), .ZN(n828) );
  NAND2_X1 U911 ( .A1(n829), .A2(n828), .ZN(n835) );
  NAND2_X1 U912 ( .A1(G67), .A2(n830), .ZN(n833) );
  NAND2_X1 U913 ( .A1(G55), .A2(n831), .ZN(n832) );
  NAND2_X1 U914 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U915 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U916 ( .A(KEYINPUT81), .B(n836), .Z(n871) );
  NOR2_X1 U917 ( .A1(n871), .A2(G868), .ZN(n837) );
  XNOR2_X1 U918 ( .A(KEYINPUT85), .B(n837), .ZN(n847) );
  XOR2_X1 U919 ( .A(G299), .B(KEYINPUT19), .Z(n839) );
  XNOR2_X1 U920 ( .A(G166), .B(n871), .ZN(n838) );
  XNOR2_X1 U921 ( .A(n839), .B(n838), .ZN(n842) );
  XNOR2_X1 U922 ( .A(G290), .B(G305), .ZN(n840) );
  XNOR2_X1 U923 ( .A(n840), .B(G288), .ZN(n841) );
  XNOR2_X1 U924 ( .A(n842), .B(n841), .ZN(n897) );
  NAND2_X1 U925 ( .A1(G559), .A2(n1014), .ZN(n843) );
  XNOR2_X1 U926 ( .A(n1018), .B(n843), .ZN(n870) );
  XNOR2_X1 U927 ( .A(n897), .B(n870), .ZN(n844) );
  NAND2_X1 U928 ( .A1(n844), .A2(G868), .ZN(n845) );
  XNOR2_X1 U929 ( .A(KEYINPUT84), .B(n845), .ZN(n846) );
  NAND2_X1 U930 ( .A1(n847), .A2(n846), .ZN(G295) );
  NAND2_X1 U931 ( .A1(G2084), .A2(G2078), .ZN(n848) );
  XOR2_X1 U932 ( .A(KEYINPUT20), .B(n848), .Z(n849) );
  NAND2_X1 U933 ( .A1(G2090), .A2(n849), .ZN(n850) );
  XNOR2_X1 U934 ( .A(KEYINPUT21), .B(n850), .ZN(n851) );
  NAND2_X1 U935 ( .A1(n851), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U936 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U937 ( .A1(G132), .A2(G82), .ZN(n852) );
  XNOR2_X1 U938 ( .A(n852), .B(KEYINPUT22), .ZN(n853) );
  XNOR2_X1 U939 ( .A(n853), .B(KEYINPUT86), .ZN(n854) );
  NOR2_X1 U940 ( .A1(G218), .A2(n854), .ZN(n855) );
  NAND2_X1 U941 ( .A1(G96), .A2(n855), .ZN(n868) );
  NAND2_X1 U942 ( .A1(n868), .A2(G2106), .ZN(n859) );
  NAND2_X1 U943 ( .A1(G69), .A2(G120), .ZN(n856) );
  NOR2_X1 U944 ( .A1(G237), .A2(n856), .ZN(n857) );
  NAND2_X1 U945 ( .A1(G108), .A2(n857), .ZN(n869) );
  NAND2_X1 U946 ( .A1(n869), .A2(G567), .ZN(n858) );
  NAND2_X1 U947 ( .A1(n859), .A2(n858), .ZN(n873) );
  NAND2_X1 U948 ( .A1(G661), .A2(G483), .ZN(n860) );
  NOR2_X1 U949 ( .A1(n873), .A2(n860), .ZN(n867) );
  NAND2_X1 U950 ( .A1(n867), .A2(G36), .ZN(n861) );
  XOR2_X1 U951 ( .A(KEYINPUT87), .B(n861), .Z(G176) );
  NOR2_X1 U952 ( .A1(n863), .A2(n862), .ZN(G160) );
  NAND2_X1 U953 ( .A1(G2106), .A2(n864), .ZN(G217) );
  AND2_X1 U954 ( .A1(G15), .A2(G2), .ZN(n865) );
  NAND2_X1 U955 ( .A1(G661), .A2(n865), .ZN(G259) );
  NAND2_X1 U956 ( .A1(G3), .A2(G1), .ZN(n866) );
  NAND2_X1 U957 ( .A1(n867), .A2(n866), .ZN(G188) );
  NOR2_X1 U958 ( .A1(n869), .A2(n868), .ZN(G325) );
  XOR2_X1 U959 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U961 ( .A(G132), .ZN(G219) );
  INV_X1 U962 ( .A(G120), .ZN(G236) );
  INV_X1 U963 ( .A(G82), .ZN(G220) );
  INV_X1 U964 ( .A(G69), .ZN(G235) );
  NOR2_X1 U965 ( .A1(n870), .A2(G860), .ZN(n872) );
  XNOR2_X1 U966 ( .A(n872), .B(n871), .ZN(G145) );
  INV_X1 U967 ( .A(n873), .ZN(G319) );
  XNOR2_X1 U968 ( .A(G2078), .B(G2072), .ZN(n874) );
  XNOR2_X1 U969 ( .A(n874), .B(KEYINPUT42), .ZN(n884) );
  XOR2_X1 U970 ( .A(KEYINPUT43), .B(G2100), .Z(n876) );
  XNOR2_X1 U971 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n876), .B(n875), .ZN(n880) );
  XOR2_X1 U973 ( .A(G2096), .B(G2090), .Z(n878) );
  XNOR2_X1 U974 ( .A(G2067), .B(G2084), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U976 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U977 ( .A(G2678), .B(KEYINPUT111), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(G227) );
  XOR2_X1 U980 ( .A(G1971), .B(G1961), .Z(n886) );
  XNOR2_X1 U981 ( .A(G1996), .B(G1991), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n896) );
  XOR2_X1 U983 ( .A(KEYINPUT114), .B(KEYINPUT112), .Z(n888) );
  XNOR2_X1 U984 ( .A(G1956), .B(G2474), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U986 ( .A(G1976), .B(G1981), .Z(n890) );
  XNOR2_X1 U987 ( .A(G1986), .B(G1966), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U989 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U990 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(G229) );
  INV_X1 U993 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U994 ( .A(n897), .B(KEYINPUT121), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n1018), .B(G286), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n1014), .B(G171), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G397) );
  NAND2_X1 U1000 ( .A1(G124), .A2(n926), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n903), .B(KEYINPUT44), .ZN(n908) );
  NAND2_X1 U1002 ( .A1(G100), .A2(n919), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G112), .A2(n927), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(KEYINPUT116), .B(n906), .Z(n907) );
  NAND2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(G136), .A2(n921), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT115), .B(n909), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(G162) );
  XOR2_X1 U1010 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n935) );
  NAND2_X1 U1011 ( .A1(G139), .A2(n921), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(G103), .A2(n919), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n918) );
  NAND2_X1 U1014 ( .A1(G127), .A2(n926), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(G115), .A2(n927), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1017 ( .A(KEYINPUT47), .B(n916), .Z(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n977) );
  XNOR2_X1 U1019 ( .A(KEYINPUT45), .B(KEYINPUT119), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(n919), .A2(G106), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n920), .B(KEYINPUT118), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(G142), .A2(n921), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n925), .B(n924), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(G130), .A2(n926), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(G118), .A2(n927), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT117), .B(n930), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n977), .B(n933), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(n935), .B(n934), .ZN(n936) );
  XOR2_X1 U1032 ( .A(n936), .B(n967), .Z(n939) );
  XOR2_X1 U1033 ( .A(n937), .B(G162), .Z(n938) );
  XNOR2_X1 U1034 ( .A(n939), .B(n938), .ZN(n945) );
  XNOR2_X1 U1035 ( .A(n941), .B(n940), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(G164), .B(G160), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n943), .B(n942), .ZN(n944) );
  XOR2_X1 U1038 ( .A(n945), .B(n944), .Z(n946) );
  NOR2_X1 U1039 ( .A1(G37), .A2(n946), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT120), .B(n947), .ZN(G395) );
  XOR2_X1 U1041 ( .A(G2451), .B(G2430), .Z(n949) );
  XNOR2_X1 U1042 ( .A(G2438), .B(G2443), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n949), .B(n948), .ZN(n955) );
  XOR2_X1 U1044 ( .A(G2435), .B(G2454), .Z(n951) );
  XNOR2_X1 U1045 ( .A(G1348), .B(G1341), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(n951), .B(n950), .ZN(n953) );
  XOR2_X1 U1047 ( .A(G2446), .B(G2427), .Z(n952) );
  XNOR2_X1 U1048 ( .A(n953), .B(n952), .ZN(n954) );
  XOR2_X1 U1049 ( .A(n955), .B(n954), .Z(n956) );
  NAND2_X1 U1050 ( .A1(G14), .A2(n956), .ZN(n962) );
  NAND2_X1 U1051 ( .A1(G319), .A2(n962), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(G227), .A2(G229), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(KEYINPUT49), .B(n957), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(G397), .A2(G395), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(G225) );
  INV_X1 U1057 ( .A(G225), .ZN(G308) );
  INV_X1 U1058 ( .A(G96), .ZN(G221) );
  INV_X1 U1059 ( .A(G108), .ZN(G238) );
  INV_X1 U1060 ( .A(n962), .ZN(G401) );
  XOR2_X1 U1061 ( .A(G2090), .B(G162), .Z(n963) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1063 ( .A(KEYINPUT122), .B(n965), .Z(n966) );
  XNOR2_X1 U1064 ( .A(KEYINPUT51), .B(n966), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G160), .B(G2084), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n984) );
  XOR2_X1 U1071 ( .A(G2072), .B(n977), .Z(n979) );
  XOR2_X1 U1072 ( .A(G164), .B(G2078), .Z(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n980), .B(KEYINPUT50), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n985), .ZN(n986) );
  INV_X1 U1078 ( .A(KEYINPUT55), .ZN(n1007) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n1007), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n987), .A2(G29), .ZN(n1067) );
  XNOR2_X1 U1081 ( .A(G2090), .B(G35), .ZN(n1002) );
  XNOR2_X1 U1082 ( .A(G2067), .B(G26), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G33), .B(G2072), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n990), .B(G27), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(G32), .B(G1996), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G1991), .B(G25), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(n995), .B(KEYINPUT123), .ZN(n996) );
  NAND2_X1 U1091 ( .A1(G28), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1092 ( .A(KEYINPUT124), .B(n997), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1094 ( .A(KEYINPUT53), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(G2084), .B(G34), .Z(n1003) );
  XNOR2_X1 U1097 ( .A(KEYINPUT54), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1099 ( .A(n1007), .B(n1006), .ZN(n1009) );
  INV_X1 U1100 ( .A(G29), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1010), .ZN(n1065) );
  XNOR2_X1 U1103 ( .A(G16), .B(KEYINPUT56), .ZN(n1037) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G168), .ZN(n1012) );
  NAND2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1106 ( .A(n1013), .B(KEYINPUT57), .ZN(n1035) );
  XNOR2_X1 U1107 ( .A(G1348), .B(n1014), .ZN(n1016) );
  XNOR2_X1 U1108 ( .A(G171), .B(G1961), .ZN(n1015) );
  NAND2_X1 U1109 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1110 ( .A(KEYINPUT125), .B(n1017), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(n1018), .B(G1341), .Z(n1020) );
  XNOR2_X1 U1112 ( .A(G166), .B(G1971), .ZN(n1019) );
  NAND2_X1 U1113 ( .A1(n1020), .A2(n1019), .ZN(n1025) );
  XNOR2_X1 U1114 ( .A(n1021), .B(G1956), .ZN(n1023) );
  NAND2_X1 U1115 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1033) );
  INV_X1 U1118 ( .A(n1028), .ZN(n1030) );
  NAND2_X1 U1119 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1120 ( .A(KEYINPUT126), .B(n1031), .ZN(n1032) );
  NOR2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1063) );
  INV_X1 U1124 ( .A(G16), .ZN(n1061) );
  XOR2_X1 U1125 ( .A(G1976), .B(G23), .Z(n1039) );
  XOR2_X1 U1126 ( .A(G1971), .B(G22), .Z(n1038) );
  NAND2_X1 U1127 ( .A1(n1039), .A2(n1038), .ZN(n1041) );
  XNOR2_X1 U1128 ( .A(G24), .B(G1986), .ZN(n1040) );
  NOR2_X1 U1129 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XOR2_X1 U1130 ( .A(KEYINPUT58), .B(n1042), .Z(n1058) );
  XOR2_X1 U1131 ( .A(G1961), .B(G5), .Z(n1053) );
  XNOR2_X1 U1132 ( .A(G20), .B(n1043), .ZN(n1047) );
  XNOR2_X1 U1133 ( .A(G1341), .B(G19), .ZN(n1045) );
  XNOR2_X1 U1134 ( .A(G6), .B(G1981), .ZN(n1044) );
  NOR2_X1 U1135 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1136 ( .A1(n1047), .A2(n1046), .ZN(n1050) );
  XOR2_X1 U1137 ( .A(KEYINPUT59), .B(G1348), .Z(n1048) );
  XNOR2_X1 U1138 ( .A(G4), .B(n1048), .ZN(n1049) );
  NOR2_X1 U1139 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XNOR2_X1 U1140 ( .A(KEYINPUT60), .B(n1051), .ZN(n1052) );
  NAND2_X1 U1141 ( .A1(n1053), .A2(n1052), .ZN(n1055) );
  XNOR2_X1 U1142 ( .A(G21), .B(G1966), .ZN(n1054) );
  NOR2_X1 U1143 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  XNOR2_X1 U1144 ( .A(KEYINPUT127), .B(n1056), .ZN(n1057) );
  NOR2_X1 U1145 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  XNOR2_X1 U1146 ( .A(KEYINPUT61), .B(n1059), .ZN(n1060) );
  NAND2_X1 U1147 ( .A1(n1061), .A2(n1060), .ZN(n1062) );
  NAND2_X1 U1148 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
  NOR2_X1 U1149 ( .A1(n1065), .A2(n1064), .ZN(n1066) );
  NAND2_X1 U1150 ( .A1(n1067), .A2(n1066), .ZN(n1068) );
  XOR2_X1 U1151 ( .A(KEYINPUT62), .B(n1068), .Z(G311) );
  INV_X1 U1152 ( .A(G311), .ZN(G150) );
endmodule

