//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G101), .ZN(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n188), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G119), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT66), .A3(G116), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(G119), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT2), .B(G113), .Z(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT71), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT65), .A3(new_n208), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n211), .B2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n215), .A2(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  INV_X1    g036(.A(G134), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G137), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(G134), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n222), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT11), .B1(new_n226), .B2(G134), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n229), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n224), .A2(G137), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT11), .A2(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n232), .A2(new_n236), .A3(new_n222), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT67), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(G134), .B1(new_n233), .B2(new_n234), .ZN(new_n239));
  INV_X1    g053(.A(new_n229), .ZN(new_n240));
  OAI21_X1  g054(.A(G131), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n232), .A2(new_n236), .A3(new_n222), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n221), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n222), .B1(new_n232), .B2(new_n236), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n250), .A2(new_n216), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n216), .A2(new_n249), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n247), .A2(new_n243), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n206), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n215), .A2(new_n217), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n218), .A2(new_n220), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n242), .B1(new_n241), .B2(new_n243), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n252), .B1(new_n250), .B2(new_n216), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n237), .B2(new_n246), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(KEYINPUT71), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n205), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n196), .B1(new_n264), .B2(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(new_n205), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n245), .A2(new_n206), .A3(new_n253), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n260), .B2(new_n262), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n241), .A2(new_n243), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n262), .B1(new_n221), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n205), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n205), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n260), .A2(new_n266), .A3(new_n262), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n260), .A2(new_n283), .A3(new_n266), .A4(new_n262), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n270), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n195), .B1(new_n272), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n260), .B2(new_n262), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n274), .A2(KEYINPUT30), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n205), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n194), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT31), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n285), .A2(new_n291), .A3(KEYINPUT31), .A4(new_n194), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n287), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n287), .A2(new_n299), .A3(new_n296), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n187), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n279), .B1(new_n284), .B2(new_n282), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n265), .B(new_n271), .C1(new_n304), .C2(new_n270), .ZN(new_n305));
  AOI221_X4 g119(.A(KEYINPUT73), .B1(new_n294), .B2(new_n295), .C1(new_n305), .C2(new_n195), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n299), .B1(new_n287), .B2(new_n296), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n187), .B(new_n302), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n272), .A2(new_n286), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n194), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT74), .B1(new_n305), .B2(new_n195), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n285), .A2(new_n291), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n195), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n205), .B1(new_n245), .B2(new_n253), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n285), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(new_n270), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(new_n272), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n195), .A2(new_n313), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G472), .ZN(new_n326));
  OAI22_X1  g140(.A1(new_n303), .A2(new_n309), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT75), .B(G217), .ZN(new_n328));
  INV_X1    g142(.A(G902), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(G234), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G902), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n207), .A2(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n200), .A2(G128), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT24), .B(G110), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n333), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n332), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n336), .B1(new_n341), .B2(G110), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT76), .B(G140), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G140), .ZN(new_n348));
  INV_X1    g162(.A(G140), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(KEYINPUT76), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT77), .B(G125), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(KEYINPUT78), .A2(G125), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT78), .A2(G125), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(G140), .A3(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n351), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT16), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n349), .ZN(new_n358));
  AOI21_X1  g172(.A(G146), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n359), .A2(KEYINPUT79), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(G146), .A3(new_n358), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n359), .B2(KEYINPUT79), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n342), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(G125), .B(G140), .Z(new_n364));
  NOR2_X1   g178(.A1(new_n341), .A2(G110), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n334), .A2(new_n335), .ZN(new_n366));
  OAI221_X1 g180(.A(new_n361), .B1(G146), .B2(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G137), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n363), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n363), .B2(new_n367), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n374), .A2(KEYINPUT81), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(KEYINPUT81), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n331), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n329), .B1(new_n372), .B2(new_n373), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n363), .A2(new_n367), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n370), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n363), .A2(new_n367), .A3(new_n371), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT25), .A3(new_n329), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n380), .A2(new_n385), .A3(KEYINPUT80), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n330), .B1(new_n380), .B2(KEYINPUT80), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n377), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n203), .A2(KEYINPUT5), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n198), .A2(KEYINPUT5), .A3(G119), .ZN(new_n391));
  INV_X1    g205(.A(G113), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n203), .A2(new_n204), .ZN(new_n395));
  INV_X1    g209(.A(G101), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G104), .ZN(new_n398));
  INV_X1    g212(.A(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n397), .B2(G104), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(new_n399), .B2(G107), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n397), .A3(G104), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(KEYINPUT83), .A3(G107), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n404), .A2(new_n405), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n402), .B1(new_n409), .B2(G101), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n394), .A2(new_n395), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G122), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT8), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n393), .B1(new_n390), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT89), .B1(new_n203), .B2(KEYINPUT5), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n395), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n410), .B1(new_n418), .B2(KEYINPUT90), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n395), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n257), .A2(new_n352), .A3(new_n353), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n261), .A2(new_n356), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT88), .B(G224), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n190), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(KEYINPUT7), .A3(new_n428), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n404), .A2(new_n405), .A3(new_n407), .A4(new_n408), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n396), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n409), .A2(G101), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(KEYINPUT4), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n409), .A2(new_n434), .A3(G101), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n205), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n401), .B1(new_n430), .B2(new_n396), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n394), .A2(new_n437), .A3(new_n395), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n438), .A3(new_n412), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n428), .A2(KEYINPUT7), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n424), .A2(new_n425), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n429), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n423), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n436), .A2(new_n438), .ZN(new_n446));
  INV_X1    g260(.A(new_n412), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n426), .B(new_n428), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n451), .A3(new_n447), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n444), .A2(new_n445), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n445), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n329), .B1(new_n422), .B2(new_n442), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G214), .B1(G237), .B2(G902), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT91), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT9), .B(G234), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n257), .A2(KEYINPUT10), .A3(new_n437), .ZN(new_n467));
  INV_X1    g281(.A(new_n432), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT4), .B1(new_n409), .B2(G101), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n261), .B(new_n435), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT84), .B(KEYINPUT1), .C1(new_n211), .C2(G146), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT84), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n474));
  OAI21_X1  g288(.A(G128), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n218), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n410), .B1(new_n476), .B2(new_n255), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT85), .B1(new_n477), .B2(KEYINPUT10), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n219), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n207), .B1(new_n480), .B2(new_n472), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT65), .B1(new_n216), .B2(new_n208), .ZN(new_n482));
  AND4_X1   g296(.A1(KEYINPUT65), .A2(new_n208), .A3(new_n210), .A4(new_n212), .ZN(new_n483));
  OAI22_X1  g297(.A1(new_n481), .A2(new_n216), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n437), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT10), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n471), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n247), .A2(new_n243), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n466), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n467), .A2(new_n470), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n486), .B1(new_n485), .B2(new_n487), .ZN(new_n494));
  AOI211_X1 g308(.A(KEYINPUT85), .B(KEYINPUT10), .C1(new_n484), .C2(new_n437), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT86), .A3(new_n490), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n492), .A2(new_n497), .B1(new_n491), .B2(new_n489), .ZN(new_n498));
  XOR2_X1   g312(.A(G110), .B(G140), .Z(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT82), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n190), .A2(G227), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT87), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n489), .A2(new_n491), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n489), .A2(new_n466), .A3(new_n491), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT86), .B1(new_n496), .B2(new_n490), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n508));
  INV_X1    g322(.A(new_n502), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n257), .A2(new_n437), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n490), .B1(new_n477), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT12), .Z(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n489), .B2(new_n491), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n503), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G469), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n329), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n502), .B1(new_n513), .B2(new_n504), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n492), .A2(new_n497), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(new_n514), .ZN(new_n521));
  OAI21_X1  g335(.A(G469), .B1(new_n521), .B2(G902), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n465), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n360), .A2(new_n362), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n189), .A2(new_n190), .A3(G214), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(G143), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n222), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n527), .A2(new_n222), .ZN(new_n529));
  MUX2_X1   g343(.A(new_n528), .B(new_n529), .S(KEYINPUT17), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G113), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(new_n399), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n527), .B1(new_n534), .B2(new_n222), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n346), .A2(new_n351), .A3(new_n354), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n209), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n364), .A2(G146), .ZN(new_n538));
  OAI221_X1 g352(.A(new_n535), .B1(new_n534), .B2(new_n529), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(KEYINPUT19), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT19), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n364), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n209), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n361), .A3(new_n528), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n539), .ZN(new_n547));
  INV_X1    g361(.A(new_n533), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G475), .A2(G902), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n524), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n551), .ZN(new_n553));
  AOI211_X1 g367(.A(KEYINPUT20), .B(new_n553), .C1(new_n540), .C2(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n531), .A2(new_n539), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n548), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n556), .B2(new_n540), .ZN(new_n557));
  INV_X1    g371(.A(G475), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n552), .A2(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n207), .A2(G143), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n211), .A2(G128), .ZN(new_n561));
  OAI21_X1  g375(.A(G134), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n560), .ZN(new_n563));
  INV_X1    g377(.A(new_n561), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n223), .ZN(new_n565));
  INV_X1    g379(.A(G122), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G116), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n198), .A2(G122), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n562), .A2(new_n565), .B1(new_n569), .B2(new_n397), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n198), .A2(G122), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n568), .B1(new_n571), .B2(KEYINPUT14), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(KEYINPUT14), .B2(new_n568), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n573), .A2(new_n574), .A3(G107), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n573), .B2(G107), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n569), .B(new_n397), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n560), .B1(new_n564), .B2(KEYINPUT13), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n560), .A2(KEYINPUT13), .ZN(new_n580));
  OAI21_X1  g394(.A(G134), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n581), .A3(new_n565), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n328), .A2(new_n463), .A3(G953), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n329), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G478), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT15), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n590), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n585), .A2(new_n329), .A3(new_n587), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT21), .B(G898), .Z(new_n595));
  NAND2_X1  g409(.A1(G234), .A2(G237), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(G902), .A3(G953), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n190), .A2(G952), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n596), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n559), .A2(new_n594), .A3(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n462), .A2(new_n523), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n327), .A2(new_n389), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT93), .B(G101), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G3));
  OAI21_X1  g421(.A(new_n329), .B1(new_n306), .B2(new_n307), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G472), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n610));
  AND4_X1   g424(.A1(new_n389), .A2(new_n609), .A3(new_n610), .A4(new_n523), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n588), .A2(new_n589), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n583), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n583), .B2(new_n614), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n616), .A2(KEYINPUT95), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(KEYINPUT95), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n585), .A2(new_n613), .A3(new_n587), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n589), .A2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n612), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n559), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n624), .A2(new_n602), .A3(new_n461), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n611), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT96), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT34), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G104), .ZN(G6));
  INV_X1    g443(.A(new_n559), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n594), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n601), .B(KEYINPUT97), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n631), .A2(new_n461), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n611), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(new_n330), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT25), .B1(new_n384), .B2(new_n329), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT80), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n380), .A2(new_n385), .A3(KEYINPUT80), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n371), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n381), .B(new_n643), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n641), .A2(new_n642), .B1(new_n331), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n298), .B2(new_n300), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n610), .B(new_n646), .C1(new_n647), .C2(new_n326), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n604), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  XOR2_X1   g466(.A(new_n600), .B(KEYINPUT99), .Z(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT98), .B(G900), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n653), .B1(new_n597), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n645), .A2(new_n461), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n327), .A2(new_n523), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XOR2_X1   g474(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n655), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n523), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT101), .Z(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT40), .Z(new_n665));
  INV_X1    g479(.A(new_n292), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n195), .B2(new_n319), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n667), .B2(G902), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n303), .B2(new_n309), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n459), .B(KEYINPUT38), .Z(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n559), .A2(new_n594), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n460), .A3(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n670), .A2(new_n646), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NOR2_X1   g491(.A1(new_n624), .A2(new_n656), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n327), .A2(new_n523), .A3(new_n658), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  AOI21_X1  g494(.A(new_n326), .B1(new_n317), .B2(new_n324), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n610), .A2(KEYINPUT32), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n681), .B1(new_n682), .B2(new_n308), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n388), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n516), .A2(new_n329), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n518), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n465), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n625), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND4_X1  g505(.A1(new_n327), .A2(new_n389), .A3(new_n634), .A4(new_n688), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NAND4_X1  g507(.A1(new_n327), .A2(new_n603), .A3(new_n658), .A4(new_n688), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  OAI21_X1  g509(.A(new_n195), .B1(new_n321), .B2(new_n272), .ZN(new_n696));
  AOI211_X1 g510(.A(G472), .B(G902), .C1(new_n696), .C2(new_n296), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n388), .B(new_n697), .C1(new_n608), .C2(G472), .ZN(new_n698));
  INV_X1    g512(.A(new_n460), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n454), .B2(new_n458), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n559), .A2(new_n700), .A3(new_n594), .A4(new_n632), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n687), .A2(new_n465), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  AOI211_X1 g518(.A(new_n645), .B(new_n697), .C1(new_n608), .C2(G472), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n686), .A2(new_n464), .A3(new_n518), .A4(new_n700), .ZN(new_n706));
  INV_X1    g520(.A(new_n624), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n655), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n705), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n516), .A2(new_n517), .A3(new_n329), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n517), .B1(new_n516), .B2(new_n329), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n464), .A3(new_n700), .A4(new_n678), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n696), .A2(new_n296), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n302), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n646), .B(new_n717), .C1(new_n647), .C2(new_n326), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT102), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  NAND2_X1  g535(.A1(new_n518), .A2(new_n522), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n459), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n460), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n465), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n518), .A2(KEYINPUT103), .A3(new_n522), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n678), .A2(new_n730), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n683), .A2(new_n729), .A3(new_n388), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n327), .A2(KEYINPUT104), .A3(new_n389), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n683), .B2(new_n388), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n729), .A2(new_n708), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n732), .B1(new_n737), .B2(KEYINPUT42), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  AND2_X1   g553(.A1(new_n724), .A2(new_n728), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n684), .A2(new_n657), .A3(new_n727), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  NAND2_X1  g556(.A1(new_n630), .A2(new_n623), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT43), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n645), .B(new_n744), .C1(new_n610), .C2(new_n609), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n726), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n746), .B1(new_n753), .B2(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g568(.A1(G469), .A2(G902), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n521), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(G469), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT105), .B1(new_n757), .B2(G469), .ZN(new_n761));
  OAI211_X1 g575(.A(KEYINPUT46), .B(new_n755), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT106), .A3(new_n518), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n758), .B(new_n759), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n755), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n763), .B1(new_n765), .B2(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT106), .B1(new_n762), .B2(new_n518), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n464), .B(new_n662), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n752), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n754), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  OAI21_X1  g586(.A(new_n464), .B1(new_n766), .B2(new_n767), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT47), .B(new_n464), .C1(new_n766), .C2(new_n767), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n683), .A2(new_n388), .A3(new_n678), .A4(new_n750), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT109), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT110), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n349), .ZN(G42));
  XNOR2_X1  g597(.A(new_n714), .B(KEYINPUT49), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n671), .A2(new_n464), .A3(new_n460), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n388), .A3(new_n743), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n670), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n744), .A2(new_n653), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n698), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n688), .A2(new_n699), .A3(new_n671), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT50), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n669), .A2(new_n388), .A3(new_n600), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n714), .A2(new_n727), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT116), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n623), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n630), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n795), .A2(new_n800), .A3(new_n788), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n800), .B1(new_n795), .B2(new_n788), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT118), .B1(new_n803), .B2(new_n718), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n803), .A2(KEYINPUT118), .A3(new_n718), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n714), .A2(new_n465), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n775), .A2(new_n776), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n789), .A2(new_n726), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT114), .Z(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n599), .B1(new_n789), .B2(new_n706), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n707), .B2(new_n796), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n733), .A2(new_n735), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(KEYINPUT48), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(KEYINPUT48), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n812), .B(new_n814), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n807), .B(KEYINPUT115), .Z(new_n820));
  OAI21_X1  g634(.A(new_n810), .B1(new_n777), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT51), .B1(new_n806), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n673), .A2(new_n700), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n823), .A2(new_n646), .A3(new_n465), .A4(new_n656), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n669), .A3(new_n740), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n720), .A2(new_n659), .A3(new_n679), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n658), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n683), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n830), .B(new_n523), .C1(new_n657), .C2(new_n678), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n720), .A4(new_n825), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n834));
  INV_X1    g648(.A(new_n732), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n834), .A2(new_n835), .A3(new_n741), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n605), .A2(new_n650), .A3(new_n703), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n688), .A2(new_n603), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n462), .A2(new_n632), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n591), .A2(new_n841), .A3(new_n593), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n591), .B2(new_n593), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n624), .A2(new_n840), .B1(new_n630), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n707), .A2(KEYINPUT111), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n839), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n830), .A2(new_n838), .B1(new_n847), .B2(new_n611), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n609), .A2(new_n717), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n729), .A2(new_n849), .A3(new_n708), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n556), .A2(new_n540), .ZN(new_n851));
  OAI21_X1  g665(.A(G475), .B1(new_n851), .B2(G902), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n842), .A2(new_n843), .A3(new_n656), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n852), .B(new_n853), .C1(new_n552), .C2(new_n554), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n726), .B1(new_n854), .B2(KEYINPUT113), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(new_n523), .C1(KEYINPUT113), .C2(new_n854), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n683), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n646), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n684), .B(new_n688), .C1(new_n625), .C2(new_n634), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n837), .A2(new_n848), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(KEYINPUT53), .A2(new_n833), .A3(new_n836), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n834), .A2(new_n835), .A3(new_n741), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n860), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n864), .B2(new_n833), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  INV_X1    g681(.A(new_n833), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n604), .A2(new_n649), .B1(new_n698), .B2(new_n702), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n847), .A2(new_n611), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n694), .A4(new_n605), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n689), .A2(new_n692), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n738), .A3(new_n741), .A4(new_n858), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n867), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n833), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n866), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n819), .A2(new_n822), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n787), .B1(new_n880), .B2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n190), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n329), .B1(new_n875), .B2(new_n877), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(G210), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n449), .A2(new_n452), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n450), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n456), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n884), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n885), .B(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n455), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n897), .B2(new_n891), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n892), .B1(new_n896), .B2(new_n900), .ZN(G51));
  AND2_X1   g715(.A1(new_n885), .A2(new_n893), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n885), .A2(new_n893), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n764), .ZN(new_n904));
  INV_X1    g718(.A(new_n516), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n866), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n875), .A2(new_n877), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(KEYINPUT122), .A3(KEYINPUT54), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n878), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n755), .B(KEYINPUT57), .Z(new_n911));
  AOI21_X1  g725(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n904), .B1(new_n912), .B2(KEYINPUT123), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n878), .B1(new_n914), .B2(KEYINPUT122), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n866), .A2(new_n906), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n516), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n883), .B1(new_n913), .B2(new_n920), .ZN(G54));
  NAND4_X1  g735(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .A4(new_n550), .ZN(new_n922));
  NAND2_X1  g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n540), .B(new_n549), .C1(new_n894), .C2(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n922), .A2(new_n924), .A3(new_n884), .ZN(G60));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n926));
  INV_X1    g740(.A(new_n620), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n910), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n866), .B2(new_n878), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n884), .B1(new_n932), .B2(new_n927), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n910), .A2(new_n927), .A3(new_n930), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n932), .A2(new_n927), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT124), .A4(new_n884), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n875), .B2(new_n877), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n644), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n375), .A2(new_n376), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n942), .B(new_n884), .C1(new_n943), .C2(new_n941), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT61), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G66));
  AOI21_X1  g761(.A(new_n190), .B1(new_n595), .B2(new_n427), .ZN(new_n948));
  INV_X1    g762(.A(new_n873), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n190), .ZN(new_n950));
  INV_X1    g764(.A(G898), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n887), .B1(new_n951), .B2(G953), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n950), .B(new_n952), .ZN(G69));
  AOI21_X1  g767(.A(new_n726), .B1(new_n845), .B2(new_n846), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n684), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n664), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n754), .B2(new_n770), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n831), .A2(new_n720), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n665), .B2(new_n675), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n957), .B(new_n960), .C1(new_n781), .C2(new_n780), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n190), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n289), .A2(new_n290), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n544), .B(KEYINPUT126), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n768), .A2(new_n815), .A3(new_n823), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(new_n958), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n771), .A2(new_n836), .A3(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n972), .A2(new_n782), .A3(G953), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n967), .B(new_n969), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n973), .A2(new_n975), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n965), .B1(new_n961), .B2(new_n190), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n968), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(G72));
  XOR2_X1   g794(.A(new_n315), .B(KEYINPUT127), .Z(new_n981));
  NOR3_X1   g795(.A1(new_n972), .A2(new_n782), .A3(new_n949), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n195), .B(new_n981), .C1(new_n982), .C2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n961), .B2(new_n949), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n981), .A2(new_n195), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n985), .B1(new_n316), .B2(new_n292), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n883), .B1(new_n908), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n986), .A2(new_n989), .A3(new_n991), .ZN(G57));
endmodule


