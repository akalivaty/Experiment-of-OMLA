//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n192), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G107), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n202), .A2(KEYINPUT3), .A3(G104), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT3), .B1(new_n202), .B2(G104), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n199), .B(new_n201), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT4), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n202), .A2(G104), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n200), .B2(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(KEYINPUT3), .A3(G104), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g027(.A(KEYINPUT73), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n206), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT73), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(new_n212), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n217), .A2(KEYINPUT4), .A3(new_n218), .A4(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT74), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n202), .B2(G104), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n202), .A2(G104), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n200), .A2(KEYINPUT74), .A3(G107), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n237), .A2(new_n205), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  OAI22_X1  g054(.A1(new_n240), .A2(new_n224), .B1(new_n222), .B2(G128), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT64), .B1(new_n228), .B2(new_n240), .ZN(new_n243));
  AND4_X1   g057(.A1(KEYINPUT64), .A2(new_n240), .A3(new_n222), .A4(new_n224), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT10), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n238), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n240), .A2(new_n222), .A3(new_n224), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n228), .A2(KEYINPUT64), .A3(new_n240), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n241), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n237), .A2(new_n205), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT10), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n220), .A2(new_n231), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n198), .B1(new_n255), .B2(KEYINPUT77), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n220), .A2(new_n231), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n254), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n257), .A2(KEYINPUT77), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT78), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n258), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT77), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n255), .A2(KEYINPUT77), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT78), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .A4(new_n198), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n198), .B(KEYINPUT75), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G110), .B(G140), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n272), .A2(G227), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n271), .B(new_n273), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n252), .B(new_n253), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(new_n198), .B1(KEYINPUT76), .B2(KEYINPUT12), .ZN(new_n279));
  OR2_X1    g093(.A1(KEYINPUT76), .A2(KEYINPUT12), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n275), .B1(new_n281), .B2(new_n270), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n187), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT79), .B(G469), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n274), .B1(new_n267), .B2(new_n269), .ZN(new_n287));
  INV_X1    g101(.A(new_n276), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(new_n281), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n284), .B(new_n286), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT80), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n270), .B1(new_n260), .B2(new_n266), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n292), .A2(new_n274), .B1(new_n288), .B2(new_n281), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT80), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n284), .A4(new_n286), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n285), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G214), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n231), .A2(G125), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n252), .B2(G125), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT81), .B(G224), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G953), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n300), .B(new_n303), .C1(new_n252), .C2(G125), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n305), .A2(KEYINPUT82), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT82), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT2), .B(G113), .Z(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G116), .B(G119), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(KEYINPUT65), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n220), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(KEYINPUT5), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G116), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n316), .B(G113), .C1(KEYINPUT5), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n310), .A2(new_n312), .ZN(new_n320));
  AND4_X1   g134(.A1(new_n205), .A2(new_n319), .A3(new_n237), .A4(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G110), .B(G122), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n323), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n313), .B(new_n310), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n215), .B2(new_n219), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n327), .B2(new_n321), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n328), .A3(KEYINPUT6), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT6), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n330), .B(new_n325), .C1(new_n327), .C2(new_n321), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n309), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n323), .B(KEYINPUT8), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n319), .A2(new_n320), .B1(new_n237), .B2(new_n205), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n321), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n301), .A2(KEYINPUT7), .A3(new_n304), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT7), .ZN(new_n337));
  OAI221_X1 g151(.A(new_n300), .B1(new_n337), .B2(new_n303), .C1(new_n252), .C2(G125), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(G902), .B1(new_n339), .B2(new_n324), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n299), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n332), .A2(new_n340), .A3(new_n299), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n298), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G221), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT9), .B(G234), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n348), .B2(new_n284), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n296), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT16), .ZN(new_n351));
  INV_X1    g165(.A(G140), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G125), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(G125), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n353), .B1(new_n357), .B2(new_n351), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n221), .ZN(new_n359));
  OAI211_X1 g173(.A(G146), .B(new_n353), .C1(new_n357), .C2(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G110), .ZN(new_n362));
  OR3_X1    g176(.A1(new_n317), .A2(KEYINPUT23), .A3(G128), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n239), .A2(G119), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT23), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n363), .A2(new_n365), .B1(new_n317), .B2(G128), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n317), .A2(G128), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n364), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT24), .B(G110), .ZN(new_n369));
  OAI221_X1 g183(.A(new_n361), .B1(new_n362), .B2(new_n366), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n366), .A2(new_n362), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n360), .B1(G146), .B2(new_n357), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT22), .B(G137), .ZN(new_n375));
  INV_X1    g189(.A(G234), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n346), .A2(new_n376), .A3(G953), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n375), .B(new_n377), .Z(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n370), .A2(new_n373), .A3(new_n378), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G217), .B1(new_n376), .B2(G902), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n383), .B(KEYINPUT69), .Z(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G902), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n385), .B(KEYINPUT70), .Z(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT25), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n382), .B2(new_n284), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n380), .A2(new_n388), .A3(new_n284), .A4(new_n381), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n384), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n387), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT71), .ZN(new_n393));
  INV_X1    g207(.A(new_n193), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n189), .A2(G137), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n197), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n252), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n195), .A2(new_n197), .B1(new_n227), .B2(new_n230), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n314), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n245), .A2(new_n197), .A3(new_n396), .ZN(new_n401));
  INV_X1    g215(.A(new_n399), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n326), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(KEYINPUT28), .C1(new_n404), .C2(new_n403), .ZN(new_n406));
  NOR2_X1   g220(.A1(G237), .A2(G953), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G210), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(G101), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n398), .A2(new_n314), .A3(new_n399), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT28), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n406), .A2(KEYINPUT29), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n398), .B2(new_n399), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n401), .A2(KEYINPUT30), .A3(new_n402), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n314), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n403), .ZN(new_n419));
  INV_X1    g233(.A(new_n411), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(new_n400), .B2(new_n403), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n412), .A2(KEYINPUT28), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n426), .A2(new_n427), .A3(new_n420), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n414), .B(new_n284), .C1(new_n423), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G472), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n418), .A2(new_n411), .A3(new_n403), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT31), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT31), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n418), .A2(new_n434), .A3(new_n411), .A4(new_n403), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(G472), .A2(G902), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT32), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(KEYINPUT32), .A3(new_n437), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n430), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n436), .A2(KEYINPUT32), .A3(new_n437), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n438), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT68), .B1(new_n445), .B2(new_n430), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n393), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT72), .ZN(new_n448));
  INV_X1    g262(.A(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n451));
  INV_X1    g265(.A(G116), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n452), .B2(G122), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n449), .A2(KEYINPUT84), .A3(G116), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n202), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT84), .B1(new_n449), .B2(G116), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n452), .A3(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(G107), .A3(new_n450), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n450), .A2(KEYINPUT14), .A3(G107), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n459), .A2(KEYINPUT14), .A3(G107), .A4(new_n450), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n223), .A2(G128), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n239), .A2(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT85), .ZN(new_n467));
  XNOR2_X1  g281(.A(G128), .B(G143), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n470), .A3(G134), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n470), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n189), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n462), .A2(new_n463), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n189), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(new_n468), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n456), .A3(new_n460), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n348), .A2(G217), .A3(new_n272), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n485));
  INV_X1    g299(.A(G478), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(KEYINPUT15), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n480), .B1(new_n474), .B2(new_n478), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n284), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n487), .B1(new_n492), .B2(KEYINPUT86), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n485), .B(new_n284), .C1(new_n490), .C2(new_n491), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n407), .A2(G143), .A3(G214), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(G143), .B1(new_n407), .B2(G214), .ZN(new_n500));
  OAI21_X1  g314(.A(G131), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n407), .A2(G214), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n223), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n196), .A3(new_n498), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(KEYINPUT17), .B(G131), .C1(new_n499), .C2(new_n500), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n360), .A3(new_n359), .A4(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n200), .ZN(new_n510));
  XNOR2_X1  g324(.A(G125), .B(G140), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n221), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n504), .B(new_n498), .C1(new_n513), .C2(new_n196), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n514), .C1(new_n501), .C2(new_n513), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n508), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n510), .B1(new_n508), .B2(new_n515), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n497), .B(new_n284), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G475), .ZN(new_n520));
  INV_X1    g334(.A(new_n506), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n359), .A2(new_n507), .A3(new_n360), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n510), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n497), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n357), .A2(KEYINPUT19), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT19), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n511), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n530), .A3(new_n221), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n499), .A2(new_n500), .A3(G131), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n196), .B1(new_n504), .B2(new_n498), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n531), .B(new_n360), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n515), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n516), .B1(new_n535), .B2(new_n510), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n520), .A2(new_n527), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT87), .B(G952), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(G953), .ZN(new_n543));
  NAND2_X1  g357(.A1(G234), .A2(G237), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT21), .B(G898), .Z(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(G902), .A3(G953), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n496), .A2(new_n541), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n441), .A2(new_n442), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n445), .A2(KEYINPUT68), .A3(new_n430), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n393), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n350), .A2(new_n448), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT88), .B(G101), .Z(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(G3));
  INV_X1    g372(.A(new_n393), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n436), .A2(new_n437), .ZN(new_n560));
  INV_X1    g374(.A(G472), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n436), .B2(new_n284), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR4_X1   g377(.A1(new_n296), .A2(new_n559), .A3(new_n349), .A4(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n332), .A2(new_n299), .A3(new_n340), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n297), .B(new_n548), .C1(new_n565), .C2(new_n341), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n526), .A2(new_n497), .ZN(new_n567));
  INV_X1    g381(.A(G475), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n526), .B2(new_n497), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n536), .A2(new_n538), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT20), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n567), .A2(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT89), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n574), .A2(KEYINPUT89), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(new_n576), .C1(new_n490), .C2(new_n491), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n482), .A2(KEYINPUT89), .A3(new_n574), .A4(new_n483), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n486), .A2(G902), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n579), .A2(new_n580), .B1(new_n486), .B2(new_n492), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n566), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT90), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n564), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT91), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT34), .B(G104), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G6));
  INV_X1    g401(.A(new_n496), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n567), .A2(new_n569), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n571), .A2(new_n590), .A3(new_n572), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n548), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT93), .ZN(new_n596));
  INV_X1    g410(.A(new_n593), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n597), .A2(new_n598), .A3(new_n496), .A4(new_n548), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n596), .A2(KEYINPUT94), .A3(new_n344), .A4(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n344), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n598), .B1(new_n594), .B2(new_n548), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n564), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n202), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G9));
  NOR2_X1   g423(.A1(new_n389), .A2(new_n391), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n379), .A2(KEYINPUT36), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n374), .B(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n386), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n563), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n350), .A2(new_n550), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT37), .B(G110), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G12));
  NAND2_X1  g431(.A1(new_n291), .A2(new_n295), .ZN(new_n618));
  INV_X1    g432(.A(new_n285), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n349), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n547), .A2(G900), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n621), .A2(KEYINPUT96), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(KEYINPUT96), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n545), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n588), .A2(new_n593), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n613), .B1(new_n551), .B2(new_n552), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n620), .A2(new_n344), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT97), .B(G128), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G30));
  NAND2_X1  g444(.A1(new_n342), .A2(new_n343), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT38), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n405), .B1(new_n404), .B2(new_n403), .ZN(new_n633));
  OAI211_X1 g447(.A(G472), .B(new_n431), .C1(new_n633), .C2(new_n411), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n561), .A2(new_n284), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT98), .Z(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n445), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n588), .A2(new_n298), .A3(new_n573), .ZN(new_n640));
  AND4_X1   g454(.A1(new_n613), .A2(new_n632), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT99), .Z(new_n642));
  XOR2_X1   g456(.A(new_n624), .B(KEYINPUT39), .Z(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n620), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n645), .A2(KEYINPUT40), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(KEYINPUT40), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n642), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G143), .ZN(G45));
  NOR2_X1   g463(.A1(new_n573), .A2(new_n581), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n624), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n620), .A2(new_n344), .A3(new_n627), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT100), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n350), .A2(new_n655), .A3(new_n627), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G146), .ZN(G48));
  INV_X1    g472(.A(new_n447), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n660));
  INV_X1    g474(.A(new_n349), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n187), .B1(new_n293), .B2(new_n284), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n660), .A2(new_n618), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(new_n291), .B2(new_n295), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n660), .B1(new_n665), .B2(new_n661), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n659), .B(new_n583), .C1(new_n664), .C2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n618), .A2(new_n661), .A3(new_n663), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT101), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n665), .A2(new_n660), .A3(new_n661), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n673), .A2(KEYINPUT102), .A3(new_n659), .A4(new_n583), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  OAI211_X1 g491(.A(new_n659), .B(new_n605), .C1(new_n664), .C2(new_n666), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT103), .B(G116), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G18));
  NOR2_X1   g494(.A1(new_n670), .A2(new_n345), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n550), .A3(new_n627), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  AND2_X1   g497(.A1(new_n562), .A2(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n432), .A2(new_n435), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n411), .B1(new_n406), .B2(new_n413), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n437), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n687), .B1(new_n562), .B2(KEYINPUT104), .ZN(new_n688));
  OR3_X1    g502(.A1(new_n684), .A2(new_n688), .A3(new_n392), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n640), .A2(new_n631), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n549), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n664), .B2(new_n666), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G122), .ZN(G24));
  NOR3_X1   g507(.A1(new_n613), .A2(new_n684), .A3(new_n688), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n652), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n696), .A2(new_n344), .A3(new_n661), .A4(new_n665), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT105), .B(G125), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G27));
  INV_X1    g513(.A(new_n392), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n441), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT108), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n342), .A2(new_n297), .A3(new_n343), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n705), .B1(new_n620), .B2(new_n707), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n296), .A2(KEYINPUT106), .A3(new_n349), .A4(new_n706), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n704), .B(new_n652), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n659), .B(new_n652), .C1(new_n708), .C2(new_n709), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT42), .B1(new_n712), .B2(KEYINPUT107), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n618), .A2(new_n619), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n661), .A3(new_n707), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT106), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n620), .A2(new_n705), .A3(new_n707), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n659), .A4(new_n652), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n711), .B1(new_n713), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n196), .ZN(G33));
  NAND2_X1  g536(.A1(new_n659), .A2(new_n626), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n716), .B2(new_n717), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n189), .ZN(G36));
  INV_X1    g539(.A(new_n580), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n577), .B2(new_n578), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n484), .A2(G478), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n573), .ZN(new_n730));
  NAND2_X1  g544(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n733));
  MUX2_X1   g547(.A(new_n732), .B(new_n730), .S(new_n733), .Z(new_n734));
  INV_X1    g548(.A(new_n613), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n563), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n707), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT110), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n736), .A2(new_n741), .A3(new_n737), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n738), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n283), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n277), .A2(KEYINPUT45), .A3(new_n282), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(G469), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n618), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(KEYINPUT46), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n661), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n743), .A2(new_n644), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  NAND2_X1  g570(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n752), .A2(new_n758), .A3(new_n661), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n553), .A2(new_n393), .A3(new_n651), .A4(new_n706), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n763));
  NOR2_X1   g577(.A1(G952), .A2(G953), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n713), .A2(new_n720), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n710), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n678), .A2(new_n682), .A3(new_n692), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n496), .A2(KEYINPUT113), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n770), .B(new_n489), .C1(new_n493), .C2(new_n495), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n772), .A2(new_n593), .A3(new_n625), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n627), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n715), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n723), .A2(new_n695), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n775), .B1(new_n718), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n566), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT114), .B1(new_n772), .B2(new_n573), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n780), .B(new_n541), .C1(new_n769), .C2(new_n771), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n778), .C1(new_n779), .C2(new_n781), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT111), .B1(new_n573), .B2(new_n581), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n541), .B(new_n787), .C1(new_n728), .C2(new_n727), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n778), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n778), .B2(new_n789), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n783), .A2(new_n785), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n564), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n556), .A3(new_n615), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n675), .A2(new_n768), .A3(new_n777), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n767), .A2(new_n797), .A3(KEYINPUT116), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n675), .A2(new_n768), .A3(new_n777), .A4(new_n796), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n721), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n697), .A2(new_n628), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n690), .A2(new_n625), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n620), .A2(new_n613), .A3(new_n639), .A4(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n657), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n657), .A2(new_n807), .A3(new_n802), .A4(new_n804), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT53), .A4(new_n809), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n765), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n806), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n721), .A3(new_n800), .ZN(new_n816));
  AOI211_X1 g630(.A(KEYINPUT54), .B(new_n816), .C1(new_n810), .C2(new_n811), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n734), .A2(new_n544), .A3(new_n543), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n689), .ZN(new_n820));
  INV_X1    g634(.A(new_n632), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n298), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n822), .A2(new_n823), .A3(new_n670), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n823), .B1(new_n822), .B2(new_n670), .ZN(new_n825));
  INV_X1    g639(.A(new_n670), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n706), .A2(new_n545), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n559), .A3(new_n639), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n729), .A2(new_n541), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n824), .A2(new_n825), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n734), .A3(new_n827), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n694), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n757), .A2(new_n759), .B1(new_n349), .B2(new_n665), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n820), .A2(new_n707), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n831), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT51), .ZN(new_n838));
  INV_X1    g652(.A(new_n702), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT48), .B1(new_n840), .B2(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n829), .A2(new_n650), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n820), .A2(new_n681), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n543), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n841), .A2(new_n842), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n838), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n764), .B1(new_n818), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n665), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n852), .A2(KEYINPUT49), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(KEYINPUT49), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n700), .A2(new_n297), .A3(new_n661), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n632), .A2(new_n639), .A3(new_n855), .A4(new_n730), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n763), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n849), .A2(new_n814), .A3(new_n817), .ZN(new_n860));
  OAI211_X1 g674(.A(KEYINPUT119), .B(new_n857), .C1(new_n860), .C2(new_n764), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(G75));
  NAND2_X1  g676(.A1(new_n329), .A2(new_n331), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(new_n309), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n816), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n812), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(KEYINPUT120), .A3(G902), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n816), .B1(new_n810), .B2(new_n811), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n284), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n299), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n867), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n272), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n872), .A2(new_n284), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n880), .B2(new_n865), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n876), .A2(new_n881), .ZN(G51));
  NOR2_X1   g696(.A1(new_n872), .A2(new_n765), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n817), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n748), .B(KEYINPUT57), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n293), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n747), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n874), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n877), .B1(new_n886), .B2(new_n888), .ZN(G54));
  NAND2_X1  g703(.A1(KEYINPUT58), .A2(G475), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT122), .Z(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n870), .B2(new_n873), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n536), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n878), .B1(new_n892), .B2(new_n536), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(G60));
  NAND2_X1  g709(.A1(G478), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT59), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n818), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n579), .ZN(new_n899));
  INV_X1    g713(.A(new_n897), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n579), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n878), .B1(new_n884), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(G63));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT60), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n869), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n382), .B(KEYINPUT123), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n869), .A2(new_n612), .A3(new_n905), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n878), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n908), .A2(KEYINPUT61), .A3(new_n878), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(G66));
  INV_X1    g728(.A(new_n546), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n915), .B2(new_n302), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n675), .A2(new_n768), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n796), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n919), .B2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n863), .B1(G898), .B2(new_n272), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G69));
  AND2_X1   g736(.A1(new_n755), .A2(new_n761), .ZN(new_n923));
  INV_X1    g737(.A(new_n645), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n779), .A2(new_n781), .A3(new_n789), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n706), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n448), .A3(new_n555), .A4(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n657), .A2(new_n802), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n648), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n648), .A3(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n928), .A2(new_n934), .A3(KEYINPUT124), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT124), .B1(new_n928), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n272), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n416), .A2(new_n417), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n528), .A2(new_n530), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n724), .ZN(new_n943));
  OR4_X1    g757(.A1(new_n643), .A2(new_n753), .A3(new_n690), .A4(new_n702), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n923), .A2(new_n943), .A3(new_n929), .A4(new_n944), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n945), .A2(G953), .A3(new_n721), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(G900), .B2(G953), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n949));
  AOI22_X1  g763(.A1(new_n946), .A2(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n948), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n951), .B(new_n952), .Z(G72));
  NOR2_X1   g767(.A1(new_n419), .A2(new_n411), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n945), .A2(new_n721), .A3(new_n918), .ZN(new_n955));
  XNOR2_X1  g769(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n635), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n878), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n928), .A2(new_n934), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n928), .A2(new_n934), .A3(KEYINPUT124), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n919), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n957), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n419), .A2(new_n411), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n959), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n812), .A2(new_n813), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n421), .A2(new_n431), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n965), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n969), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(G57));
endmodule


