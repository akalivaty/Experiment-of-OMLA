//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT5), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n206), .A2(new_n208), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n211), .A2(G148gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n209), .A2(G141gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n205), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n207), .A2(new_n204), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT74), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT2), .B1(new_n210), .B2(new_n212), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n223));
  XNOR2_X1  g022(.A(G155gat), .B(G162gat), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n214), .B(new_n216), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G134gat), .ZN(new_n227));
  INV_X1    g026(.A(G127gat), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G113gat), .ZN(new_n230));
  INV_X1    g029(.A(G113gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n228), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI211_X1 g034(.A(KEYINPUT1), .B(G127gat), .C1(new_n230), .C2(new_n232), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n227), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238));
  OAI21_X1  g037(.A(G127gat), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n233), .A2(new_n234), .A3(new_n228), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(G134gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n223), .B1(new_n222), .B2(new_n224), .ZN(new_n244));
  XNOR2_X1  g043(.A(G141gat), .B(G148gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n220), .B(KEYINPUT74), .C1(new_n245), .C2(KEYINPUT2), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n213), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n226), .B(new_n242), .C1(new_n243), .C2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT76), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n246), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(new_n251), .B2(new_n214), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n253), .A2(KEYINPUT76), .A3(new_n242), .A4(new_n226), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n214), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n242), .B2(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n239), .A2(new_n240), .A3(G134gat), .ZN(new_n260));
  AOI21_X1  g059(.A(G134gat), .B1(new_n239), .B2(new_n240), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(KEYINPUT4), .A3(new_n247), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  AND4_X1   g063(.A1(new_n203), .A2(new_n255), .A3(new_n256), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n256), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n242), .A2(new_n258), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n247), .B1(new_n241), .B2(new_n237), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n263), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n250), .B2(new_n254), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n272), .B2(new_n256), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G57gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G85gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  NOR3_X1   g078(.A1(new_n274), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(KEYINPUT79), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI211_X1 g081(.A(new_n213), .B(new_n215), .C1(new_n244), .C2(new_n246), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n252), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT76), .B1(new_n284), .B2(new_n242), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n248), .A2(new_n249), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n256), .B(new_n264), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n270), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n203), .A3(new_n256), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n289), .A2(KEYINPUT81), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT81), .B1(new_n289), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n282), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT82), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT81), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n265), .B2(new_n273), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n289), .A2(KEYINPUT81), .A3(new_n290), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n282), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT6), .B1(new_n274), .B2(new_n279), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n280), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G15gat), .B(G43gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G227gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  OR3_X1    g110(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G183gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(G190gat), .B1(new_n318), .B2(KEYINPUT67), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT28), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n321), .A2(new_n326), .A3(G190gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n311), .B(new_n316), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  OR3_X1    g127(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n329), .A2(new_n330), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n317), .A2(new_n334), .A3(KEYINPUT66), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT66), .B1(new_n317), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(KEYINPUT25), .B(new_n331), .C1(new_n337), .C2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n342));
  INV_X1    g141(.A(new_n330), .ZN(new_n343));
  NOR3_X1   g142(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n344));
  OAI22_X1  g143(.A1(new_n343), .A2(new_n344), .B1(new_n314), .B2(new_n315), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n317), .A2(new_n334), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n333), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n342), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n262), .A2(new_n328), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n262), .B1(new_n328), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n310), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT68), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n349), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n242), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n350), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n310), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n307), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n357), .B2(new_n310), .ZN(new_n363));
  INV_X1    g162(.A(new_n310), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT68), .B(new_n364), .C1(new_n356), .C2(new_n350), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT32), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n356), .A2(new_n364), .A3(new_n350), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT34), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT34), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n356), .A2(new_n369), .A3(new_n364), .A4(new_n350), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n360), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n362), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n361), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n373), .A2(new_n374), .B1(new_n376), .B2(new_n306), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G228gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(new_n309), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n226), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n383), .A2(KEYINPUT70), .ZN(new_n384));
  XNOR2_X1  g183(.A(G197gat), .B(G204gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(KEYINPUT70), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT71), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G211gat), .B(G218gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n392), .A2(KEYINPUT72), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT72), .B1(new_n392), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n382), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT70), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n383), .B(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT71), .B1(new_n398), .B2(new_n385), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n393), .B(new_n381), .C1(new_n399), .C2(new_n390), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n392), .A2(KEYINPUT77), .A3(new_n381), .A4(new_n393), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n402), .A2(new_n243), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n380), .B(new_n396), .C1(new_n404), .C2(new_n247), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n392), .A2(new_n393), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n382), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n390), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n398), .A2(new_n391), .A3(new_n385), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n381), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n247), .B1(new_n410), .B2(new_n216), .ZN(new_n411));
  OAI22_X1  g210(.A1(new_n407), .A2(new_n411), .B1(new_n379), .B2(new_n309), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G22gat), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n405), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n415), .B1(new_n405), .B2(new_n412), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT78), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n414), .A2(new_n422), .A3(new_n416), .A4(new_n420), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT35), .ZN(new_n427));
  XNOR2_X1  g226(.A(G8gat), .B(G36gat), .ZN(new_n428));
  INV_X1    g227(.A(G64gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G92gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n394), .A2(new_n395), .ZN(new_n433));
  AND2_X1   g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n328), .B2(new_n349), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT73), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n355), .A2(new_n381), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n435), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(new_n438), .B2(new_n435), .ZN(new_n441));
  INV_X1    g240(.A(new_n406), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n432), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n355), .A2(new_n434), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT73), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n436), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n439), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n433), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n450), .A2(new_n451), .B1(new_n441), .B2(new_n442), .ZN(new_n452));
  INV_X1    g251(.A(new_n432), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n445), .A2(new_n454), .A3(KEYINPUT30), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n378), .A2(new_n426), .A3(new_n427), .A4(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n202), .B1(new_n303), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n299), .B1(new_n298), .B2(new_n282), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT82), .B(new_n281), .C1(new_n296), .C2(new_n297), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n302), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n280), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND4_X1   g264(.A1(new_n427), .A2(new_n378), .A3(new_n426), .A4(new_n458), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT84), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n302), .B1(new_n279), .B2(new_n274), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n464), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n458), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n378), .A2(new_n426), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n460), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n426), .ZN(new_n474));
  OR3_X1    g273(.A1(new_n267), .A2(new_n268), .A3(new_n266), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT39), .B(new_n475), .C1(new_n272), .C2(new_n256), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n255), .A2(new_n264), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n266), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n479), .A3(new_n281), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT80), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n455), .A3(new_n457), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n294), .B2(new_n300), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT40), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n474), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI22_X1  g286(.A1(new_n450), .A2(new_n451), .B1(new_n441), .B2(new_n442), .ZN(new_n488));
  AOI211_X1 g287(.A(KEYINPUT38), .B(new_n453), .C1(new_n488), .C2(KEYINPUT37), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n452), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n454), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n450), .A2(new_n451), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n494), .B2(new_n443), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT83), .B1(new_n495), .B2(new_n453), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n432), .C1(new_n452), .C2(new_n490), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n493), .B1(new_n499), .B2(KEYINPUT38), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n463), .A2(new_n464), .A3(new_n492), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n487), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT36), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n503), .A2(KEYINPUT36), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n378), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n503), .B(KEYINPUT36), .C1(new_n375), .C2(new_n377), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n426), .B1(new_n469), .B2(new_n458), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n473), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G230gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n309), .ZN(new_n514));
  NAND2_X1  g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  INV_X1    g314(.A(G71gat), .ZN(new_n516));
  INV_X1    g315(.A(G78gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n519));
  AND2_X1   g318(.A1(G57gat), .A2(G64gat), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n515), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(KEYINPUT9), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(KEYINPUT95), .A2(G57gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n429), .ZN(new_n526));
  NAND3_X1  g325(.A1(KEYINPUT95), .A2(G57gat), .A3(G64gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n521), .B(KEYINPUT101), .C1(new_n524), .C2(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT97), .B(G85gat), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n533), .A2(new_n431), .B1(KEYINPUT8), .B2(new_n531), .ZN(new_n534));
  AND3_X1   g333(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n532), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n431), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n531), .A2(KEYINPUT8), .ZN(new_n542));
  AND4_X1   g341(.A1(new_n532), .A2(new_n537), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n529), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT10), .ZN(new_n545));
  INV_X1    g344(.A(new_n529), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n518), .A2(new_n515), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n515), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n547), .A2(new_n549), .A3(new_n526), .A4(new_n527), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT101), .B1(new_n550), .B2(new_n521), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n531), .A3(new_n530), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n532), .A3(new_n537), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n544), .B(new_n545), .C1(new_n552), .C2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n550), .A2(new_n521), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n514), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n544), .B1(new_n552), .B2(new_n556), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n514), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n315), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G204gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n563), .A2(new_n565), .A3(new_n569), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G113gat), .B(G141gat), .Z(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G169gat), .B(G197gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT12), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT16), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(G1gat), .ZN(new_n582));
  INV_X1    g381(.A(G15gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G22gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n415), .A2(G15gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n586), .B(new_n587), .C1(G1gat), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT89), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n586), .B(new_n591), .C1(G1gat), .C2(new_n588), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(G8gat), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G8gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(KEYINPUT89), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT17), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(KEYINPUT17), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G50gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G43gat), .ZN(new_n602));
  INV_X1    g401(.A(G43gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(G50gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n604), .A3(KEYINPUT15), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(KEYINPUT88), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT88), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G43gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n608), .A3(new_n601), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT15), .B1(new_n609), .B2(new_n604), .ZN(new_n610));
  OR2_X1    g409(.A1(KEYINPUT87), .A2(G29gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(KEYINPUT87), .A2(G29gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(G36gat), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT14), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(G29gat), .B2(G36gat), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n614), .A2(G29gat), .A3(G36gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n605), .B1(new_n610), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n605), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n619), .A2(new_n615), .A3(new_n613), .A4(new_n616), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n598), .B(new_n600), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  AND4_X1   g420(.A1(new_n597), .A2(new_n618), .A3(KEYINPUT17), .A4(new_n620), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n596), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT92), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n618), .A2(new_n620), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n627));
  AOI21_X1  g426(.A(G1gat), .B1(new_n584), .B2(new_n585), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n628), .B1(new_n588), .B2(new_n582), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n591), .B1(new_n629), .B2(new_n587), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n592), .A2(G8gat), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n627), .B(new_n595), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n627), .B1(new_n593), .B2(new_n595), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n626), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n598), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n625), .A2(new_n637), .A3(new_n599), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n618), .A2(new_n620), .A3(new_n597), .A4(KEYINPUT17), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT92), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n596), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n624), .A2(new_n635), .A3(new_n636), .A4(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT18), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n643), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n636), .B(KEYINPUT13), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n634), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n625), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n650), .B2(new_n635), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT86), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n580), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n647), .ZN(new_n655));
  INV_X1    g454(.A(new_n651), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(KEYINPUT86), .A3(new_n579), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n512), .A2(new_n573), .A3(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n596), .A2(KEYINPUT93), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n632), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(G183gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n649), .A2(new_n317), .A3(new_n668), .ZN(new_n671));
  XOR2_X1   g470(.A(G127gat), .B(G155gat), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n670), .B2(new_n671), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT96), .B(G211gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(G231gat), .A2(G233gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n675), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n670), .A2(new_n671), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n672), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n683), .B2(new_n674), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n666), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n679), .B1(new_n675), .B2(new_n676), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n681), .A3(new_n674), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n665), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n640), .A2(new_n556), .ZN(new_n689));
  XNOR2_X1  g488(.A(G190gat), .B(G218gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT98), .ZN(new_n691));
  AND2_X1   g490(.A1(G232gat), .A2(G233gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT41), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n626), .A2(new_n558), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n689), .A2(new_n691), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n698));
  INV_X1    g497(.A(new_n691), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n695), .A2(new_n696), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n695), .A2(new_n696), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT100), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n692), .A2(KEYINPUT41), .ZN(new_n705));
  XNOR2_X1  g504(.A(G134gat), .B(G162gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n697), .B(new_n700), .C1(KEYINPUT100), .C2(new_n709), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n685), .A2(new_n688), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n662), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n469), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G1gat), .ZN(G1324gat));
  INV_X1    g515(.A(new_n458), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n581), .A2(new_n594), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n662), .A2(new_n711), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n581), .A2(new_n594), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G8gat), .B1(new_n712), .B2(new_n458), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT102), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n722), .A2(new_n727), .A3(new_n723), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(G1325gat));
  NOR3_X1   g528(.A1(new_n712), .A2(new_n583), .A3(new_n509), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n378), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n583), .B2(new_n731), .ZN(G1326gat));
  NOR2_X1   g531(.A1(new_n712), .A2(new_n426), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT43), .B(G22gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT103), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n733), .B(new_n735), .ZN(G1327gat));
  NAND2_X1  g535(.A1(new_n708), .A2(new_n710), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n460), .A2(new_n472), .A3(new_n467), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n511), .B(new_n508), .C1(new_n487), .C2(new_n501), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n685), .A2(new_n688), .ZN(new_n743));
  INV_X1    g542(.A(new_n573), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n660), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n469), .B1(new_n611), .B2(new_n612), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT45), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n741), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n512), .A2(KEYINPUT44), .A3(new_n738), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(new_n745), .A3(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n611), .B(new_n612), .C1(new_n754), .C2(new_n469), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n755), .ZN(G1328gat));
  NOR3_X1   g555(.A1(new_n746), .A2(G36gat), .A3(new_n458), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g557(.A(G36gat), .B1(new_n754), .B2(new_n458), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1329gat));
  AND2_X1   g559(.A1(new_n606), .A2(new_n608), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n754), .B2(new_n509), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT47), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n378), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(new_n761), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n746), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n764), .B(new_n767), .ZN(G1330gat));
  NOR2_X1   g567(.A1(new_n426), .A2(G50gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT105), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n474), .A3(new_n745), .A4(new_n753), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n747), .A2(new_n770), .B1(new_n771), .B2(G50gat), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g572(.A1(new_n512), .A2(new_n711), .A3(new_n660), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n744), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n714), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n744), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n458), .B(new_n778), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1333gat));
  NAND4_X1  g580(.A1(new_n775), .A2(KEYINPUT106), .A3(G71gat), .A4(new_n508), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n774), .A2(G71gat), .A3(new_n744), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n509), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n516), .B1(new_n778), .B2(new_n765), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT50), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n790), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1334gat));
  NOR2_X1   g591(.A1(new_n778), .A2(new_n426), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(new_n517), .ZN(G1335gat));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  INV_X1    g594(.A(new_n743), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n660), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n741), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n661), .A2(new_n743), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n512), .A2(KEYINPUT51), .A3(new_n738), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n801), .A2(new_n799), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT108), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT108), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n533), .B(new_n744), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n752), .A2(new_n744), .A3(new_n753), .A4(new_n800), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n469), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n806), .A2(new_n469), .B1(new_n533), .B2(new_n808), .ZN(G1336gat));
  OAI21_X1  g608(.A(G92gat), .B1(new_n807), .B2(new_n458), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT109), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n798), .A2(new_n801), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n458), .A2(G92gat), .A3(new_n573), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n815), .B(G92gat), .C1(new_n807), .C2(new_n458), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT52), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n813), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n810), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(G1337gat));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n823));
  OR3_X1    g622(.A1(new_n807), .A2(new_n823), .A3(new_n509), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n807), .B2(new_n509), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(G99gat), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(G99gat), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(new_n744), .C1(new_n804), .C2(new_n805), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n828), .B2(new_n765), .ZN(G1338gat));
  OR2_X1    g628(.A1(new_n807), .A2(new_n426), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n426), .A2(G106gat), .A3(new_n573), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n802), .A2(new_n803), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n830), .A2(G106gat), .B1(new_n812), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n832), .ZN(G1339gat));
  NOR2_X1   g636(.A1(new_n469), .A2(new_n717), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n557), .A2(new_n561), .A3(new_n514), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n563), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI211_X1 g641(.A(KEYINPUT112), .B(new_n569), .C1(new_n562), .C2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n557), .A2(new_n561), .ZN(new_n845));
  INV_X1    g644(.A(new_n514), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n570), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n841), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(KEYINPUT55), .B(new_n841), .C1(new_n843), .C2(new_n848), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n572), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n851), .A2(KEYINPUT113), .A3(new_n572), .A4(new_n852), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n855), .A2(new_n654), .A3(new_n659), .A4(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n624), .A2(new_n642), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n636), .B1(new_n858), .B2(new_n635), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n650), .A2(new_n635), .A3(new_n648), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n652), .A2(new_n579), .B1(new_n861), .B2(new_n578), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n744), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n738), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n738), .A2(new_n855), .A3(new_n856), .A4(new_n862), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n796), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n711), .A2(new_n660), .A3(new_n573), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT111), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n711), .A2(new_n660), .A3(new_n869), .A4(new_n573), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n866), .A2(new_n871), .A3(KEYINPUT114), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n426), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n874), .A2(KEYINPUT115), .A3(new_n426), .A4(new_n875), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n765), .B(new_n839), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n231), .B1(new_n880), .B2(new_n661), .ZN(new_n881));
  INV_X1    g680(.A(new_n471), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n874), .A2(new_n882), .A3(new_n875), .A4(new_n838), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(G113gat), .A3(new_n660), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n881), .A2(new_n884), .ZN(G1340gat));
  AOI21_X1  g684(.A(new_n229), .B1(new_n880), .B2(new_n744), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n883), .A2(G120gat), .A3(new_n573), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(G1341gat));
  AOI21_X1  g687(.A(new_n839), .B1(new_n878), .B2(new_n879), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n889), .A2(G127gat), .A3(new_n743), .A4(new_n378), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n880), .A2(KEYINPUT116), .A3(G127gat), .A4(new_n743), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n228), .B1(new_n883), .B2(new_n796), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G1342gat));
  NOR2_X1   g694(.A1(new_n737), .A2(G134gat), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT56), .B1(new_n883), .B2(new_n897), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n897), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n880), .A2(new_n738), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n227), .ZN(G1343gat));
  OAI21_X1  g700(.A(new_n863), .B1(new_n660), .B2(new_n853), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n865), .B1(new_n737), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n871), .B1(new_n903), .B2(new_n743), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(KEYINPUT57), .A3(new_n474), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n874), .A2(new_n875), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n426), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n839), .A2(new_n508), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n909), .A2(G141gat), .A3(new_n661), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n907), .A2(new_n910), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n211), .B1(new_n912), .B2(new_n660), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n911), .A2(KEYINPUT58), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1344gat));
  INV_X1    g717(.A(new_n912), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n209), .A3(new_n744), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n909), .A2(new_n744), .A3(new_n910), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(G148gat), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n874), .A2(new_n474), .A3(new_n875), .A4(new_n908), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  INV_X1    g724(.A(new_n867), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n902), .A2(new_n737), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n862), .A2(new_n738), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n853), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n926), .B1(new_n929), .B2(new_n796), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n930), .B2(new_n426), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n744), .A3(new_n910), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n209), .B1(new_n933), .B2(KEYINPUT118), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n932), .A2(new_n935), .A3(new_n744), .A4(new_n910), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n922), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n920), .B1(new_n923), .B2(new_n937), .ZN(G1345gat));
  AOI21_X1  g737(.A(G155gat), .B1(new_n919), .B2(new_n743), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n909), .A2(new_n910), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n743), .A2(G155gat), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT119), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n939), .B1(new_n941), .B2(new_n943), .ZN(G1346gat));
  OAI21_X1  g743(.A(KEYINPUT121), .B1(new_n940), .B2(new_n737), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n909), .A2(new_n946), .A3(new_n738), .A4(new_n910), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(G162gat), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n737), .A2(G162gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n919), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n919), .A2(KEYINPUT120), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n948), .A2(new_n954), .ZN(G1347gat));
  NAND2_X1  g754(.A1(new_n882), .A2(new_n717), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT122), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n874), .A2(new_n469), .A3(new_n875), .A4(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n314), .A3(new_n661), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n714), .A2(new_n458), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n878), .B2(new_n879), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n661), .A3(new_n378), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT123), .B1(new_n964), .B2(G169gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(G1348gat));
  NAND4_X1  g766(.A1(new_n963), .A2(G176gat), .A3(new_n744), .A4(new_n378), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n315), .B1(new_n958), .B2(new_n573), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(G1349gat));
  XNOR2_X1  g769(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n878), .A2(new_n879), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n972), .A2(new_n743), .A3(new_n378), .A4(new_n961), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G183gat), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n796), .A3(new_n321), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n971), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n971), .ZN(new_n978));
  AOI211_X1 g777(.A(new_n978), .B(new_n975), .C1(new_n973), .C2(G183gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n977), .A2(new_n979), .ZN(G1350gat));
  NAND3_X1  g779(.A1(new_n959), .A2(new_n334), .A3(new_n738), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n738), .A3(new_n378), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n982), .A2(new_n983), .A3(G190gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n982), .B2(G190gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  NOR2_X1   g785(.A1(new_n962), .A2(new_n508), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n932), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n661), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(G197gat), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n906), .A2(new_n714), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n508), .A2(new_n426), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n991), .A2(new_n717), .A3(new_n992), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n993), .A2(G197gat), .A3(new_n660), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(G1352gat));
  INV_X1    g797(.A(G204gat), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n991), .A2(new_n999), .A3(new_n717), .A4(new_n992), .ZN(new_n1000));
  OAI21_X1  g799(.A(KEYINPUT62), .B1(new_n1000), .B2(new_n573), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n932), .A2(new_n744), .A3(new_n987), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(G204gat), .ZN(new_n1003));
  INV_X1    g802(.A(new_n992), .ZN(new_n1004));
  NOR4_X1   g803(.A1(new_n906), .A2(new_n714), .A3(new_n458), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n1005), .A2(new_n1006), .A3(new_n999), .A4(new_n744), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1001), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n1001), .A2(new_n1003), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1353gat));
  OR3_X1    g811(.A1(new_n993), .A2(G211gat), .A3(new_n796), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n988), .A2(new_n743), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1014), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1015));
  AOI21_X1  g814(.A(KEYINPUT63), .B1(new_n1014), .B2(G211gat), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(G1354gat));
  AOI21_X1  g816(.A(G218gat), .B1(new_n1005), .B2(new_n738), .ZN(new_n1018));
  AND2_X1   g817(.A1(new_n1018), .A2(KEYINPUT127), .ZN(new_n1019));
  AND3_X1   g818(.A1(new_n988), .A2(G218gat), .A3(new_n738), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1018), .A2(KEYINPUT127), .ZN(new_n1021));
  NOR3_X1   g820(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(G1355gat));
endmodule


