//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n203), .A2(new_n216), .B1(new_n208), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  AOI211_X1 g0020(.A(new_n218), .B(new_n220), .C1(G77), .C2(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n206), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n215), .B(new_n228), .C1(new_n235), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT67), .B(G250), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  INV_X1    g0052(.A(G50), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n202), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n257), .A2(new_n229), .A3(G1), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  XOR2_X1   g0059(.A(KEYINPUT8), .B(G58), .Z(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n234), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G20), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n265), .B2(new_n260), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n233), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n229), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT7), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(new_n275), .A3(G68), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G58), .A2(G68), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n204), .A2(new_n205), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT74), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G159), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n278), .A2(new_n286), .A3(G20), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n276), .A2(new_n280), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT16), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n263), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n278), .A2(new_n286), .A3(G20), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n286), .B1(new_n278), .B2(G20), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n291), .A2(new_n292), .A3(new_n284), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n233), .A2(new_n269), .A3(KEYINPUT7), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n274), .A2(new_n270), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n203), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT16), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n266), .B1(new_n290), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G223), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G226), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n308), .C1(new_n267), .C2(new_n268), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G41), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(G1), .A3(G13), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n303), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n313), .A2(G232), .A3(new_n301), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n300), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n313), .B1(new_n309), .B2(new_n310), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NOR4_X1   g0120(.A1(new_n319), .A2(new_n320), .A3(new_n316), .A4(new_n303), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT75), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n315), .A2(G179), .A3(new_n317), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n319), .A2(new_n303), .A3(new_n316), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n300), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n299), .A2(new_n327), .A3(KEYINPUT18), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT18), .B1(new_n299), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT76), .B(G190), .Z(new_n331));
  NAND3_X1  g0131(.A1(new_n315), .A2(new_n331), .A3(new_n317), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n325), .B2(G200), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n266), .B(new_n333), .C1(new_n290), .C2(new_n298), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n280), .A2(new_n285), .A3(new_n287), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n289), .B1(new_n337), .B2(new_n296), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n291), .A2(new_n292), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n339), .A2(KEYINPUT16), .A3(new_n285), .A4(new_n276), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n263), .A3(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n341), .A2(KEYINPUT17), .A3(new_n266), .A4(new_n333), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n330), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g0144(.A(new_n344), .B(KEYINPUT77), .Z(new_n345));
  INV_X1    g0145(.A(new_n263), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n347));
  INV_X1    g0147(.A(G33), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n230), .B2(new_n232), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n260), .B1(G150), .B2(new_n281), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n346), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n265), .A2(G50), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n259), .A2(G50), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n272), .A2(new_n273), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n305), .A2(G222), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(new_n357), .C1(new_n304), .C2(new_n305), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n314), .C1(G77), .C2(new_n356), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n313), .A2(new_n301), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G226), .ZN(new_n361));
  INV_X1    g0161(.A(new_n303), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(G200), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n355), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n367), .A2(KEYINPUT10), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT10), .B1(new_n367), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n363), .A2(new_n300), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G179), .B2(new_n363), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n354), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G238), .A2(G1698), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n356), .B(new_n377), .C1(new_n222), .C2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n314), .C1(G107), .C2(new_n356), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n360), .A2(G244), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n362), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(G179), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n300), .B2(new_n381), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(KEYINPUT69), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(KEYINPUT69), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(new_n349), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT65), .B(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n260), .A2(new_n281), .B1(new_n388), .B2(G77), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(new_n263), .B1(G77), .B2(new_n265), .ZN(new_n391));
  INV_X1    g0191(.A(G77), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n258), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT70), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n383), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n372), .A2(new_n376), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n360), .A2(G238), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n356), .A2(G232), .A3(G1698), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n348), .B2(new_n208), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n356), .A2(new_n401), .A3(G226), .A4(new_n305), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n356), .A2(G226), .A3(new_n305), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT71), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n362), .B(new_n398), .C1(new_n405), .C2(new_n313), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT13), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n404), .A2(new_n402), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n314), .B1(new_n408), .B2(new_n400), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n362), .A4(new_n398), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G169), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT14), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(G179), .A3(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n416), .A3(G169), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n349), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT72), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n281), .A2(G50), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n420), .B1(new_n425), .B2(new_n346), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n263), .A3(new_n419), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n265), .A2(G68), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n257), .A2(G1), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(G20), .A3(new_n203), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT12), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n418), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n412), .A2(new_n364), .ZN(new_n434));
  INV_X1    g0234(.A(G200), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n407), .B2(new_n411), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n381), .A2(new_n364), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n381), .A2(G200), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n391), .A3(new_n394), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n433), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n345), .A2(new_n397), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT84), .ZN(new_n444));
  NAND2_X1  g0244(.A1(KEYINPUT6), .A2(G97), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT78), .B1(new_n445), .B2(G107), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(new_n209), .A3(KEYINPUT6), .A4(G97), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G97), .A2(G107), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT6), .B1(new_n210), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n452), .A2(new_n233), .B1(new_n392), .B2(new_n282), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n209), .B1(new_n294), .B2(new_n295), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n263), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n258), .B1(new_n264), .B2(G33), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n346), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n258), .A2(new_n208), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n455), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1698), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(G244), .C1(new_n268), .C2(new_n267), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  INV_X1    g0266(.A(G244), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n272), .B2(new_n273), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n465), .B(new_n466), .C1(new_n468), .C2(KEYINPUT4), .ZN(new_n469));
  OAI21_X1  g0269(.A(G250), .B1(new_n267), .B2(new_n268), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n305), .B1(new_n470), .B2(KEYINPUT4), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n314), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G41), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n264), .B(G45), .C1(new_n473), .C2(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G41), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(new_n313), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n234), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(new_n312), .B1(KEYINPUT5), .B2(new_n473), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(G41), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT79), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n264), .A4(G45), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n479), .A2(new_n480), .A3(G274), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n472), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n462), .B1(new_n485), .B2(new_n364), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(G200), .ZN(new_n487));
  INV_X1    g0287(.A(new_n484), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n224), .B1(new_n272), .B2(new_n273), .ZN(new_n489));
  OAI21_X1  g0289(.A(G1698), .B1(new_n489), .B2(new_n463), .ZN(new_n490));
  OAI21_X1  g0290(.A(G244), .B1(new_n267), .B2(new_n268), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(new_n463), .B1(G33), .B2(G283), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n492), .A3(new_n465), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n493), .B2(new_n314), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(KEYINPUT80), .A3(G190), .A4(new_n477), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n461), .A2(new_n486), .A3(new_n487), .A4(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n472), .A2(new_n320), .A3(new_n477), .A4(new_n484), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT81), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n455), .A2(new_n459), .A3(new_n460), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT81), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n494), .A2(new_n500), .A3(new_n320), .A4(new_n477), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n485), .A2(new_n300), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n498), .A2(new_n499), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n388), .A2(new_n505), .B1(G87), .B2(new_n210), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n356), .A2(new_n233), .A3(G68), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT19), .B1(new_n349), .B2(G97), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n263), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n385), .A2(new_n386), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n258), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n456), .A2(new_n385), .A3(new_n346), .A4(new_n386), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n216), .A2(new_n305), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n467), .A2(G1698), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n517), .C1(new_n267), .C2(new_n268), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n314), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n264), .A2(G45), .ZN(new_n522));
  AND2_X1   g0322(.A1(G33), .A2(G41), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(G250), .C1(new_n523), .C2(new_n234), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT82), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n313), .A2(KEYINPUT82), .A3(G250), .A4(new_n522), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n264), .A2(G45), .A3(G274), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n521), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n521), .A2(new_n528), .A3(G179), .A4(new_n529), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n510), .A2(new_n534), .A3(new_n512), .A4(new_n513), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n515), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n510), .A2(new_n512), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(G200), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n521), .A2(new_n528), .A3(G190), .A4(new_n529), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n458), .A2(G87), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n444), .B1(new_n504), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n229), .A2(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n429), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n457), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n545), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n348), .A2(G97), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n233), .A2(new_n466), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT86), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n230), .A2(new_n232), .B1(G33), .B2(G283), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT86), .B1(new_n554), .B2(new_n550), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n263), .B(new_n549), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(new_n552), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n554), .A2(KEYINPUT86), .A3(new_n550), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n346), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(KEYINPUT20), .A3(new_n549), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n548), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n305), .A2(G257), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G264), .A2(G1698), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n267), .C2(new_n268), .ZN(new_n566));
  XNOR2_X1  g0366(.A(KEYINPUT85), .B(G303), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n314), .C1(new_n356), .C2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G270), .B(new_n313), .C1(new_n474), .C2(new_n476), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n484), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G169), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n544), .B1(new_n563), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT87), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n571), .A2(new_n544), .B1(new_n320), .B2(new_n570), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n573), .B1(new_n575), .B2(new_n563), .ZN(new_n576));
  INV_X1    g0376(.A(new_n548), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n556), .A2(new_n557), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n561), .B2(new_n549), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n574), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n570), .A2(new_n331), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(G200), .B2(new_n570), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n563), .A2(new_n583), .ZN(new_n584));
  AND4_X1   g0384(.A1(new_n572), .A2(new_n576), .A3(new_n581), .A4(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n536), .A2(new_n541), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(KEYINPUT84), .A3(new_n503), .A4(new_n496), .ZN(new_n587));
  OAI211_X1 g0387(.A(G264), .B(new_n313), .C1(new_n474), .C2(new_n476), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n224), .A2(new_n305), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n217), .A2(G1698), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n267), .C2(new_n268), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(KEYINPUT89), .B(new_n588), .C1(new_n593), .C2(new_n313), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT89), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n313), .B1(new_n591), .B2(new_n592), .ZN(new_n596));
  INV_X1    g0396(.A(new_n588), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G179), .A3(new_n484), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n484), .B(new_n588), .C1(new_n593), .C2(new_n313), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT88), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n596), .A2(new_n597), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(new_n484), .ZN(new_n605));
  OAI21_X1  g0405(.A(G169), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(KEYINPUT23), .A2(G107), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(G20), .ZN(new_n610));
  NOR2_X1   g0410(.A1(KEYINPUT23), .A2(G107), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n388), .B2(new_n611), .ZN(new_n612));
  NOR4_X1   g0412(.A1(new_n269), .A2(new_n388), .A3(KEYINPUT22), .A4(new_n223), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT22), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n230), .A2(new_n232), .B1(new_n272), .B2(new_n273), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(G87), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n612), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT24), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n612), .B(KEYINPUT24), .C1(new_n613), .C2(new_n616), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n263), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n458), .A2(G107), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n258), .A2(new_n209), .ZN(new_n623));
  XOR2_X1   g0423(.A(new_n623), .B(KEYINPUT25), .Z(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n607), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n594), .A2(new_n598), .A3(new_n484), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n435), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n604), .A2(new_n603), .A3(new_n484), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n364), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(new_n622), .A3(new_n624), .A4(new_n621), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n543), .A2(new_n585), .A3(new_n587), .A4(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n443), .A2(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n372), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n336), .A2(new_n342), .ZN(new_n638));
  INV_X1    g0438(.A(new_n432), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n416), .B1(new_n412), .B2(G169), .ZN(new_n640));
  AOI211_X1 g0440(.A(KEYINPUT14), .B(new_n300), .C1(new_n407), .C2(new_n411), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n415), .ZN(new_n643));
  INV_X1    g0443(.A(new_n396), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n438), .B(new_n638), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n318), .A2(new_n321), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n299), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n299), .A2(KEYINPUT18), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n637), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT91), .B1(new_n653), .B2(new_n375), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT91), .ZN(new_n655));
  INV_X1    g0455(.A(new_n652), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n437), .B1(new_n433), .B2(new_n396), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n638), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n655), .B(new_n376), .C1(new_n658), .C2(new_n637), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n580), .A2(new_n574), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n627), .A2(new_n320), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n300), .B1(new_n629), .B2(new_n630), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n572), .B(new_n661), .C1(new_n662), .C2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n496), .A2(new_n503), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n541), .A4(new_n633), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n498), .A2(new_n501), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n499), .A2(new_n502), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n541), .A4(new_n536), .ZN(new_n671));
  XNOR2_X1  g0471(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n533), .A2(new_n514), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n541), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n503), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n671), .A2(new_n672), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n668), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n443), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n660), .A2(new_n678), .ZN(G369));
  NOR2_X1   g0479(.A1(new_n388), .A2(new_n257), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT27), .B1(new_n681), .B2(G1), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n683), .A3(new_n264), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT92), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(G343), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT92), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n563), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n572), .A2(new_n661), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n576), .A2(new_n581), .A3(new_n572), .A4(new_n584), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n692), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n662), .A2(new_n665), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n688), .A2(new_n690), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n625), .A2(new_n698), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n626), .A2(new_n633), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n702), .A3(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n691), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n576), .A2(new_n581), .A3(new_n572), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n634), .A2(new_n705), .A3(new_n691), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n213), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n210), .A2(G87), .A3(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n714), .B(new_n715), .C1(new_n236), .C2(new_n710), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n677), .A2(new_n718), .A3(new_n691), .ZN(new_n719));
  INV_X1    g0519(.A(new_n673), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n671), .A2(new_n672), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n626), .A2(new_n572), .A3(new_n576), .A4(new_n581), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n667), .A3(new_n541), .A4(new_n633), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n698), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n719), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n485), .A2(new_n320), .A3(new_n570), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n627), .A2(new_n530), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT96), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n485), .A2(new_n320), .A3(new_n570), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n627), .A2(new_n530), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT96), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n472), .A2(new_n477), .A3(new_n484), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n532), .A2(new_n570), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n736), .A2(new_n599), .A3(new_n737), .A4(KEYINPUT30), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT94), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n594), .A2(new_n598), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n485), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT94), .A3(KEYINPUT30), .A4(new_n737), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n737), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT95), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n494), .A2(new_n477), .A3(new_n598), .A4(new_n594), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n532), .A2(new_n570), .ZN(new_n749));
  OAI211_X1 g0549(.A(KEYINPUT95), .B(new_n746), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n735), .B(new_n744), .C1(new_n747), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT97), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n750), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(KEYINPUT97), .A3(new_n735), .A4(new_n744), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n754), .A2(new_n698), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n635), .A2(new_n691), .ZN(new_n763));
  INV_X1    g0563(.A(new_n744), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n755), .B1(new_n732), .B2(new_n733), .ZN(new_n765));
  OAI211_X1 g0565(.A(KEYINPUT31), .B(new_n698), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n727), .B1(G330), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n717), .B1(new_n768), .B2(G1), .ZN(G364));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n696), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n234), .B1(G20), .B2(new_n300), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n255), .A2(G45), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n708), .A2(new_n356), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n236), .B2(G45), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n777), .A2(new_n779), .B1(G116), .B2(new_n213), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n356), .A2(new_n213), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G87), .B2(new_n210), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n776), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n435), .A2(G179), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G20), .A3(G190), .ZN(new_n785));
  INV_X1    g0585(.A(G303), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n233), .A2(new_n320), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT98), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n331), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n790), .A2(new_n435), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G322), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n790), .A2(new_n364), .A3(new_n435), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G311), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n233), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n388), .A2(new_n364), .A3(new_n784), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n788), .A2(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G190), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n364), .A2(G179), .A3(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n233), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n356), .B1(new_n809), .B2(G294), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n794), .A2(new_n797), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n803), .A2(new_n331), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n787), .B(new_n811), .C1(G326), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n798), .A2(G159), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(KEYINPUT32), .ZN(new_n815));
  INV_X1    g0615(.A(new_n804), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n816), .B2(new_n203), .ZN(new_n817));
  INV_X1    g0617(.A(new_n785), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G87), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n793), .A2(G58), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n809), .A2(G97), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n796), .A2(G77), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n801), .A2(new_n209), .ZN(new_n824));
  INV_X1    g0624(.A(new_n812), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n356), .B1(KEYINPUT32), .B2(new_n814), .C1(new_n825), .C2(new_n253), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n775), .B1(new_n813), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n264), .B1(new_n680), .B2(G45), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n709), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n774), .A2(new_n783), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n696), .A2(G330), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n696), .A2(G330), .ZN(new_n834));
  INV_X1    g0634(.A(new_n831), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n836), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n698), .A2(new_n395), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n441), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n396), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n644), .A2(new_n691), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n677), .A2(new_n691), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n677), .A2(KEYINPUT101), .A3(new_n691), .A4(new_n843), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n677), .A2(new_n691), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n842), .ZN(new_n850));
  INV_X1    g0650(.A(G330), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n760), .A2(new_n761), .B1(new_n635), .B2(new_n691), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n766), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT102), .Z(new_n855));
  AOI21_X1  g0655(.A(new_n831), .B1(new_n850), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n793), .A2(G143), .B1(G150), .B2(new_n804), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n859), .B2(new_n825), .C1(new_n283), .C2(new_n795), .ZN(new_n860));
  XNOR2_X1  g0660(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n202), .A2(new_n808), .B1(new_n801), .B2(new_n203), .ZN(new_n863));
  INV_X1    g0663(.A(new_n798), .ZN(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n356), .B1(new_n253), .B2(new_n785), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n795), .A2(new_n547), .B1(new_n800), .B2(new_n816), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n356), .B1(new_n868), .B2(KEYINPUT99), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n869), .B1(new_n209), .B2(new_n785), .C1(new_n786), .C2(new_n825), .ZN(new_n870));
  INV_X1    g0670(.A(G311), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n801), .A2(new_n223), .ZN(new_n873));
  INV_X1    g0673(.A(G294), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n821), .B1(new_n874), .B2(new_n792), .C1(new_n868), .C2(KEYINPUT99), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n870), .A2(new_n872), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n775), .B1(new_n867), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n775), .A2(new_n770), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n392), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n842), .A2(new_n770), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n877), .A2(new_n831), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n857), .A2(new_n881), .ZN(G384));
  INV_X1    g0682(.A(new_n841), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n846), .B2(new_n847), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n432), .A2(new_n698), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n433), .A2(new_n438), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n432), .B(new_n698), .C1(new_n437), .C2(new_n418), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n288), .A2(new_n289), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n340), .A3(new_n263), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n266), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n686), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n299), .A2(new_n327), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n649), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n299), .A2(new_n327), .A3(KEYINPUT18), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n899), .B2(new_n638), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n646), .B1(new_n893), .B2(new_n266), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n895), .A3(new_n334), .ZN(new_n903));
  INV_X1    g0703(.A(new_n334), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n685), .B1(new_n341), .B2(new_n266), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT37), .B1(new_n299), .B2(new_n327), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n903), .A2(KEYINPUT37), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n891), .B1(new_n900), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n685), .B1(new_n893), .B2(new_n266), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n330), .B2(new_n343), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n299), .A2(new_n686), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n334), .A3(new_n912), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n904), .A2(new_n901), .A3(new_n910), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n890), .A2(new_n918), .B1(new_n656), .B2(new_n685), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n433), .A2(new_n698), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n912), .B1(new_n652), .B2(new_n638), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n648), .A2(new_n912), .A3(new_n334), .ZN(new_n924));
  AOI22_X1  g0724(.A1(KEYINPUT37), .A2(new_n924), .B1(new_n906), .B2(new_n907), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n891), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n927), .A3(new_n917), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT103), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n918), .A2(KEYINPUT39), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT103), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n926), .A2(new_n917), .A3(new_n931), .A4(new_n927), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT104), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n929), .A2(new_n930), .A3(new_n935), .A4(new_n932), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n922), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n920), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n443), .A2(new_n727), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n660), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n698), .A4(new_n759), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n762), .A2(new_n763), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n842), .B1(new_n886), .B2(new_n887), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n926), .B2(new_n917), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n943), .A2(new_n918), .A3(new_n944), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n945), .A2(new_n947), .B1(new_n948), .B2(new_n946), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n443), .A2(new_n943), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(G330), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n941), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n264), .B2(new_n680), .ZN(new_n954));
  INV_X1    g0754(.A(new_n452), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n547), .B1(new_n955), .B2(KEYINPUT35), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(new_n235), .C1(KEYINPUT35), .C2(new_n955), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT36), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n277), .A2(G77), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n236), .A2(new_n959), .B1(G50), .B2(new_n203), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n257), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n958), .A3(new_n961), .ZN(G367));
  OAI22_X1  g0762(.A1(new_n795), .A2(new_n253), .B1(new_n202), .B2(new_n785), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n864), .A2(new_n859), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n801), .A2(new_n392), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n812), .A2(G143), .B1(G68), .B2(new_n809), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n966), .A2(new_n356), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(G150), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n968), .B1(new_n969), .B2(new_n792), .C1(new_n283), .C2(new_n816), .ZN(new_n970));
  INV_X1    g0770(.A(new_n567), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n792), .A2(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n795), .A2(new_n800), .B1(new_n209), .B2(new_n808), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n973), .A2(new_n974), .B1(G294), .B2(new_n804), .ZN(new_n975));
  INV_X1    g0775(.A(new_n801), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(G97), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n975), .B(new_n977), .C1(new_n978), .C2(new_n864), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT111), .B(G311), .Z(new_n980));
  AOI211_X1 g0780(.A(new_n972), .B(new_n979), .C1(new_n812), .C2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n973), .A2(new_n974), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n269), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT112), .B1(new_n818), .B2(G116), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT46), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n970), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT47), .Z(new_n987));
  INV_X1    g0787(.A(new_n775), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n778), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n776), .B1(new_n213), .B2(new_n511), .C1(new_n246), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n537), .A2(new_n540), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n698), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(new_n541), .A3(new_n673), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n673), .B2(new_n993), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n831), .B(new_n991), .C1(new_n995), .C2(new_n773), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n989), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n705), .A2(new_n691), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(new_n699), .A3(new_n701), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n706), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(new_n834), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT107), .B1(new_n768), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT107), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n853), .A2(new_n727), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n706), .A2(new_n704), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  OR3_X1    g0810(.A1(new_n691), .A2(new_n503), .A3(KEYINPUT105), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT105), .B1(new_n691), .B2(new_n503), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n698), .A2(new_n499), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1011), .A2(new_n1012), .B1(new_n667), .B2(new_n1013), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1009), .A2(new_n1010), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1010), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1014), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1018), .A2(KEYINPUT45), .A3(new_n704), .A4(new_n706), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT45), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1017), .A2(new_n703), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n703), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n999), .B1(new_n1008), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n767), .A2(G330), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n727), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1006), .B1(new_n1029), .B2(new_n1003), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n768), .A2(KEYINPUT107), .A3(new_n1004), .ZN(new_n1031));
  AND4_X1   g0831(.A1(new_n999), .A2(new_n1030), .A3(new_n1025), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n768), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n830), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT109), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT106), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n703), .A2(new_n1014), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  NAND2_X1  g0840(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1014), .A2(new_n706), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT42), .Z(new_n1043));
  NAND2_X1  g0843(.A1(new_n1018), .A2(new_n697), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n698), .B1(new_n1044), .B2(new_n503), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1041), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1040), .B(new_n1046), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1035), .A2(new_n1036), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1008), .A2(new_n999), .A3(new_n1025), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1030), .A2(new_n1025), .A3(new_n1031), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT108), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1029), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1034), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n829), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1047), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT109), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n998), .B1(new_n1048), .B2(new_n1056), .ZN(G387));
  OAI22_X1  g0857(.A1(new_n978), .A2(new_n792), .B1(new_n795), .B2(new_n971), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT113), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n812), .A2(G322), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n804), .A2(new_n980), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT48), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n809), .A2(G283), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n818), .A2(G294), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1064), .A2(new_n1069), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n356), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n798), .A2(G326), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n547), .C2(new_n801), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n796), .A2(G68), .B1(G150), .B2(new_n798), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n260), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n816), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n785), .A2(new_n392), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n511), .A2(new_n808), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n792), .A2(new_n253), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n812), .A2(G159), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1080), .A2(new_n356), .A3(new_n977), .A4(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n988), .B1(new_n1073), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(G45), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n778), .B1(new_n242), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n711), .B2(new_n781), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n260), .A2(new_n253), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT50), .Z(new_n1088));
  NAND2_X1  g0888(.A1(G68), .A2(G77), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1088), .A2(new_n1084), .A3(new_n1089), .A4(new_n711), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n708), .A2(new_n209), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n772), .B(new_n775), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n702), .A2(new_n773), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1083), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1095), .A2(new_n831), .B1(new_n830), .B2(new_n1004), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1008), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n709), .C1(new_n768), .C2(new_n1004), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(G393));
  INV_X1    g0899(.A(new_n1025), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n709), .B(new_n1101), .C1(new_n1026), .C2(new_n1032), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1025), .A2(new_n830), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n792), .A2(new_n871), .B1(new_n978), .B2(new_n825), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  AOI211_X1 g0905(.A(new_n824), .B(new_n1105), .C1(G294), .C2(new_n796), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n808), .A2(new_n547), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n356), .B(new_n1107), .C1(G322), .C2(new_n798), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(new_n971), .C2(new_n816), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G283), .B2(new_n818), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n798), .A2(G143), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n253), .B2(new_n816), .C1(new_n795), .C2(new_n1075), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT51), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n792), .A2(new_n283), .B1(new_n969), .B2(new_n825), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .C1(new_n392), .C2(new_n808), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n785), .A2(new_n203), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1116), .A2(new_n269), .A3(new_n873), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n775), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1014), .A2(new_n772), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n251), .A2(new_n778), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n776), .C1(new_n208), .C2(new_n213), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n831), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1102), .A2(new_n1103), .A3(new_n1123), .ZN(G390));
  AOI21_X1  g0924(.A(new_n888), .B1(new_n853), .B2(new_n843), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n943), .A2(G330), .A3(new_n944), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1125), .A2(new_n1127), .B1(new_n883), .B2(new_n848), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n853), .A2(new_n843), .A3(new_n888), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n943), .A2(G330), .A3(new_n843), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n889), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n883), .B1(new_n726), .B2(new_n840), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n443), .A2(G330), .A3(new_n943), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n660), .A2(new_n939), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n922), .B1(new_n884), .B2(new_n889), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n936), .A3(new_n934), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n921), .B1(new_n917), .B2(new_n926), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n889), .B2(new_n1132), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1126), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1129), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1139), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1137), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT114), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1137), .A2(new_n1143), .A3(KEYINPUT114), .A4(new_n1145), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n660), .A2(new_n939), .A3(new_n1135), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1139), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1127), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1148), .A2(new_n709), .A3(new_n1149), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n830), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT115), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n934), .A2(new_n770), .A3(new_n936), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n878), .A2(new_n1075), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n792), .A2(new_n865), .B1(new_n1161), .B2(new_n825), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT116), .Z(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT54), .B(G143), .Z(new_n1164));
  AOI211_X1 g0964(.A(new_n269), .B(new_n1163), .C1(new_n796), .C2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n283), .B2(new_n808), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n816), .A2(new_n859), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n818), .A2(G150), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n798), .A2(G125), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n253), .B2(new_n801), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .A4(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n793), .A2(G116), .B1(G87), .B2(new_n818), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G77), .A2(new_n809), .B1(new_n976), .B2(G68), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n208), .C2(new_n795), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n816), .A2(new_n209), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n825), .A2(new_n800), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n269), .B1(new_n864), .B2(new_n874), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n775), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1159), .A2(new_n831), .A3(new_n1160), .A4(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1155), .A2(new_n1158), .A3(new_n1181), .ZN(G378));
  NAND2_X1  g0982(.A1(new_n1154), .A2(new_n1136), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n948), .A2(new_n946), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(G330), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT118), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n372), .A2(new_n376), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT117), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT117), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n372), .A2(new_n1190), .A3(new_n376), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n354), .A2(new_n685), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1189), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1190), .B1(new_n372), .B2(new_n376), .ZN(new_n1195));
  AOI211_X1 g0995(.A(KEYINPUT117), .B(new_n375), .C1(new_n370), .C2(new_n371), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1192), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1198), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1187), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1186), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n1184), .A3(G330), .A4(new_n1185), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n934), .A2(new_n936), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n921), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n919), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1204), .A2(new_n1208), .A3(new_n1205), .A4(new_n919), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1212), .ZN(new_n1213));
  AND4_X1   g1013(.A1(new_n1208), .A2(new_n1204), .A3(new_n919), .A4(new_n1205), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1205), .A2(new_n1204), .B1(new_n1208), .B2(new_n919), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT119), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT119), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1211), .A2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1216), .A2(new_n1218), .B1(new_n1136), .B2(new_n1154), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n709), .B(new_n1213), .C1(new_n1219), .C2(KEYINPUT57), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G50), .B1(new_n273), .B2(new_n473), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G41), .B1(new_n798), .B2(G124), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1164), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n785), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n795), .A2(new_n859), .B1(new_n969), .B2(new_n808), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(G125), .C2(new_n812), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n1161), .B2(new_n792), .C1(new_n865), .C2(new_n816), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n348), .B(new_n1222), .C1(new_n1227), .C2(KEYINPUT59), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G159), .B2(new_n976), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1221), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n976), .A2(G58), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n800), .B2(new_n864), .C1(new_n795), .C2(new_n511), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1077), .B(new_n1234), .C1(G107), .C2(new_n793), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n269), .B1(new_n816), .B2(new_n208), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G41), .B(new_n1236), .C1(G116), .C2(new_n812), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1235), .B(new_n1237), .C1(new_n203), .C2(new_n808), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT58), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n988), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1201), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n771), .B1(new_n1241), .B2(new_n1199), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n878), .A2(new_n253), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(new_n1240), .A2(new_n1242), .A3(new_n835), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n830), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1220), .A2(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n878), .A2(new_n203), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1233), .B1(new_n283), .B2(new_n785), .C1(new_n795), .C2(new_n969), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G132), .B2(new_n812), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n859), .B2(new_n792), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n269), .B(new_n1252), .C1(G128), .C2(new_n798), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n253), .B2(new_n808), .C1(new_n816), .C2(new_n1223), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n965), .B1(new_n812), .B2(G294), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n511), .B2(new_n808), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n269), .B1(new_n547), .B2(new_n816), .C1(new_n792), .C2(new_n800), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(G303), .C2(new_n798), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1258), .B1(new_n208), .B2(new_n785), .C1(new_n209), .C2(new_n795), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n988), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n888), .A2(new_n771), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1260), .A2(new_n835), .A3(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1134), .A2(new_n830), .B1(new_n1249), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1128), .A2(new_n1150), .A3(new_n1133), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1034), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1265), .B2(new_n1151), .ZN(G381));
  OAI21_X1  g1066(.A(new_n1036), .B1(new_n1035), .B2(new_n1047), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1054), .A2(KEYINPUT109), .A3(new_n1055), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G390), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n998), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G396), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1096), .A2(new_n1272), .A3(new_n1098), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G384), .A2(new_n1271), .A3(G381), .A4(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1274), .A2(KEYINPUT120), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G375), .A2(G378), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(KEYINPUT120), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(G407));
  NAND2_X1  g1078(.A1(new_n689), .A2(G213), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(KEYINPUT121), .Z(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G407), .A2(G213), .A3(new_n1282), .ZN(G409));
  AND3_X1   g1083(.A1(new_n1096), .A2(new_n1272), .A3(new_n1098), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1272), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT125), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1273), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1270), .B1(new_n1269), .B2(new_n998), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n997), .B(G390), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(G390), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1271), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT122), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1220), .A2(G378), .A3(new_n1247), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1217), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1218), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1183), .B(new_n1034), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1245), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1212), .A2(new_n830), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1306), .A2(new_n1155), .A3(new_n1181), .A4(new_n1158), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1300), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1279), .ZN(new_n1309));
  INV_X1    g1109(.A(G384), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT60), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1264), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1264), .A2(new_n1311), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1312), .A2(new_n709), .A3(new_n1137), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1263), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(G384), .A3(new_n1263), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1299), .B1(new_n1309), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1279), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1300), .B2(new_n1307), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1318), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(KEYINPUT122), .A3(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1320), .A3(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1308), .A2(new_n1280), .A3(new_n1323), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1326), .B2(KEYINPUT62), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1318), .A2(new_n1281), .ZN(new_n1329));
  INV_X1    g1129(.A(G2897), .ZN(new_n1330));
  OR2_X1    g1130(.A1(new_n1330), .A2(KEYINPUT124), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(KEYINPUT124), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1321), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  OAI22_X1  g1134(.A1(new_n1329), .A2(new_n1330), .B1(new_n1318), .B2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(new_n1280), .B2(new_n1308), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1298), .B1(new_n1328), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT123), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1322), .A2(new_n1338), .ZN(new_n1339));
  AOI211_X1 g1139(.A(KEYINPUT123), .B(new_n1321), .C1(new_n1300), .C2(new_n1307), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1335), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1308), .A2(KEYINPUT63), .A3(new_n1323), .A4(new_n1280), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1297), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1341), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  AND4_X1   g1146(.A1(KEYINPUT122), .A2(new_n1308), .A3(new_n1279), .A4(new_n1323), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT122), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1346), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT126), .B1(new_n1345), .B2(new_n1349), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1297), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1309), .A2(KEYINPUT123), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1335), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1322), .A2(new_n1338), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  AND4_X1   g1155(.A1(KEYINPUT126), .A2(new_n1349), .A3(new_n1351), .A4(new_n1355), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1337), .B1(new_n1350), .B2(new_n1356), .ZN(G405));
  XNOR2_X1  g1157(.A(G375), .B(G378), .ZN(new_n1358));
  XNOR2_X1  g1158(.A(new_n1358), .B(new_n1323), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1359), .B(new_n1297), .ZN(G402));
endmodule


