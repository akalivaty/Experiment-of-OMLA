//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  XNOR2_X1  g0043(.A(KEYINPUT8), .B(G58), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n245), .A2(new_n247), .B1(G150), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n249), .A2(KEYINPUT65), .B1(G20), .B2(new_n203), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(KEYINPUT65), .B2(new_n249), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n216), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n206), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n256), .B(KEYINPUT66), .Z(new_n257));
  NAND3_X1  g0057(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(new_n216), .A3(new_n252), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n258), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n257), .A2(new_n260), .B1(new_n202), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n246), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(G223), .B1(new_n273), .B2(G77), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n268), .A2(new_n269), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G222), .A3(new_n266), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n265), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(new_n265), .A3(G274), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n265), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n263), .B(new_n288), .C1(G179), .C2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(G232), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n266), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n266), .A2(G238), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n273), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n216), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n275), .B2(G107), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n265), .A2(G244), .A3(new_n283), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n281), .A2(new_n299), .ZN(new_n300));
  OR3_X1    g0100(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(G200), .B1(new_n297), .B2(new_n300), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G20), .A2(G77), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n207), .A2(G33), .ZN(new_n305));
  INV_X1    g0105(.A(new_n248), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n303), .B1(new_n304), .B2(new_n305), .C1(new_n244), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n307), .A2(new_n253), .B1(new_n308), .B2(new_n261), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n255), .A2(G77), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n259), .A2(KEYINPUT67), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT67), .B1(new_n259), .B2(new_n310), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n301), .A2(new_n302), .A3(new_n309), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n313), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n297), .A2(new_n300), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n287), .B1(new_n297), .B2(new_n300), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n286), .A2(new_n298), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G200), .B2(new_n286), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT9), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n254), .A2(new_n325), .A3(new_n262), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n254), .B2(new_n262), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n323), .B(new_n324), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n326), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n324), .B1(new_n332), .B2(new_n323), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n289), .B(new_n321), .C1(new_n330), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n268), .A2(new_n207), .A3(new_n269), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n269), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G58), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n336), .ZN(new_n343));
  OAI21_X1  g0143(.A(G20), .B1(new_n343), .B2(new_n201), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n248), .A2(G159), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n335), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n253), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n339), .A2(new_n340), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n346), .B1(new_n351), .B2(G68), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n352), .B2(KEYINPUT16), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT71), .B(new_n335), .C1(new_n341), .C2(new_n346), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n245), .A2(new_n255), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n356), .A2(new_n259), .B1(new_n258), .B2(new_n245), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n282), .A2(G1698), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n360), .B1(G223), .B2(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G87), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n265), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n281), .B1(new_n290), .B2(new_n284), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G179), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n287), .B2(new_n365), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT18), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n361), .A2(new_n362), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n295), .ZN(new_n371));
  INV_X1    g0171(.A(new_n364), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n287), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n363), .A2(new_n364), .A3(new_n317), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n355), .B2(new_n358), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n365), .A2(new_n298), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G200), .B2(new_n365), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n355), .A2(new_n358), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n355), .A2(KEYINPUT17), .A3(new_n380), .A4(new_n358), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n369), .A2(new_n378), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n334), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n261), .A2(new_n336), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT12), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n336), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n308), .B2(new_n305), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n260), .A2(G68), .A3(new_n255), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT11), .B1(new_n390), .B2(new_n253), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n265), .A2(G238), .A3(new_n283), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT69), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n281), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n281), .B2(new_n397), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n282), .A2(new_n266), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n290), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n271), .C2(new_n272), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(KEYINPUT68), .A3(new_n405), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n295), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT13), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n401), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n401), .B2(new_n410), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n396), .B(G169), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n408), .A2(new_n409), .A3(new_n295), .ZN(new_n415));
  INV_X1    g0215(.A(new_n400), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n281), .A2(new_n397), .A3(new_n398), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT13), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n401), .A2(new_n410), .A3(new_n411), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(G179), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n420), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n396), .B1(new_n423), .B2(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT70), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n412), .A2(new_n413), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT14), .B1(new_n426), .B2(new_n287), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT70), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n421), .A4(new_n414), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n395), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n423), .A2(G200), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n395), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n386), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g0236(.A(KEYINPUT78), .B(KEYINPUT21), .Z(new_n437));
  NOR2_X1   g0237(.A1(new_n261), .A2(G116), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n350), .B(new_n258), .C1(G1), .C2(new_n246), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(G116), .ZN(new_n440));
  AOI21_X1  g0240(.A(G20), .B1(new_n246), .B2(G97), .ZN(new_n441));
  INV_X1    g0241(.A(G283), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n246), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G116), .ZN(new_n444));
  AOI221_X4 g0244(.A(KEYINPUT76), .B1(new_n444), .B2(G20), .C1(new_n252), .C2(new_n216), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(G20), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n253), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n443), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT20), .B(new_n443), .C1(new_n445), .C2(new_n448), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n440), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n279), .A2(G1), .ZN(new_n454));
  NAND2_X1  g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G274), .B1(new_n294), .B2(new_n216), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT72), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n206), .A2(G45), .ZN(new_n462));
  OR2_X1    g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n455), .ZN(new_n464));
  INV_X1    g0264(.A(G274), .ZN(new_n465));
  AND2_X1   g0265(.A1(G1), .A2(G13), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n264), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT72), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n266), .A2(G264), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G257), .A2(G1698), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n470), .A2(new_n471), .B1(new_n271), .B2(new_n272), .ZN(new_n472));
  INV_X1    g0272(.A(G303), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n268), .A2(new_n473), .A3(new_n269), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n295), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n458), .A2(G270), .A3(new_n265), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(G169), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n437), .B1(new_n453), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n437), .C1(new_n453), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n253), .A2(new_n447), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT76), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n253), .A2(new_n446), .A3(new_n447), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT20), .B1(new_n487), .B2(new_n443), .ZN(new_n488));
  INV_X1    g0288(.A(new_n452), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n259), .B1(new_n206), .B2(G33), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n444), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n488), .A2(new_n489), .B1(new_n491), .B2(new_n438), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n469), .A2(new_n317), .A3(new_n477), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(KEYINPUT77), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT77), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n475), .A2(new_n476), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n460), .B1(new_n458), .B2(new_n459), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n464), .A2(KEYINPUT72), .A3(new_n467), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(G179), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n495), .B1(new_n453), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n453), .A2(new_n478), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n494), .A2(new_n501), .B1(new_n502), .B2(KEYINPUT21), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  INV_X1    g0305(.A(G107), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(G20), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n507), .C1(new_n444), .C2(new_n305), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT80), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n247), .A2(G116), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(KEYINPUT80), .A3(new_n507), .A4(new_n504), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n207), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT22), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n275), .A2(new_n517), .A3(new_n207), .A4(G87), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n513), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n514), .B1(new_n513), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n253), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT25), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n258), .B2(G107), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n258), .A2(new_n523), .A3(G107), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n439), .A2(new_n506), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G250), .B(new_n266), .C1(new_n271), .C2(new_n272), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  OAI211_X1 g0331(.A(G257), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT81), .B1(new_n270), .B2(G257), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n295), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n458), .A2(G264), .A3(new_n265), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(new_n537), .A3(new_n499), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n458), .A2(KEYINPUT82), .A3(G264), .A4(new_n265), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n542), .A3(new_n499), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n538), .A2(new_n287), .B1(new_n543), .B2(new_n317), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n529), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n483), .A2(new_n503), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n207), .B1(new_n405), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  INV_X1    g0349(.A(G87), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n207), .B(G68), .C1(new_n271), .C2(new_n272), .ZN(new_n553));
  INV_X1    g0353(.A(G97), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n547), .B1(new_n305), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n253), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT15), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n561), .A2(new_n258), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n557), .A2(KEYINPUT75), .A3(new_n563), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n490), .A2(G87), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT74), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT74), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n275), .A2(new_n572), .A3(G244), .A4(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G238), .B(new_n266), .C1(new_n271), .C2(new_n272), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G116), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n265), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(G250), .B1(new_n206), .B2(G45), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n295), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G274), .B2(new_n462), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(G200), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n575), .A2(new_n576), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n573), .B2(new_n571), .ZN(new_n585));
  OAI211_X1 g0385(.A(G190), .B(new_n581), .C1(new_n585), .C2(new_n265), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n568), .A2(new_n569), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n490), .A2(new_n561), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT75), .B1(new_n557), .B2(new_n563), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n565), .B(new_n562), .C1(new_n556), .C2(new_n253), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n581), .B1(new_n585), .B2(new_n265), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n287), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n317), .B(new_n581), .C1(new_n585), .C2(new_n265), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g0396(.A(KEYINPUT5), .B(G41), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n454), .B1(new_n466), .B2(new_n264), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G257), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n461), .B2(new_n468), .ZN(new_n600));
  OAI211_X1 g0400(.A(G244), .B(new_n266), .C1(new_n271), .C2(new_n272), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n246), .A2(new_n442), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G250), .A2(G1698), .ZN(new_n605));
  NAND2_X1  g0405(.A1(KEYINPUT4), .A2(G244), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n275), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n265), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n600), .A2(KEYINPUT73), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT73), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n497), .A2(new_n498), .B1(new_n598), .B2(G257), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n603), .A2(new_n608), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n295), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n287), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n600), .A2(new_n609), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n506), .A2(KEYINPUT6), .A3(G97), .ZN(new_n618));
  XNOR2_X1  g0418(.A(G97), .B(G107), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT6), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n621), .A2(new_n207), .B1(new_n308), .B2(new_n306), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n506), .B1(new_n339), .B2(new_n340), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n253), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n258), .A2(G97), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n490), .B2(G97), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n617), .A2(new_n317), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n626), .ZN(new_n628));
  INV_X1    g0428(.A(G200), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n612), .B2(new_n614), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT73), .B1(new_n600), .B2(new_n609), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n612), .A2(new_n614), .A3(new_n611), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G190), .A3(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n616), .A2(new_n627), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n532), .A2(new_n533), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n275), .A2(KEYINPUT81), .A3(G257), .A4(G1698), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n530), .A4(new_n531), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(new_n295), .B1(new_n540), .B2(new_n541), .ZN(new_n639));
  AOI21_X1  g0439(.A(G200), .B1(new_n639), .B2(new_n499), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n298), .A2(new_n536), .A3(new_n537), .A4(new_n499), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n522), .B(new_n528), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(G200), .B1(new_n469), .B2(new_n477), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n496), .A2(G190), .A3(new_n499), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n453), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n596), .A2(new_n635), .A3(new_n642), .A4(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n436), .A2(new_n546), .A3(new_n646), .ZN(G372));
  AND3_X1   g0447(.A1(new_n642), .A2(new_n595), .A3(new_n587), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n546), .A2(new_n648), .A3(new_n635), .ZN(new_n649));
  INV_X1    g0449(.A(new_n595), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n587), .A2(new_n595), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n616), .A2(new_n627), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n612), .A2(new_n614), .A3(new_n317), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n628), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n632), .A2(new_n633), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n287), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n595), .A4(new_n587), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n650), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n436), .B1(new_n649), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n377), .B1(new_n359), .B2(new_n367), .ZN(new_n662));
  AOI211_X1 g0462(.A(KEYINPUT18), .B(new_n375), .C1(new_n355), .C2(new_n358), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n425), .A2(new_n429), .ZN(new_n666));
  INV_X1    g0466(.A(new_n395), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n434), .B2(new_n320), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n383), .A2(new_n384), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n330), .A2(new_n333), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n289), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n661), .A2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n483), .A2(new_n503), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(G213), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n453), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n676), .B(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n645), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n545), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n529), .A2(new_n682), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n642), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n545), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n682), .B1(new_n483), .B2(new_n503), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n689), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n210), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n549), .A2(new_n550), .A3(new_n444), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT83), .Z(new_n701));
  OR3_X1    g0501(.A1(new_n699), .A2(new_n701), .A3(new_n206), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT84), .ZN(new_n703));
  INV_X1    g0503(.A(new_n699), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n702), .A2(new_n703), .B1(new_n214), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n703), .B2(new_n702), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT28), .Z(new_n707));
  INV_X1    g0507(.A(KEYINPUT88), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n660), .A2(new_n649), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n683), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n649), .A2(KEYINPUT87), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n596), .A2(new_n635), .A3(new_n642), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT87), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n546), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n716), .A3(new_n660), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n683), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(new_n708), .A3(KEYINPUT29), .A4(new_n683), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n536), .A2(new_n542), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n722), .A2(new_n592), .A3(new_n500), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n610), .A2(new_n615), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT30), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(G179), .B1(new_n496), .B2(new_n499), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n612), .A2(new_n614), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n543), .A2(new_n726), .A3(new_n727), .A4(new_n592), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n632), .A2(KEYINPUT30), .A3(new_n633), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n572), .B1(new_n270), .B2(G244), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n570), .A2(KEYINPUT74), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n577), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n582), .B1(new_n732), .B2(new_n295), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n493), .A2(new_n733), .A3(new_n639), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n728), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT31), .B(new_n682), .C1(new_n725), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(KEYINPUT85), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n682), .B1(new_n725), .B2(new_n735), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT86), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT86), .A3(new_n740), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n743), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n745), .A2(new_n741), .B1(KEYINPUT85), .B2(new_n737), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n483), .A2(new_n545), .A3(new_n503), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n714), .A2(new_n747), .A3(new_n645), .A4(new_n683), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n721), .B1(G330), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n707), .B1(new_n750), .B2(G1), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT89), .ZN(G364));
  AND2_X1   g0552(.A1(new_n207), .A2(G13), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n206), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n699), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n698), .A2(new_n275), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n279), .B2(new_n215), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n279), .B2(new_n239), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n698), .A2(new_n273), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(G355), .B1(new_n444), .B2(new_n698), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT90), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n216), .B1(G20), .B2(new_n287), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n757), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n768), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n207), .A2(new_n629), .A3(G179), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(new_n298), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(new_n317), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n298), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n317), .A2(G200), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(G20), .A3(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(new_n783), .B2(G322), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n776), .A2(new_n442), .B1(KEYINPUT94), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(KEYINPUT94), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n207), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G179), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n781), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n273), .B1(new_n789), .B2(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n772), .A2(G190), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n207), .B1(new_n788), .B2(G190), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n794), .A2(new_n473), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n798), .A2(KEYINPUT91), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(KEYINPUT91), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT93), .B(G326), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n793), .B(new_n797), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n789), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT32), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n550), .B2(new_n794), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n275), .B1(new_n792), .B2(new_n308), .C1(new_n342), .C2(new_n782), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n806), .A2(new_n807), .B1(new_n336), .B2(new_n778), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n796), .A2(new_n554), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n776), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n814), .A2(G107), .B1(G50), .B2(new_n802), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n786), .A2(new_n804), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n767), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n770), .B1(new_n771), .B2(new_n816), .C1(new_n686), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n688), .A2(new_n756), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n686), .A2(G330), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n749), .A2(G330), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n315), .A2(new_n682), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n314), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n320), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n320), .A2(new_n682), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT99), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n710), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n828), .B(KEYINPUT99), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n709), .A2(new_n683), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n823), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT100), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n823), .A2(new_n834), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT101), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n756), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n836), .B(new_n841), .C1(new_n838), .C2(new_n837), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n768), .A2(new_n765), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n756), .B1(G77), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n789), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n273), .B1(new_n845), .B2(G132), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n814), .A2(G68), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n202), .B2(new_n794), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT97), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n846), .B1(new_n342), .B2(new_n796), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n852), .A2(KEYINPUT98), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(KEYINPUT98), .ZN(new_n854));
  XNOR2_X1  g0654(.A(KEYINPUT95), .B(G143), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n792), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n783), .A2(new_n856), .B1(new_n857), .B2(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n859), .B2(new_n778), .C1(new_n801), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT96), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n853), .A2(new_n854), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n814), .A2(G87), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n792), .A2(new_n444), .B1(new_n789), .B2(new_n791), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n275), .B(new_n866), .C1(G294), .C2(new_n783), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n778), .A2(new_n442), .ZN(new_n868));
  INV_X1    g0668(.A(new_n794), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n812), .B(new_n868), .C1(G107), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n802), .A2(G303), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n865), .A2(new_n867), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n844), .B1(new_n873), .B2(new_n768), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n766), .B2(new_n832), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n842), .A2(new_n875), .ZN(G384));
  INV_X1    g0676(.A(new_n621), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n217), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  OR3_X1    g0681(.A1(new_n214), .A2(new_n308), .A3(new_n343), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n202), .A2(G68), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n206), .B(G13), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n436), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT30), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n734), .B2(new_n657), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n888), .B(new_n728), .C1(new_n734), .C2(new_n729), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT31), .B1(new_n889), .B2(new_n682), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n737), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n748), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT104), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  INV_X1    g0695(.A(new_n680), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n359), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n368), .A2(new_n897), .A3(new_n381), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT103), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n368), .A2(new_n897), .A3(new_n901), .A4(new_n381), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n680), .B1(new_n355), .B2(new_n358), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n385), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n898), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n352), .A2(KEYINPUT16), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n910), .A2(new_n253), .A3(new_n347), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(new_n357), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n896), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n385), .A2(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n911), .A2(new_n357), .B1(new_n367), .B2(new_n896), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n381), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n902), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n646), .A2(new_n546), .A3(new_n682), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n739), .A2(new_n740), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n736), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n832), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n395), .A2(new_n683), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n668), .A2(new_n433), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n430), .B2(new_n434), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n895), .B1(new_n921), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n913), .B1(new_n670), .B2(new_n664), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n901), .B1(new_n916), .B2(new_n381), .ZN(new_n933));
  INV_X1    g0733(.A(new_n381), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n934), .A2(new_n376), .A3(new_n904), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(new_n901), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n908), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n920), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n928), .A2(new_n929), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n830), .B1(new_n891), .B2(new_n748), .ZN(new_n940));
  AND4_X1   g0740(.A1(new_n895), .A2(new_n938), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n931), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n894), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n894), .A2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(G330), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n674), .B1(new_n721), .B2(new_n886), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n935), .A2(new_n901), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n950), .A2(KEYINPUT103), .B1(new_n385), .B2(new_n904), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT38), .B1(new_n951), .B2(new_n903), .ZN(new_n952));
  AOI221_X4 g0752(.A(new_n908), .B1(new_n902), .B2(new_n918), .C1(new_n385), .C2(new_n914), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT102), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n430), .A2(new_n955), .A3(new_n683), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n955), .B1(new_n430), .B2(new_n683), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n937), .A2(new_n920), .A3(KEYINPUT39), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n833), .A2(new_n827), .B1(new_n928), .B2(new_n929), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n938), .B1(new_n665), .B2(new_n680), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n948), .B(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n947), .A2(new_n966), .B1(new_n206), .B2(new_n753), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n947), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n885), .B1(new_n967), .B2(new_n968), .ZN(G367));
  NOR2_X1   g0769(.A1(new_n759), .A2(new_n235), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n769), .B1(new_n210), .B2(new_n304), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n756), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n814), .A2(G77), .B1(new_n802), .B2(new_n856), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n792), .A2(new_n202), .B1(new_n789), .B2(new_n860), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n273), .B(new_n974), .C1(G150), .C2(new_n783), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n796), .A2(new_n336), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n778), .A2(new_n805), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(G58), .C2(new_n869), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(G317), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n792), .A2(new_n442), .B1(new_n789), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n275), .B(new_n981), .C1(G303), .C2(new_n783), .ZN(new_n982));
  INV_X1    g0782(.A(new_n796), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n779), .A2(G294), .B1(new_n983), .B2(G107), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n869), .A2(KEYINPUT46), .A3(G116), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT46), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n794), .B2(new_n444), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n982), .A2(new_n984), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n814), .A2(G97), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n791), .B2(new_n801), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n979), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT47), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n972), .B1(new_n992), .B2(new_n768), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n683), .B1(new_n568), .B2(new_n569), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n650), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n652), .B2(new_n994), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(new_n817), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n628), .A2(new_n682), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n635), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n653), .B2(new_n683), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n695), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1001), .B(KEYINPUT105), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(new_n545), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1006), .A2(new_n653), .ZN(new_n1007));
  OAI211_X1 g0807(.A(KEYINPUT107), .B(new_n1004), .C1(new_n1007), .C2(new_n682), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT107), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1004), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n682), .B1(new_n1006), .B2(new_n653), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT108), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1008), .A2(new_n1012), .A3(new_n1016), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n996), .B(KEYINPUT43), .Z(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n693), .B2(new_n1005), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n693), .A2(new_n1005), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1024), .A3(new_n1021), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n699), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(KEYINPUT109), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n696), .A2(new_n1028), .A3(new_n1001), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT45), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1028), .B1(new_n696), .B2(new_n1001), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n696), .A2(new_n1001), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT44), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1037), .A2(new_n688), .A3(new_n692), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n687), .A2(KEYINPUT110), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n692), .B(new_n694), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n750), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1033), .A2(new_n693), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1038), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1027), .B1(new_n1045), .B2(new_n750), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n755), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n998), .B1(new_n1026), .B2(new_n1047), .ZN(G387));
  NOR2_X1   g0848(.A1(new_n1043), .A2(new_n704), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n750), .B2(new_n1041), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n701), .B(KEYINPUT111), .Z(new_n1051));
  OAI21_X1  g0851(.A(new_n279), .B1(new_n336), .B2(new_n308), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n245), .A2(new_n202), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(KEYINPUT50), .B2(new_n1053), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n758), .B1(new_n232), .B2(new_n279), .C1(new_n1051), .C2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n762), .A2(new_n701), .B1(new_n506), .B2(new_n698), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n757), .B1(new_n1058), .B2(new_n769), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n692), .B2(new_n817), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n792), .A2(new_n336), .B1(new_n789), .B2(new_n859), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n273), .B(new_n1061), .C1(G50), .C2(new_n783), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n778), .A2(new_n244), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n794), .A2(new_n308), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n561), .C2(new_n983), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n802), .A2(G159), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n989), .A2(new_n1062), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n783), .A2(G317), .B1(new_n857), .B2(G303), .ZN(new_n1068));
  INV_X1    g0868(.A(G322), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1068), .B1(new_n791), .B2(new_n778), .C1(new_n801), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n869), .A2(G294), .B1(new_n983), .B2(G283), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT112), .Z(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT49), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n275), .B1(new_n845), .B2(new_n803), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n444), .C2(new_n776), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1076), .A2(KEYINPUT49), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1067), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1060), .B1(new_n1081), .B2(new_n768), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1041), .B2(new_n755), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1050), .A2(new_n1083), .ZN(G393));
  NAND2_X1  g0884(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1042), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n699), .A3(new_n1045), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1038), .A2(new_n755), .A3(new_n1044), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n759), .A2(new_n242), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n769), .B1(new_n554), .B2(new_n210), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n756), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n801), .A2(new_n980), .B1(new_n791), .B2(new_n782), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  AOI22_X1  g0893(.A1(new_n869), .A2(G283), .B1(new_n983), .B2(G116), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n473), .B2(new_n778), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n273), .B1(new_n789), .B2(new_n1069), .C1(new_n795), .C2(new_n792), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n506), .B2(new_n776), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n802), .A2(G150), .B1(G159), .B2(new_n783), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n794), .A2(new_n336), .B1(new_n308), .B2(new_n796), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n275), .B1(new_n789), .B2(new_n855), .C1(new_n244), .C2(new_n792), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G50), .C2(new_n779), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n865), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1093), .A2(new_n1098), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1091), .B1(new_n1107), .B2(new_n768), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1005), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n817), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1087), .A2(new_n1088), .A3(new_n1110), .ZN(G390));
  AOI21_X1  g0911(.A(new_n927), .B1(new_n668), .B2(new_n433), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n430), .A2(new_n434), .A3(new_n926), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n892), .A2(G330), .A3(new_n832), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT115), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n928), .A2(KEYINPUT115), .A3(new_n929), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n717), .A2(new_n683), .A3(new_n832), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1118), .A2(new_n1119), .B1(new_n1120), .B2(new_n827), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n958), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(KEYINPUT114), .A3(new_n956), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT114), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n957), .B2(new_n958), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n921), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n833), .A2(new_n827), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n939), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n954), .A2(new_n961), .B1(new_n1129), .B2(new_n959), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1116), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT39), .B1(new_n909), .B2(new_n920), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n937), .A2(KEYINPUT39), .A3(new_n920), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1132), .A2(new_n1133), .B1(new_n960), .B2(new_n963), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n749), .A2(G330), .A3(new_n832), .A4(new_n939), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n1121), .C2(new_n1126), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1118), .A2(new_n1119), .A3(new_n1115), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1138), .A3(new_n827), .A4(new_n1120), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n749), .A2(G330), .A3(new_n832), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1116), .B1(new_n1140), .B2(new_n1114), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1128), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n436), .B1(new_n719), .B2(new_n720), .ZN(new_n1144));
  AND4_X1   g0944(.A1(G330), .A2(new_n386), .A3(new_n435), .A4(new_n892), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1144), .A2(new_n674), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1137), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1131), .A2(new_n1136), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n699), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1131), .A2(new_n755), .A3(new_n1136), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n756), .B1(new_n245), .B2(new_n843), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n273), .B1(new_n794), .B2(new_n550), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT117), .Z(new_n1154));
  NAND2_X1  g0954(.A1(new_n802), .A2(G283), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n782), .A2(new_n444), .B1(new_n792), .B2(new_n554), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n778), .A2(new_n506), .B1(new_n796), .B2(new_n308), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(G294), .C2(new_n845), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n847), .A2(new_n1154), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n275), .B1(new_n776), .B2(new_n202), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT116), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n802), .A2(G128), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n794), .A2(new_n859), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  INV_X1    g0964(.A(G132), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n782), .A2(new_n1165), .B1(new_n789), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n857), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n779), .A2(G137), .B1(new_n983), .B2(G159), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1162), .A2(new_n1164), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1159), .B1(new_n1161), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1152), .B1(new_n1173), .B2(new_n768), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1133), .B1(new_n921), .B2(new_n949), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n766), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1150), .A2(new_n1151), .A3(new_n1176), .ZN(G378));
  NAND2_X1  g0977(.A1(new_n672), .A2(new_n289), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n263), .A2(new_n896), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1180), .B(new_n1181), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1128), .A2(new_n938), .A3(new_n939), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n665), .A2(new_n680), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1175), .B2(new_n960), .ZN(new_n1187));
  OAI21_X1  g0987(.A(G330), .B1(new_n931), .B2(new_n941), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n953), .B1(new_n908), .B2(new_n907), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n940), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT40), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n930), .A2(new_n895), .A3(new_n938), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n946), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(new_n965), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1183), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n965), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(new_n1182), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1145), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT119), .B1(new_n948), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT119), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1144), .A2(new_n1203), .A3(new_n674), .A4(new_n1145), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1149), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(KEYINPUT57), .A3(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1196), .A2(new_n1199), .B1(new_n1149), .B2(new_n1205), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n699), .C1(KEYINPUT57), .C2(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1183), .A2(new_n766), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n756), .B1(G50), .B2(new_n843), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n814), .A2(G58), .B1(G116), .B2(new_n802), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n273), .A2(new_n278), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n792), .A2(new_n304), .B1(new_n789), .B2(new_n442), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G107), .C2(new_n783), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n976), .B(new_n1064), .C1(G97), .C2(new_n779), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1212), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G50), .B1(new_n246), .B2(new_n278), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1217), .A2(KEYINPUT58), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G33), .B(G41), .C1(new_n845), .C2(G124), .ZN(new_n1220));
  INV_X1    g1020(.A(G128), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n782), .A2(new_n1221), .B1(new_n792), .B2(new_n860), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G132), .B2(new_n779), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n869), .A2(new_n1169), .B1(new_n983), .B2(G150), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n1166), .C2(new_n801), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT118), .Z(new_n1226));
  INV_X1    g1026(.A(KEYINPUT59), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1220), .B1(new_n805), .B2(new_n776), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1226), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1219), .B1(KEYINPUT58), .B2(new_n1217), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1211), .B1(new_n1231), .B2(new_n768), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1200), .A2(new_n755), .B1(new_n1210), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1209), .A2(new_n1233), .ZN(G375));
  INV_X1    g1034(.A(new_n1027), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1147), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT120), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n778), .A2(new_n1168), .B1(new_n782), .B2(new_n860), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n802), .B2(G132), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT123), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n275), .B1(new_n789), .B2(new_n1221), .C1(new_n859), .C2(new_n792), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n794), .A2(new_n805), .B1(new_n202), .B2(new_n796), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n814), .C2(G58), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n778), .A2(new_n444), .B1(new_n792), .B2(new_n506), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(KEYINPUT121), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(KEYINPUT121), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n802), .C2(G294), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n273), .B1(new_n473), .B2(new_n789), .C1(new_n794), .C2(new_n554), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n782), .A2(new_n442), .B1(new_n796), .B2(new_n304), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT122), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1250), .B(new_n1252), .C1(G77), .C2(new_n814), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1242), .A2(new_n1245), .B1(new_n1249), .B2(new_n1253), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n756), .B1(G68), .B2(new_n843), .C1(new_n1254), .C2(new_n771), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n765), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1143), .B2(new_n755), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1239), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(G381));
  INV_X1    g1060(.A(G387), .ZN(new_n1261));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  INV_X1    g1062(.A(G396), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1050), .A2(new_n1263), .A3(new_n1083), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(G390), .A2(G384), .A3(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1261), .A2(new_n1262), .A3(new_n1259), .A4(new_n1265), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1266), .A2(G375), .ZN(G407));
  NAND4_X1  g1067(.A1(new_n1209), .A2(new_n681), .A3(new_n1262), .A4(new_n1233), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(G407), .A2(G213), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT124), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT124), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(G407), .A2(new_n1271), .A3(G213), .A4(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(G409));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1264), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(G387), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(new_n1276), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(G390), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G390), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1280), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1278), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1237), .A2(KEYINPUT60), .A3(new_n1147), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n699), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1237), .B1(KEYINPUT60), .B2(new_n1147), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1258), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n875), .A3(new_n842), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G384), .B(new_n1258), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n681), .A2(G213), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(G2897), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1291), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1295), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1208), .A2(new_n1235), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G378), .B1(new_n1299), .B2(new_n1233), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1197), .A2(new_n1182), .A3(new_n1198), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1182), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT57), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1149), .A2(new_n1205), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n699), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1206), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G378), .B(new_n1233), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT125), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1209), .A2(new_n1309), .A3(G378), .A4(new_n1233), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1300), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1298), .B1(new_n1311), .B2(new_n1294), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1311), .A2(new_n1313), .A3(new_n1294), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1286), .B(new_n1312), .C1(new_n1314), .C2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1300), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1313), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1293), .ZN(new_n1322));
  XOR2_X1   g1122(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1285), .B1(new_n1317), .B2(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1312), .A2(new_n1286), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1322), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1314), .A2(KEYINPUT63), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1326), .A2(new_n1328), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1325), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1262), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1318), .A2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1313), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1335), .B(new_n1329), .ZN(G402));
endmodule


