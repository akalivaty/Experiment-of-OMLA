//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  AOI21_X1  g0045(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT67), .B(G223), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT66), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT65), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n249), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT65), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT65), .B1(new_n256), .B2(new_n257), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT66), .A3(G1698), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n248), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G222), .A3(new_n260), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(new_n223), .B2(new_n264), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n246), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n273), .A2(new_n246), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n246), .A2(new_n272), .ZN(new_n276));
  XOR2_X1   g0076(.A(KEYINPUT64), .B(G226), .Z(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G169), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n210), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(KEYINPUT68), .A3(new_n210), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n289), .A2(new_n211), .A3(G1), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT8), .ZN(new_n299));
  INV_X1    g0099(.A(G58), .ZN(new_n300));
  OR3_X1    g0100(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT69), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(KEYINPUT69), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n211), .A2(G33), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n288), .B1(new_n202), .B2(new_n290), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n281), .B(new_n307), .C1(G179), .C2(new_n279), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n296), .A2(new_n306), .A3(new_n310), .A4(new_n311), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n279), .A2(G200), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n269), .A2(G190), .A3(new_n278), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n315), .B2(new_n316), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n308), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n246), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G232), .A3(new_n273), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT77), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n276), .A2(new_n324), .A3(G232), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n275), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT76), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(new_n251), .A3(G33), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n329), .A3(new_n256), .ZN(new_n330));
  OR2_X1    g0130(.A1(G223), .A2(G1698), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(G226), .B2(new_n260), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n330), .A2(new_n332), .B1(new_n253), .B2(new_n219), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n246), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n326), .A2(G179), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n326), .A2(new_n334), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n280), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n300), .A2(new_n217), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n338), .B2(new_n201), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n297), .A2(G159), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n330), .A2(new_n343), .A3(new_n211), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G68), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n330), .B2(new_n211), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT16), .B(new_n342), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n256), .A2(new_n257), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n211), .ZN(new_n349));
  NOR2_X1   g0149(.A1(KEYINPUT7), .A2(G20), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n259), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n341), .B1(new_n351), .B2(G68), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n347), .B(new_n288), .C1(new_n352), .C2(KEYINPUT16), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n303), .B1(new_n292), .B2(G20), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n291), .A2(new_n354), .B1(new_n290), .B2(new_n303), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n337), .A2(new_n356), .A3(KEYINPUT18), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT78), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT78), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n337), .A2(new_n356), .A3(new_n359), .A4(KEYINPUT18), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n337), .A2(new_n356), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT18), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n326), .A2(G190), .A3(new_n334), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n326), .B2(new_n334), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n365), .B1(new_n369), .B2(new_n356), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n366), .A2(new_n368), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n371), .A2(KEYINPUT17), .A3(new_n353), .A4(new_n355), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n364), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n291), .A2(G77), .A3(new_n293), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G20), .A2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  INV_X1    g0177(.A(new_n297), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT8), .B(G58), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n376), .B1(new_n377), .B2(new_n304), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n288), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n290), .A2(new_n223), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n375), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n218), .B1(new_n261), .B2(new_n265), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n264), .A2(G232), .A3(new_n260), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n225), .B2(new_n264), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n246), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n275), .B1(G244), .B2(new_n276), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(G179), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n384), .B1(new_n391), .B2(KEYINPUT71), .ZN(new_n392));
  AOI21_X1  g0192(.A(G169), .B1(new_n388), .B2(new_n389), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT71), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(new_n390), .B2(G179), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n383), .B1(new_n390), .B2(G200), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n388), .A2(G190), .A3(new_n389), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n320), .A2(new_n374), .A3(new_n400), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n223), .B2(new_n304), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n288), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g0204(.A(new_n404), .B(KEYINPUT11), .Z(new_n405));
  OR2_X1    g0205(.A1(new_n405), .A2(KEYINPUT75), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(KEYINPUT75), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n217), .B1(new_n292), .B2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(new_n290), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT12), .B1(new_n409), .B2(G68), .ZN(new_n410));
  OR3_X1    g0210(.A1(new_n409), .A2(KEYINPUT12), .A3(G68), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n291), .A2(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n406), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n264), .A2(KEYINPUT73), .A3(G226), .A4(new_n260), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n255), .A2(G226), .A3(new_n260), .A4(new_n258), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n255), .A2(G232), .A3(G1698), .A4(new_n258), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT74), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n417), .B2(new_n420), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT74), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n430), .A3(new_n246), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n275), .B1(G238), .B2(new_n276), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n416), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n246), .B1(new_n429), .B2(KEYINPUT74), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n427), .B(new_n424), .C1(new_n420), .C2(new_n417), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n416), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n415), .B(G169), .C1(new_n433), .C2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT13), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(G179), .A3(new_n436), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n436), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n415), .B1(new_n443), .B2(G169), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n414), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(G200), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n413), .C1(new_n447), .C2(new_n443), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n401), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n271), .A2(G1), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n246), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G257), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n451), .A2(new_n450), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n246), .A2(new_n274), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n255), .A2(G250), .A3(G1698), .A4(new_n258), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT4), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n224), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n255), .A2(new_n260), .A3(new_n258), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n260), .A2(G244), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n330), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n458), .A2(new_n461), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n457), .B1(new_n465), .B2(new_n246), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI211_X1 g0268(.A(KEYINPUT81), .B(new_n457), .C1(new_n246), .C2(new_n465), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n280), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n225), .A2(KEYINPUT6), .ZN(new_n471));
  INV_X1    g0271(.A(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT79), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G97), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g0276(.A(G97), .B(G107), .Z(new_n477));
  OAI22_X1  g0277(.A1(new_n476), .A2(KEYINPUT80), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n479));
  OAI21_X1  g0279(.A(G20), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n297), .A2(G77), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n350), .B1(new_n262), .B2(new_n263), .ZN(new_n482));
  INV_X1    g0282(.A(new_n349), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n288), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n409), .A2(G97), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n292), .A2(G33), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n287), .A2(new_n409), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(G97), .ZN(new_n491));
  INV_X1    g0291(.A(G179), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n486), .A2(new_n491), .B1(new_n466), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n470), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n224), .A2(G1698), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G238), .B2(G1698), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n330), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT82), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(new_n495), .C1(new_n330), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n246), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n321), .B(G250), .C1(G1), .C2(new_n271), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n455), .A2(new_n450), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n280), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n321), .B1(new_n499), .B2(new_n501), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n509), .A2(new_n492), .A3(new_n506), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT83), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(G169), .B1(new_n509), .B2(new_n506), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT83), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n503), .A2(new_n507), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n492), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT79), .B(G97), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n219), .A3(new_n225), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n211), .B1(new_n423), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n516), .B2(new_n304), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n330), .A2(G20), .A3(new_n217), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n288), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n377), .A2(new_n290), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n489), .A2(new_n377), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n511), .A2(new_n515), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n486), .A2(new_n491), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n466), .A2(new_n367), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n465), .A2(new_n246), .ZN(new_n534));
  INV_X1    g0334(.A(new_n457), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT81), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n466), .A2(new_n467), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(G190), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n490), .A2(G87), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n524), .A2(new_n541), .A3(new_n525), .ZN(new_n542));
  OAI21_X1  g0342(.A(G200), .B1(new_n509), .B2(new_n506), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n447), .C2(new_n514), .ZN(new_n544));
  AND4_X1   g0344(.A1(new_n494), .A2(new_n530), .A3(new_n540), .A4(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n287), .A2(G116), .A3(new_n409), .A4(new_n488), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n289), .A2(G1), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n211), .A2(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G116), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n282), .A2(new_n210), .B1(G20), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(G33), .B1(new_n473), .B2(new_n475), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n464), .A2(new_n211), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT20), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n553), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n516), .B2(G33), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT20), .B1(new_n557), .B2(new_n551), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n546), .B(new_n549), .C1(new_n555), .C2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(G303), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n255), .B2(new_n258), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n226), .A2(G1698), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G257), .B2(G1698), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n330), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n246), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n452), .A2(G270), .B1(new_n454), .B2(new_n455), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(new_n567), .A3(G169), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n567), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n559), .A3(G179), .ZN(new_n573));
  INV_X1    g0373(.A(new_n570), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n559), .A2(new_n567), .A3(G169), .A4(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(G303), .B1(new_n262), .B2(new_n263), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n327), .A2(new_n329), .A3(new_n256), .ZN(new_n577));
  INV_X1    g0377(.A(new_n563), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n321), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n451), .A2(new_n450), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n321), .A3(G270), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n456), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(G200), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n565), .A2(G190), .A3(new_n566), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n557), .A2(new_n551), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n554), .B1(new_n547), .B2(new_n548), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n584), .A2(new_n585), .A3(new_n589), .A4(new_n546), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n571), .A2(new_n573), .A3(new_n575), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n220), .A2(new_n260), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G257), .B2(new_n260), .ZN(new_n594));
  INV_X1    g0394(.A(G294), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n330), .A2(new_n594), .B1(new_n253), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n246), .B1(new_n452), .B2(G264), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n456), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n280), .ZN(new_n599));
  INV_X1    g0399(.A(new_n598), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n492), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n255), .A2(new_n211), .A3(G87), .A4(new_n258), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(KEYINPUT22), .A2(G87), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n495), .B1(new_n330), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n211), .ZN(new_n607));
  OAI211_X1 g0407(.A(KEYINPUT85), .B(KEYINPUT23), .C1(new_n211), .C2(G107), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n225), .A2(G20), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT85), .B1(new_n610), .B2(KEYINPUT23), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n609), .A2(new_n611), .B1(KEYINPUT23), .B2(new_n610), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n604), .A2(new_n607), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT24), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n602), .B2(new_n603), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT24), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n607), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n287), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n489), .A2(new_n225), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n290), .A2(new_n225), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT25), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n599), .B(new_n601), .C1(new_n619), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n614), .A2(KEYINPUT24), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n617), .B1(new_n616), .B2(new_n607), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n288), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n597), .A2(new_n447), .A3(new_n456), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n600), .B2(G200), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n631), .A3(new_n623), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n618), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n624), .B1(new_n634), .B2(new_n288), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT86), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n631), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n626), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n449), .A2(new_n545), .A3(new_n592), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n510), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n528), .B1(new_n640), .B2(new_n512), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT87), .B1(new_n542), .B2(new_n543), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n514), .A2(new_n447), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n542), .A2(KEYINPUT87), .A3(new_n543), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n633), .A2(new_n637), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n470), .A2(new_n493), .B1(new_n533), .B2(new_n539), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n573), .A2(new_n575), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n625), .A2(new_n571), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n646), .A2(new_n647), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n494), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n470), .A2(KEYINPUT88), .A3(new_n493), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n646), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n641), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n530), .A2(new_n544), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n658), .B2(new_n494), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n651), .A2(new_n656), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n449), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n373), .ZN(new_n662));
  INV_X1    g0462(.A(new_n396), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n448), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n445), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n363), .A2(new_n357), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n665), .A2(new_n667), .B1(new_n319), .B2(new_n318), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n668), .A2(KEYINPUT89), .A3(new_n308), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT89), .B1(new_n668), .B2(new_n308), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n661), .B1(new_n669), .B2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(KEYINPUT90), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n636), .B1(new_n635), .B2(new_n631), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n547), .A2(new_n211), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n635), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n625), .B1(new_n675), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n626), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n649), .A2(new_n571), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n682), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n672), .B1(new_n691), .B2(new_n685), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n672), .A3(new_n685), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n559), .A2(new_n681), .ZN(new_n696));
  MUX2_X1   g0496(.A(new_n688), .B(new_n592), .S(new_n696), .Z(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n687), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(G399));
  NOR2_X1   g0501(.A1(new_n517), .A2(G116), .ZN(new_n702));
  INV_X1    g0502(.A(new_n207), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n705), .A3(G1), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n215), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n646), .A2(new_n653), .A3(new_n655), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT26), .ZN(new_n711));
  INV_X1    g0511(.A(new_n494), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n654), .A3(new_n544), .A4(new_n530), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n711), .A2(new_n657), .A3(new_n651), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n709), .B1(new_n714), .B2(new_n682), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n591), .A2(new_n681), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n545), .A2(new_n717), .A3(new_n638), .A4(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n718), .B(new_n625), .C1(new_n673), .C2(new_n674), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n494), .A2(new_n530), .A3(new_n540), .A4(new_n544), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT91), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n597), .A2(new_n565), .A3(G179), .A4(new_n566), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n514), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n537), .A3(new_n538), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n725), .A2(KEYINPUT30), .A3(new_n537), .A4(new_n538), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n600), .A2(new_n572), .A3(G179), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n536), .A3(new_n514), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT31), .B1(new_n732), .B2(new_n681), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n716), .B1(new_n723), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n660), .A2(new_n709), .A3(new_n682), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n715), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n708), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n697), .A2(G330), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n289), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n292), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n704), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n698), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n210), .B1(G20), .B2(new_n280), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n577), .A2(new_n703), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G45), .B2(new_n215), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(G45), .B2(new_n244), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n264), .A2(new_n207), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n207), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n752), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(G317), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT33), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT33), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n211), .B1(new_n766), .B2(G190), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n765), .B1(new_n595), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n367), .A2(G179), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n211), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n766), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G283), .A2(new_n772), .B1(new_n774), .B2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n770), .A2(G179), .A3(new_n367), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n211), .A2(new_n447), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G179), .A3(new_n367), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n775), .B1(new_n776), .B2(new_n777), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n760), .A2(new_n447), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n768), .B(new_n781), .C1(G326), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n779), .A2(new_n769), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n259), .B1(new_n560), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT94), .Z(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(G159), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT32), .ZN(new_n788));
  INV_X1    g0588(.A(new_n761), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n789), .A2(new_n217), .B1(new_n767), .B2(new_n472), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n782), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n264), .B1(new_n792), .B2(new_n202), .ZN(new_n793));
  INV_X1    g0593(.A(new_n784), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G87), .A2(new_n794), .B1(new_n772), .B2(G107), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n300), .B2(new_n780), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n777), .A2(KEYINPUT93), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n777), .A2(KEYINPUT93), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n793), .B(new_n796), .C1(G77), .C2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n783), .A2(new_n786), .B1(new_n791), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n751), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n759), .B(new_n745), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT95), .Z(new_n805));
  INV_X1    g0605(.A(new_n750), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n697), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n747), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n660), .A2(new_n682), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n384), .A2(new_n682), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n392), .A2(new_n395), .A3(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n392), .A2(new_n395), .B1(new_n398), .B2(new_n397), .ZN(new_n813));
  INV_X1    g0613(.A(new_n811), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n812), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n400), .B2(new_n811), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n818), .A2(new_n660), .A3(new_n682), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n736), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n745), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  INV_X1    g0623(.A(new_n780), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G143), .B1(G137), .B2(new_n782), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  INV_X1    g0626(.A(new_n800), .ZN(new_n827));
  INV_X1    g0627(.A(G159), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n825), .B1(new_n826), .B2(new_n789), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n784), .A2(new_n202), .B1(new_n771), .B2(new_n217), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n577), .B1(new_n300), .B2(new_n767), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(G132), .C2(new_n774), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G107), .A2(new_n794), .B1(new_n774), .B2(G311), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n835), .B1(new_n219), .B2(new_n771), .C1(new_n827), .C2(new_n550), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n780), .A2(new_n595), .B1(new_n767), .B2(new_n472), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT96), .Z(new_n838));
  INV_X1    g0638(.A(G283), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n259), .B1(new_n792), .B2(new_n560), .C1(new_n839), .C2(new_n789), .ZN(new_n840));
  OR3_X1    g0640(.A1(new_n836), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n803), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n751), .A2(new_n748), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n746), .B(new_n842), .C1(new_n223), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n818), .B2(new_n749), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n823), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  NAND2_X1  g0647(.A1(new_n414), .A2(new_n681), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n445), .A2(new_n448), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(G169), .B1(new_n433), .B2(new_n437), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT14), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n441), .A3(new_n438), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n413), .B1(new_n443), .B2(new_n447), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n367), .B1(new_n440), .B2(new_n436), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n414), .B(new_n681), .C1(new_n852), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n371), .A2(new_n353), .A3(new_n355), .ZN(new_n859));
  INV_X1    g0659(.A(new_n679), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n356), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n361), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n347), .A2(new_n288), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT7), .B1(new_n577), .B2(G20), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(G68), .A3(new_n344), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT16), .B1(new_n866), .B2(new_n342), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n355), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n860), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT97), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT97), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n871), .A3(new_n860), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n337), .A2(new_n868), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n870), .A2(new_n859), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n863), .B1(new_n874), .B2(KEYINPUT37), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n364), .A2(new_n373), .B1(new_n872), .B2(new_n870), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n858), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n870), .A2(new_n872), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n374), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(KEYINPUT37), .B2(new_n862), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n815), .B1(new_n723), .B2(new_n735), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n857), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT99), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n863), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n861), .B1(new_n373), .B2(new_n666), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n858), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n886), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n857), .A3(new_n884), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n401), .A2(new_n445), .A3(new_n448), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n723), .B2(new_n735), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n896), .A2(new_n898), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n900), .A2(new_n716), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n669), .A2(new_n670), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n449), .B1(new_n715), .B2(new_n737), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT98), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT98), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n449), .B(new_n906), .C1(new_n715), .C2(new_n737), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n877), .A2(new_n882), .A3(KEYINPUT39), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n882), .A2(new_n893), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(KEYINPUT39), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n852), .A2(new_n414), .A3(new_n682), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n396), .A2(new_n681), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n819), .A2(new_n918), .B1(new_n849), .B2(new_n856), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n883), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n667), .A2(new_n679), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n909), .B(new_n922), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n902), .A2(new_n923), .B1(new_n292), .B2(new_n742), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n923), .B2(new_n902), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n478), .A2(new_n479), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n550), .B(new_n213), .C1(new_n927), .C2(KEYINPUT35), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(KEYINPUT35), .B2(new_n927), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT36), .Z(new_n930));
  OR3_X1    g0730(.A1(new_n215), .A2(new_n223), .A3(new_n338), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n202), .A2(G68), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n292), .B(G13), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n925), .A2(new_n930), .A3(new_n933), .ZN(G367));
  OR2_X1    g0734(.A1(new_n542), .A2(new_n682), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n646), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n657), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g0738(.A(new_n531), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n648), .B1(new_n939), .B2(new_n682), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n712), .A2(new_n681), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n687), .A2(new_n690), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n494), .B1(new_n940), .B2(new_n625), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT100), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT100), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n682), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n938), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n942), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n700), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n704), .B(KEYINPUT41), .Z(new_n957));
  INV_X1    g0757(.A(new_n700), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n693), .A2(new_n694), .A3(new_n954), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT45), .B1(new_n695), .B2(new_n942), .ZN(new_n963));
  INV_X1    g0763(.A(new_n694), .ZN(new_n964));
  OAI211_X1 g0764(.A(KEYINPUT45), .B(new_n942), .C1(new_n964), .C2(new_n692), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n958), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n695), .A2(new_n942), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n965), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n959), .B(new_n960), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n700), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n686), .B(new_n689), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n699), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n968), .A2(new_n974), .A3(new_n738), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n957), .B1(new_n977), .B2(new_n738), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n956), .B1(new_n978), .B2(new_n744), .ZN(new_n979));
  INV_X1    g0779(.A(new_n753), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n752), .B1(new_n207), .B2(new_n377), .C1(new_n980), .C2(new_n237), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n745), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT102), .Z(new_n983));
  OAI22_X1  g0783(.A1(new_n789), .A2(new_n828), .B1(new_n767), .B2(new_n217), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n259), .B(new_n984), .C1(G143), .C2(new_n782), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n771), .A2(new_n223), .ZN(new_n986));
  INV_X1    g0786(.A(G137), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n780), .A2(new_n826), .B1(new_n773), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(G58), .C2(new_n794), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n985), .B(new_n989), .C1(new_n202), .C2(new_n827), .ZN(new_n990));
  INV_X1    g0790(.A(new_n516), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n824), .A2(G303), .B1(new_n772), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n762), .B2(new_n773), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n794), .A2(G116), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT46), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n995), .A2(new_n996), .B1(new_n595), .B2(new_n789), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n792), .A2(new_n776), .B1(new_n767), .B2(new_n225), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n800), .A2(G283), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n577), .B1(new_n995), .B2(new_n996), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n994), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n990), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1004), .A2(KEYINPUT47), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n751), .B1(new_n1004), .B2(KEYINPUT47), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n983), .B1(new_n1005), .B2(new_n1006), .C1(new_n937), .C2(new_n806), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n979), .A2(new_n1007), .ZN(G387));
  OAI22_X1  g0808(.A1(new_n756), .A2(new_n702), .B1(G107), .B2(new_n207), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n702), .B(new_n271), .C1(new_n217), .C2(new_n223), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT103), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT103), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n379), .A2(G50), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n980), .B1(new_n234), .B2(G45), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n752), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n745), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n771), .A2(new_n472), .B1(new_n773), .B2(new_n826), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G50), .B2(new_n824), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n303), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n761), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n217), .A2(new_n777), .B1(new_n784), .B2(new_n223), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n330), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n767), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n377), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1027), .A2(new_n1028), .B1(G159), .B2(new_n782), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n800), .A2(G303), .B1(G317), .B2(new_n824), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n789), .A2(new_n776), .B1(new_n792), .B2(new_n778), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT104), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT104), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n784), .A2(new_n595), .B1(new_n767), .B2(new_n839), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(G326), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n330), .B1(new_n773), .B2(new_n1041), .C1(new_n550), .C2(new_n771), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT105), .Z(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT49), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1030), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT106), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n803), .B1(new_n1046), .B2(KEYINPUT106), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1020), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n687), .B2(new_n806), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT107), .Z(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n744), .B2(new_n976), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n976), .A2(new_n738), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n976), .A2(new_n738), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n704), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1052), .B1(new_n1053), .B2(new_n1055), .ZN(G393));
  NAND2_X1  g0856(.A1(new_n968), .A2(new_n974), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1054), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n704), .A3(new_n977), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n968), .A2(new_n974), .A3(new_n744), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n752), .B1(new_n207), .B2(new_n516), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n241), .B2(new_n753), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n577), .B1(new_n223), .B2(new_n767), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G50), .B2(new_n761), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n784), .A2(new_n217), .B1(new_n771), .B2(new_n219), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G143), .B2(new_n774), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(new_n827), .C2(new_n379), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n824), .A2(G159), .B1(G150), .B2(new_n782), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n264), .B1(G303), .B2(new_n761), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n784), .A2(new_n839), .B1(new_n771), .B2(new_n225), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n777), .A2(new_n595), .B1(new_n773), .B2(new_n778), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1070), .B(new_n1073), .C1(new_n550), .C2(new_n767), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n762), .A2(new_n792), .B1(new_n780), .B2(new_n776), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT108), .B(KEYINPUT52), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1067), .A2(new_n1069), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n746), .B(new_n1062), .C1(new_n1078), .C2(new_n751), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n942), .B2(new_n806), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1060), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1059), .A2(new_n1081), .ZN(G390));
  NOR3_X1   g0882(.A1(new_n821), .A2(new_n897), .A3(KEYINPUT110), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT110), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n449), .B2(new_n736), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n903), .A2(new_n908), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n736), .A2(new_n818), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n857), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT111), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n857), .A2(new_n736), .A3(new_n818), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n819), .A2(new_n918), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1088), .A2(new_n1089), .A3(KEYINPUT111), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n494), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(KEYINPUT26), .B2(new_n710), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n651), .A2(new_n657), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n681), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n917), .B1(new_n1100), .B2(new_n818), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT109), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n857), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n849), .A2(new_n856), .A3(KEYINPUT109), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1088), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1092), .B(new_n1101), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1096), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n912), .B1(new_n915), .B2(new_n919), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1101), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n911), .A2(new_n915), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1092), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1109), .B(new_n1092), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1087), .A2(new_n1108), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1116), .A2(new_n704), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1087), .A2(new_n1108), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(KEYINPUT112), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT112), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1117), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1114), .A2(new_n744), .A3(new_n1115), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n843), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n784), .A2(new_n826), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n264), .B1(new_n1128), .B2(KEYINPUT53), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n824), .A2(G132), .B1(new_n774), .B2(G125), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n202), .B2(new_n771), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1129), .B(new_n1131), .C1(new_n800), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n792), .A2(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n789), .A2(new_n987), .B1(new_n767), .B2(new_n828), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(KEYINPUT53), .C2(new_n1128), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n789), .A2(new_n225), .B1(new_n792), .B2(new_n839), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n264), .B(new_n1139), .C1(G77), .C2(new_n1027), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n784), .A2(new_n219), .B1(new_n771), .B2(new_n217), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n780), .A2(new_n550), .B1(new_n773), .B2(new_n595), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n800), .C2(new_n991), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1134), .A2(new_n1138), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n745), .B1(new_n1023), .B2(new_n1126), .C1(new_n1144), .C2(new_n803), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT113), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n913), .B2(new_n749), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1125), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1124), .A2(new_n1149), .ZN(G378));
  AND2_X1   g0950(.A1(new_n895), .A2(G330), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n887), .B2(new_n888), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT115), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g0954(.A(KEYINPUT115), .B(new_n1151), .C1(new_n887), .C2(new_n888), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n307), .A2(new_n860), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n320), .B(new_n1156), .Z(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1154), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n922), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n889), .A2(KEYINPUT115), .A3(new_n1151), .A4(new_n1159), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1116), .A2(new_n1087), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT57), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n922), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1116), .B2(new_n1087), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n704), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1159), .A2(new_n748), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n745), .B1(new_n1126), .B2(G50), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n577), .A2(G41), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G50), .B(new_n1179), .C1(new_n253), .C2(new_n270), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n780), .A2(new_n225), .B1(new_n784), .B2(new_n223), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G68), .B2(new_n1027), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n777), .A2(new_n377), .B1(new_n773), .B2(new_n839), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G58), .B2(new_n772), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G97), .A2(new_n761), .B1(new_n782), .B2(G116), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .A4(new_n1179), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT58), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G132), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n789), .A2(new_n1189), .B1(new_n777), .B2(new_n987), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT114), .Z(new_n1191));
  AND2_X1   g0991(.A1(new_n782), .A2(G125), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n767), .A2(new_n826), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n780), .A2(new_n1135), .B1(new_n784), .B2(new_n1132), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n253), .B(new_n270), .C1(new_n771), .C2(new_n828), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G124), .B2(new_n774), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT59), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1199), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1188), .B1(new_n1187), .B2(new_n1186), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1178), .B1(new_n1202), .B2(new_n751), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1177), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1166), .B2(new_n744), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1176), .A2(new_n1206), .ZN(G375));
  AOI21_X1  g1007(.A(new_n746), .B1(new_n217), .B2(new_n843), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n800), .A2(G107), .B1(G116), .B2(new_n761), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT116), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n824), .A2(G283), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT117), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT117), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1210), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n259), .B1(new_n792), .B2(new_n595), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n986), .B1(G303), .B2(new_n774), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n472), .B2(new_n784), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(new_n1209), .C2(KEYINPUT116), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n777), .A2(new_n826), .B1(new_n767), .B2(new_n202), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT118), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n784), .A2(new_n828), .B1(new_n773), .B2(new_n1135), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT119), .Z(new_n1223));
  OAI22_X1  g1023(.A1(new_n1189), .A2(new_n792), .B1(new_n789), .B2(new_n1132), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n780), .A2(new_n987), .B1(new_n771), .B2(new_n300), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1223), .A2(new_n330), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1215), .A2(new_n1219), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1208), .B1(new_n803), .B2(new_n1227), .C1(new_n1105), .C2(new_n749), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1108), .B2(new_n744), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n957), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1118), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1087), .A2(new_n1108), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1230), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  INV_X1    g1034(.A(G375), .ZN(new_n1235));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT120), .Z(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1239), .A2(G387), .A3(G381), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1124), .A2(new_n1149), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1235), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT121), .ZN(G407));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1206), .C1(new_n1168), .C2(new_n1175), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1170), .A2(new_n1231), .A3(new_n1173), .A4(new_n1167), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1170), .A2(new_n744), .A3(new_n1173), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1204), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1241), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1245), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n903), .A2(new_n908), .A3(new_n1086), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1257), .A2(KEYINPUT60), .A3(new_n1096), .A4(new_n1107), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n704), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1087), .B2(new_n1108), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n1233), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1230), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n846), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G384), .B(new_n1230), .C1(new_n1259), .C2(new_n1262), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1255), .A2(new_n1256), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1246), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1268), .A2(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  XOR2_X1   g1072(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AND4_X1   g1074(.A1(G2897), .A2(new_n1264), .A3(new_n1245), .A4(new_n1265), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1264), .A2(new_n1265), .B1(G2897), .B2(new_n1246), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1249), .B1(new_n1272), .B2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(new_n808), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(new_n1236), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n979), .A2(G390), .A3(new_n1007), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(G387), .A2(KEYINPUT123), .A3(new_n1236), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n979), .A2(G390), .A3(KEYINPUT124), .A4(new_n1007), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1285), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT123), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1280), .B1(new_n1282), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1284), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n1245), .B(new_n1266), .C1(new_n1250), .C2(new_n1254), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(KEYINPUT62), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1246), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1255), .A2(new_n1296), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1273), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1295), .A2(KEYINPUT126), .A3(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1279), .A2(new_n1292), .A3(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1291), .A2(new_n1288), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1284), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT61), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1294), .A2(KEYINPUT63), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1270), .A2(KEYINPUT63), .A3(new_n1267), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1298), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .A4(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1301), .A2(new_n1309), .ZN(G405));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1241), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1250), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(KEYINPUT127), .A3(new_n1267), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1267), .A2(KEYINPUT127), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1311), .A2(new_n1250), .A3(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1313), .A2(new_n1292), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1292), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


