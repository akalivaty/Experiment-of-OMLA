//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT64), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n474), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT65), .B1(new_n462), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n493), .A2(KEYINPUT66), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n474), .A2(G138), .A3(new_n494), .A4(new_n462), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n496));
  INV_X1    g071(.A(new_n494), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n495), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(new_n504), .A2(new_n507), .A3(G89), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(KEYINPUT67), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(new_n510), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G168));
  XOR2_X1   g104(.A(KEYINPUT69), .B(G90), .Z(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT68), .B(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n508), .A2(new_n530), .B1(new_n510), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n514), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n532), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  XOR2_X1   g111(.A(KEYINPUT70), .B(G81), .Z(new_n537));
  NOR2_X1   g112(.A1(new_n508), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n514), .ZN(new_n540));
  AOI211_X1 g115(.A(new_n538), .B(new_n540), .C1(G43), .C2(new_n526), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT72), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n501), .A2(new_n503), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n555), .B2(new_n508), .ZN(new_n556));
  OAI211_X1 g131(.A(G53), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n559), .A2(KEYINPUT74), .A3(new_n561), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n556), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n528), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n528), .A2(new_n568), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND3_X1  g149(.A1(new_n504), .A2(new_n507), .A3(G87), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT76), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n526), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  AOI22_X1  g154(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n514), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n504), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(new_n507), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n508), .A2(new_n587), .B1(new_n510), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n514), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n504), .A2(new_n507), .A3(G92), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT10), .Z(new_n596));
  NAND2_X1  g171(.A1(new_n526), .A2(G54), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n514), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n594), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n572), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n566), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT77), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(KEYINPUT77), .B2(new_n604), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(KEYINPUT77), .B2(new_n604), .ZN(G280));
  XNOR2_X1  g183(.A(KEYINPUT78), .B(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n600), .B1(G860), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT79), .Z(G148));
  NAND2_X1  g186(.A1(new_n600), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n476), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n478), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT80), .Z(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n635), .B(new_n637), .Z(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n638), .A2(new_n639), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n647), .B(KEYINPUT84), .Z(new_n651));
  OAI21_X1  g226(.A(KEYINPUT17), .B1(new_n651), .B2(new_n646), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n646), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n664), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n662), .B2(new_n663), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n661), .A2(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1986), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n674), .B(new_n678), .ZN(G229));
  NOR2_X1   g254(.A1(G29), .A2(G32), .ZN(new_n680));
  AOI22_X1  g255(.A1(new_n476), .A2(G141), .B1(new_n478), .B2(G129), .ZN(new_n681));
  NAND3_X1  g256(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT26), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT97), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n680), .B1(new_n689), .B2(G29), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT27), .B(G1996), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(G160), .A2(G29), .ZN(new_n693));
  NOR2_X1   g268(.A1(KEYINPUT24), .A2(G34), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(KEYINPUT24), .A2(G34), .ZN(new_n696));
  AOI21_X1  g271(.A(G29), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n693), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G2084), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G5), .A2(G16), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G171), .B2(G16), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n692), .B(new_n702), .C1(G1961), .C2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT99), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT31), .B(G11), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n690), .A2(new_n691), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NOR2_X1   g284(.A1(G164), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G27), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G2078), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n709), .A2(G33), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G139), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n475), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI22_X1  g297(.A1(new_n720), .A2(new_n721), .B1(new_n462), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n714), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2072), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI22_X1  g301(.A1(new_n724), .A2(new_n725), .B1(new_n712), .B2(new_n711), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n708), .A2(new_n713), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n709), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n709), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2090), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1966), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n621), .A2(new_n709), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n704), .A2(G1961), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n700), .A2(new_n701), .ZN(new_n739));
  INV_X1    g314(.A(G28), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n741), .A2(new_n742), .A3(new_n709), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n732), .A2(new_n736), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n706), .A2(new_n707), .A3(new_n728), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n733), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n541), .B2(new_n733), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1341), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT91), .B1(G4), .B2(G16), .ZN(new_n751));
  OR3_X1    g326(.A1(KEYINPUT91), .A2(G4), .A3(G16), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n733), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1348), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n709), .A2(G26), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n476), .A2(G140), .B1(new_n478), .B2(G128), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n462), .A2(G116), .ZN(new_n758));
  OR3_X1    g333(.A1(KEYINPUT93), .A2(G104), .A3(G2105), .ZN(new_n759));
  OAI21_X1  g334(.A(KEYINPUT93), .B1(G104), .B2(G2105), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n759), .A2(G2104), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n757), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(G29), .ZN(new_n763));
  MUX2_X1   g338(.A(new_n756), .B(new_n763), .S(KEYINPUT28), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2067), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n750), .A2(new_n755), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n733), .A2(G20), .ZN(new_n769));
  OAI211_X1 g344(.A(KEYINPUT23), .B(new_n769), .C1(new_n566), .C2(new_n733), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT23), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n746), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n766), .A2(new_n767), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G16), .B2(G23), .ZN(new_n777));
  OR3_X1    g352(.A1(new_n776), .A2(G16), .A3(G23), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n777), .B(new_n778), .C1(G288), .C2(new_n733), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT33), .B(G1976), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n733), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n733), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1971), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n733), .A2(G6), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n585), .B2(new_n733), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT32), .B(G1981), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n781), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT89), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n733), .A2(G24), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n592), .B2(new_n733), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1986), .Z(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(KEYINPUT90), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n790), .B2(KEYINPUT34), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(KEYINPUT90), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n709), .A2(G25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n476), .A2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n478), .A2(G119), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n709), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT35), .B(G1991), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n791), .A2(new_n797), .A3(new_n798), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n791), .A2(new_n809), .A3(new_n797), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n811), .A2(KEYINPUT90), .A3(new_n795), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n774), .A2(new_n775), .A3(new_n810), .A4(new_n812), .ZN(G150));
  INV_X1    g388(.A(G150), .ZN(G311));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n508), .A2(new_n815), .B1(new_n510), .B2(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n514), .ZN(new_n819));
  OAI21_X1  g394(.A(G860), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n600), .A2(G559), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT39), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n817), .A2(new_n819), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n541), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n821), .B1(new_n828), .B2(G860), .ZN(G145));
  NAND2_X1  g404(.A1(new_n478), .A2(G130), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n476), .A2(G142), .ZN(new_n832));
  NOR2_X1   g407(.A1(G106), .A2(G2105), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n689), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n723), .B(new_n624), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n492), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n490), .A2(KEYINPUT101), .A3(new_n491), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n498), .A2(new_n495), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n837), .A2(new_n843), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n836), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n687), .A2(new_n688), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n835), .ZN(new_n849));
  INV_X1    g424(.A(new_n844), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n845), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n762), .B(new_n804), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n847), .A2(new_n851), .A3(new_n853), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n621), .B(G160), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n482), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(G37), .B1(new_n859), .B2(KEYINPUT103), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(new_n856), .ZN(new_n861));
  INV_X1    g436(.A(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n855), .A2(new_n856), .A3(new_n864), .A4(new_n858), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n826), .A2(G868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n612), .B(KEYINPUT104), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n827), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n600), .A2(new_n566), .ZN(new_n873));
  NAND2_X1  g448(.A1(G299), .A2(new_n753), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n827), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n871), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n875), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G166), .B(new_n592), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G305), .ZN(new_n884));
  INV_X1    g459(.A(G288), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT42), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n887), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n868), .B(new_n870), .C1(new_n890), .C2(new_n603), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n603), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT105), .B1(new_n892), .B2(new_n869), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(G295));
  OAI21_X1  g469(.A(new_n870), .B1(new_n890), .B2(new_n603), .ZN(G331));
  OAI21_X1  g470(.A(G171), .B1(new_n570), .B2(new_n571), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n528), .A2(G171), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n877), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(G168), .A2(KEYINPUT75), .ZN(new_n900));
  AOI21_X1  g475(.A(G301), .B1(new_n900), .B2(new_n569), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n827), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n875), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n880), .A2(new_n902), .A3(new_n899), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n886), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT107), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n904), .A2(new_n886), .A3(new_n905), .A4(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(new_n886), .ZN(new_n913));
  INV_X1    g488(.A(new_n904), .ZN(new_n914));
  INV_X1    g489(.A(new_n905), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n911), .A2(KEYINPUT108), .A3(new_n912), .A4(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n914), .A2(new_n915), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n908), .C1(new_n918), .C2(new_n906), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n906), .B2(KEYINPUT107), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(new_n912), .A3(new_n916), .A4(new_n910), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n911), .A2(KEYINPUT43), .A3(new_n916), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n920), .A2(new_n912), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(G397));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n842), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n467), .A2(new_n468), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G2105), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n470), .A2(new_n471), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n462), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n940), .A3(G40), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n936), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n848), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n762), .B(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n808), .B2(new_n805), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n804), .A2(new_n807), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n956));
  INV_X1    g531(.A(new_n946), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n957), .A2(G1986), .A3(G290), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT48), .Z(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n689), .B2(new_n950), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n946), .A2(new_n947), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(KEYINPUT125), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n963), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(KEYINPUT125), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n762), .A2(G2067), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n951), .B2(new_n953), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n960), .B(new_n969), .C1(new_n957), .C2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n945), .A2(new_n934), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n978));
  NOR2_X1   g553(.A1(G305), .A2(G1981), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n585), .A2(new_n676), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT49), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n978), .B(new_n983), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n976), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n885), .ZN(new_n987));
  INV_X1    g562(.A(new_n979), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n842), .A2(new_n990), .A3(new_n933), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n991), .A2(new_n992), .A3(new_n943), .A4(new_n944), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(G2090), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n995));
  INV_X1    g570(.A(G40), .ZN(new_n996));
  NOR4_X1   g571(.A1(new_n469), .A2(new_n472), .A3(new_n942), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n490), .A2(new_n491), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n841), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT110), .B(new_n935), .C1(G164), .C2(G1384), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1971), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT55), .Z(new_n1011));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n994), .A2(new_n1007), .A3(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1009), .A2(G8), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G288), .A2(new_n986), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT52), .B1(new_n977), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(G288), .B2(new_n986), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n976), .B(new_n1018), .C1(new_n986), .C2(G288), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n985), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n989), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1020), .A2(KEYINPUT63), .A3(new_n1014), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1009), .A2(G8), .A3(new_n1013), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1011), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1966), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n841), .A2(new_n1000), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(new_n943), .A3(new_n944), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT45), .B1(new_n842), .B2(new_n933), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n998), .A2(new_n701), .A3(new_n992), .A4(new_n991), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n572), .A2(G8), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1026), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT113), .B(KEYINPUT63), .Z(new_n1037));
  OAI21_X1  g612(.A(new_n1021), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1034), .A2(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n528), .A2(G8), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT51), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1044), .B(G8), .C1(new_n1034), .C2(new_n528), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT120), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1040), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1047), .B(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(KEYINPUT121), .A3(new_n1045), .A4(new_n1043), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1049), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1050), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1005), .B2(G2078), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT123), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(new_n1057), .C1(new_n1005), .C2(G2078), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n936), .A2(new_n998), .A3(new_n712), .A4(new_n1029), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1057), .B1(new_n1063), .B2(KEYINPUT122), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n712), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1064), .A2(new_n1067), .B1(new_n1068), .B2(new_n993), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1039), .B1(new_n1056), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n993), .A2(new_n1068), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1031), .A2(G2078), .A3(new_n941), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1004), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1004), .A2(new_n1003), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(new_n712), .A3(new_n998), .A4(new_n1002), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1060), .B1(new_n1079), .B2(new_n1057), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1061), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1075), .B(new_n1077), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1071), .B(new_n1074), .C1(G171), .C2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1062), .A2(new_n1069), .A3(G301), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(G171), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1062), .A2(new_n1069), .A3(KEYINPUT124), .A4(G301), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1083), .B1(new_n1089), .B2(new_n1074), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT56), .B(G2072), .Z(new_n1091));
  NOR2_X1   g666(.A1(new_n1005), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n556), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n559), .B2(new_n561), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n566), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n990), .B1(new_n842), .B2(new_n933), .ZN(new_n1100));
  NOR3_X1   g675(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n945), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1102), .A2(KEYINPUT114), .A3(G1956), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1001), .A2(new_n990), .ZN(new_n1105));
  INV_X1    g680(.A(new_n934), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n998), .B(new_n1105), .C1(new_n1106), .C2(new_n990), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1104), .B1(new_n1107), .B2(new_n772), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1093), .B(new_n1099), .C1(new_n1103), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1098), .B(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT114), .B1(new_n1102), .B2(G1956), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1104), .A3(new_n772), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1114), .B2(new_n1093), .ZN(new_n1115));
  INV_X1    g690(.A(G1348), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n993), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n998), .A2(new_n1106), .A3(new_n949), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n753), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1109), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1078), .A2(new_n947), .A3(new_n998), .A4(new_n1002), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n945), .B2(new_n934), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1122), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1122), .B(new_n1125), .C1(new_n1005), .C2(G1996), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n541), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  OAI221_X1 g708(.A(new_n541), .B1(new_n1130), .B2(new_n1131), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(KEYINPUT119), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1136), .A2(KEYINPUT119), .A3(new_n753), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n753), .B1(new_n1136), .B2(KEYINPUT119), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1099), .B1(new_n1114), .B2(new_n1093), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1098), .B(new_n1092), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1135), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1109), .A2(KEYINPUT61), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT118), .B1(new_n1148), .B2(new_n1115), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1093), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1111), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1152), .A2(new_n1153), .A3(KEYINPUT61), .A4(new_n1109), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1121), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1090), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1073), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(G2090), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1160), .A2(new_n1102), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1024), .B1(new_n1161), .B2(new_n975), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1020), .A2(new_n1014), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1038), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n952), .A2(new_n953), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n592), .B(G1986), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n957), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n973), .B1(new_n1164), .B2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g743(.A(G227), .B1(new_n642), .B2(new_n643), .ZN(new_n1170));
  AND2_X1   g744(.A1(new_n866), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g745(.A1(G229), .A2(new_n460), .ZN(new_n1172));
  AND3_X1   g746(.A1(new_n1171), .A2(new_n926), .A3(new_n1172), .ZN(G308));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n926), .A3(new_n1172), .ZN(G225));
endmodule


