//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n187), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n201), .B(new_n203), .C1(G119), .C2(new_n202), .ZN(new_n204));
  XNOR2_X1  g018(.A(G119), .B(G128), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT24), .B(G110), .Z(new_n206));
  AOI22_X1  g020(.A1(new_n204), .A2(G110), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n198), .A2(new_n207), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n204), .A2(G110), .B1(new_n205), .B2(new_n206), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n209), .B(new_n197), .C1(G146), .C2(new_n193), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G137), .ZN(new_n212));
  INV_X1    g026(.A(G221), .ZN(new_n213));
  INV_X1    g027(.A(G234), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n213), .A2(new_n214), .A3(G953), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n212), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n208), .A2(new_n210), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(G217), .B1(new_n214), .B2(G902), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(KEYINPUT76), .ZN(new_n222));
  INV_X1    g036(.A(G902), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n224), .B(KEYINPUT78), .Z(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n223), .A3(new_n219), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n227), .A2(KEYINPUT25), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n222), .B(KEYINPUT77), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n227), .B2(KEYINPUT25), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(KEYINPUT79), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n234));
  NOR2_X1   g048(.A1(G237), .A2(G953), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G210), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n234), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G101), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n200), .A2(G116), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g058(.A(G116), .B(G119), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT2), .B(G113), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n245), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G128), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT64), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n195), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n255), .A2(new_n257), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(G137), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  INV_X1    g089(.A(G131), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(new_n272), .A3(new_n276), .A4(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n252), .B1(new_n267), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT1), .B1(new_n259), .B2(G146), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n259), .A2(G146), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n195), .A2(G143), .ZN(new_n282));
  OAI211_X1 g096(.A(G128), .B(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n269), .A2(G137), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n271), .A2(G134), .ZN(new_n285));
  OAI21_X1  g099(.A(G131), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n258), .B(new_n260), .C1(KEYINPUT1), .C2(new_n202), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n283), .A2(new_n277), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT28), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n288), .B(KEYINPUT68), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n279), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n271), .A2(G134), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n276), .B1(new_n295), .B2(new_n273), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT11), .B1(new_n271), .B2(G134), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n285), .A2(G131), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(KEYINPUT68), .A3(new_n287), .A4(new_n283), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n288), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n299), .A2(new_n300), .B1(new_n274), .B2(G131), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n249), .B(new_n251), .C1(new_n266), .C2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT69), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n294), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT65), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n266), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n255), .A2(new_n265), .A3(KEYINPUT65), .A4(new_n257), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n278), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n283), .A2(new_n287), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n301), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n252), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n309), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n291), .B1(new_n321), .B2(KEYINPUT28), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n294), .A2(new_n308), .B1(new_n319), .B2(new_n252), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n323), .A2(new_n290), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n239), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n267), .A2(new_n278), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(KEYINPUT30), .A3(new_n304), .A4(new_n302), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n306), .B1(new_n266), .B2(new_n310), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n329), .A2(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n252), .C1(new_n330), .C2(KEYINPUT30), .ZN(new_n331));
  INV_X1    g145(.A(new_n239), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n309), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT31), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(KEYINPUT31), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n326), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G472), .A2(G902), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n233), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n321), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n340));
  INV_X1    g154(.A(new_n289), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n323), .B2(new_n324), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n332), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n336), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n344), .A2(new_n334), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n338), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT32), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT75), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n337), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n339), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n239), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n327), .A2(new_n304), .A3(new_n302), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n294), .A2(new_n308), .B1(new_n252), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n341), .B(new_n356), .C1(new_n358), .C2(new_n324), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n359), .A2(KEYINPUT74), .A3(new_n223), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT74), .B1(new_n359), .B2(new_n223), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n331), .A2(new_n309), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n239), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n340), .A2(new_n343), .A3(new_n332), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n355), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n366), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G472), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n232), .B1(new_n354), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G107), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT80), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n374), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(G107), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n377), .A2(KEYINPUT80), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G104), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n380), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n376), .A2(new_n378), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n383), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n382), .A2(G104), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n374), .B2(new_n376), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(KEYINPUT4), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n387), .B2(new_n389), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(new_n252), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n240), .A2(new_n242), .A3(new_n246), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n246), .B1(new_n240), .B2(new_n242), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT5), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G113), .ZN(new_n400));
  INV_X1    g214(.A(new_n240), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n399), .A2(new_n403), .B1(new_n250), .B2(new_n245), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n390), .B1(new_n383), .B2(new_n380), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n379), .A2(new_n384), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n390), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G122), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n372), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n394), .A2(new_n393), .B1(new_n249), .B2(new_n251), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n413), .A2(new_n392), .B1(new_n404), .B2(new_n407), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT86), .B1(new_n414), .B2(new_n410), .ZN(new_n415));
  AND4_X1   g229(.A1(KEYINPUT86), .A2(new_n396), .A3(new_n408), .A4(new_n410), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n372), .A3(new_n411), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n266), .A2(G125), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n283), .A2(new_n287), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n191), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G953), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G224), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n422), .B(new_n424), .Z(new_n425));
  NAND3_X1  g239(.A1(new_n417), .A2(new_n418), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n409), .B2(new_n411), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n414), .A2(KEYINPUT86), .A3(new_n410), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n403), .A2(new_n431), .B1(new_n250), .B2(new_n245), .ZN(new_n432));
  INV_X1    g246(.A(new_n405), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n391), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT87), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n407), .A2(new_n436), .A3(new_n432), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n435), .B(new_n437), .C1(new_n407), .C2(new_n404), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n410), .B(KEYINPUT8), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n422), .A2(KEYINPUT7), .A3(new_n424), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n419), .A2(new_n421), .A3(new_n441), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n438), .A2(new_n439), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n430), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n426), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G210), .B1(G237), .B2(G902), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(KEYINPUT88), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n426), .A2(new_n444), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT85), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT94), .B1(new_n259), .B2(G128), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT94), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n202), .A3(G143), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n259), .A2(G128), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n259), .A2(KEYINPUT13), .A3(G128), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G134), .ZN(new_n464));
  INV_X1    g278(.A(G122), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT93), .B1(new_n465), .B2(G116), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n241), .A3(G122), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n241), .A2(G122), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n382), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n382), .B1(new_n469), .B2(new_n471), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n464), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n456), .B1(new_n202), .B2(G143), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n259), .A2(KEYINPUT94), .A3(G128), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n459), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT95), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n458), .A2(new_n480), .A3(new_n459), .ZN(new_n481));
  AOI21_X1  g295(.A(G134), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n469), .A2(KEYINPUT14), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n466), .A2(new_n468), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n471), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n487), .A2(new_n488), .A3(G107), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n487), .B2(G107), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n458), .A2(new_n480), .A3(new_n459), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n480), .B1(new_n458), .B2(new_n459), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n269), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n479), .A2(G134), .A3(new_n481), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n473), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n483), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT9), .B(G234), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(G217), .A3(new_n423), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT98), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n494), .A2(new_n495), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n466), .A2(new_n468), .A3(new_n485), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n485), .B1(new_n466), .B2(new_n468), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n504), .A2(new_n505), .A3(new_n470), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT96), .B1(new_n506), .B2(new_n382), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n487), .A2(new_n488), .A3(G107), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n503), .A2(new_n507), .A3(new_n472), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n483), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT98), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n497), .B2(new_n501), .ZN(new_n515));
  AND4_X1   g329(.A1(new_n514), .A2(new_n509), .A3(new_n510), .A4(new_n501), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n502), .B(new_n513), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n223), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n517), .B2(new_n223), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n525));
  NOR2_X1   g339(.A1(G475), .A2(G902), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n526), .B(KEYINPUT90), .Z(new_n527));
  AND3_X1   g341(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT19), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT19), .B1(new_n190), .B2(new_n192), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n195), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n235), .A2(G143), .A3(G214), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(G143), .B1(new_n235), .B2(G214), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n532), .A2(new_n533), .A3(G131), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n235), .A2(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n259), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n276), .B1(new_n536), .B2(new_n531), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n530), .B(new_n197), .C1(new_n534), .C2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n193), .B(G146), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT18), .B(G131), .C1(new_n532), .C2(new_n533), .ZN(new_n540));
  NAND2_X1  g354(.A1(KEYINPUT18), .A2(G131), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n536), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n545));
  XNOR2_X1  g359(.A(G113), .B(G122), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(new_n373), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n538), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT17), .ZN(new_n552));
  OAI211_X1 g366(.A(KEYINPUT17), .B(G131), .C1(new_n532), .C2(new_n533), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n196), .A2(new_n553), .A3(new_n197), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n547), .B(new_n543), .C1(new_n552), .C2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n527), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n525), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n555), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n550), .A2(new_n548), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n560), .B2(new_n545), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n561), .C2(new_n527), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n551), .A2(new_n555), .ZN(new_n563));
  INV_X1    g377(.A(new_n527), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n543), .B1(new_n552), .B2(new_n554), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n548), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n568), .B2(new_n555), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT92), .B(G475), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n423), .A2(G952), .ZN(new_n574));
  NAND2_X1  g388(.A1(G234), .A2(G237), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT99), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT21), .B(G898), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(G902), .A3(G953), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n524), .A2(new_n573), .A3(KEYINPUT100), .A4(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n517), .A2(new_n223), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n519), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n521), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n566), .A2(new_n571), .A3(new_n583), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n213), .B1(new_n499), .B2(new_n223), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G140), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n423), .A2(G227), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n392), .A2(new_n267), .A3(new_n395), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n407), .B2(new_n314), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n379), .A2(new_n384), .A3(G101), .ZN(new_n600));
  NOR4_X1   g414(.A1(new_n600), .A2(new_n420), .A3(KEYINPUT10), .A4(new_n405), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n306), .B(new_n597), .C1(new_n599), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT81), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n407), .A2(new_n598), .A3(new_n314), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n391), .A2(new_n433), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT10), .B1(new_n605), .B2(new_n420), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT81), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n306), .A4(new_n597), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT82), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n278), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n407), .A2(new_n314), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n420), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n610), .A2(new_n616), .A3(KEYINPUT83), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n596), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n595), .B1(new_n603), .B2(new_n609), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n266), .B1(new_n394), .B2(new_n393), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n606), .A2(new_n604), .B1(new_n623), .B2(new_n392), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n306), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n223), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G469), .ZN(new_n630));
  INV_X1    g444(.A(G469), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n610), .A2(new_n616), .A3(new_n596), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n596), .B1(new_n610), .B2(new_n626), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n631), .B(new_n223), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT84), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n616), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n625), .B1(new_n609), .B2(new_n603), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(new_n596), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n639), .A2(KEYINPUT84), .A3(new_n631), .A4(new_n223), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n592), .B1(new_n630), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n371), .A2(new_n454), .A3(new_n591), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G101), .ZN(G3));
  INV_X1    g458(.A(G472), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n337), .B2(new_n223), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n344), .A2(new_n345), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n347), .B1(new_n647), .B2(new_n335), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n646), .A2(new_n648), .A3(new_n232), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT101), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n586), .A2(new_n518), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n517), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n509), .A2(new_n510), .A3(new_n501), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(new_n511), .A3(new_n653), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n518), .A2(G902), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n652), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n572), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n426), .A2(new_n447), .A3(new_n444), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n447), .B1(new_n426), .B2(new_n444), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n453), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n583), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n651), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n565), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n556), .A2(KEYINPUT102), .A3(new_n557), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n673), .A2(new_n558), .A3(new_n562), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n571), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n667), .A2(new_n524), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n651), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT35), .B(G107), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  NOR2_X1   g494(.A1(new_n216), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n211), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n225), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n228), .B2(new_n230), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n449), .A2(new_n666), .A3(new_n450), .A4(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n646), .A2(new_n648), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n642), .A2(new_n591), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  AOI22_X1  g503(.A1(new_n629), .A2(G469), .B1(new_n636), .B2(new_n640), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n578), .B1(new_n691), .B2(new_n581), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n588), .A2(new_n571), .A3(new_n675), .A4(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n690), .A2(new_n592), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n351), .A2(new_n353), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n337), .A2(new_n338), .ZN(new_n697));
  INV_X1    g511(.A(new_n233), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n370), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n685), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n695), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT103), .B(G128), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G30));
  XOR2_X1   g518(.A(new_n692), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n642), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  INV_X1    g521(.A(new_n363), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n239), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n357), .A2(new_n252), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n309), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n223), .B1(new_n711), .B2(new_n332), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n346), .A2(KEYINPUT75), .A3(new_n350), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n352), .B1(new_n337), .B2(new_n349), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n699), .B(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n684), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n453), .B1(new_n566), .B2(new_n571), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n588), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n451), .B(KEYINPUT38), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n719), .B2(new_n720), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n707), .A2(new_n716), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  AOI211_X1 g539(.A(new_n656), .B(new_n660), .C1(new_n517), .C2(new_n653), .ZN(new_n726));
  AOI21_X1  g540(.A(G478), .B1(new_n517), .B2(new_n223), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n572), .B(new_n693), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n700), .A2(new_n642), .A3(new_n701), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  INV_X1    g545(.A(new_n232), .ZN(new_n732));
  INV_X1    g546(.A(new_n592), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n639), .A2(new_n223), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G469), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n732), .A2(new_n641), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n700), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n668), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT105), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n738), .B(new_n740), .ZN(G15));
  NAND3_X1  g555(.A1(new_n700), .A2(new_n677), .A3(new_n736), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT106), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n700), .A2(new_n736), .A3(new_n744), .A4(new_n677), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT107), .B(G116), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G18));
  AOI21_X1  g562(.A(new_n717), .B1(new_n584), .B2(new_n590), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n454), .A2(new_n641), .A3(new_n733), .A4(new_n735), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n700), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT108), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n700), .A2(new_n749), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT109), .B(G119), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G21));
  AOI21_X1  g571(.A(new_n289), .B1(new_n711), .B2(KEYINPUT28), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n336), .B1(new_n758), .B2(new_n332), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(KEYINPUT110), .B(new_n336), .C1(new_n758), .C2(new_n332), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n335), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n338), .ZN(new_n764));
  INV_X1    g578(.A(new_n231), .ZN(new_n765));
  OAI21_X1  g579(.A(G472), .B1(new_n346), .B2(G902), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n641), .A2(new_n735), .A3(new_n733), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n588), .A2(new_n665), .A3(new_n718), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n767), .A2(new_n768), .A3(new_n582), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n465), .ZN(G24));
  AND3_X1   g585(.A1(new_n764), .A2(new_n766), .A3(new_n684), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n728), .A2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n661), .A2(new_n774), .A3(new_n572), .A4(new_n693), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n750), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  NAND2_X1  g591(.A1(new_n451), .A2(new_n666), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n642), .A2(new_n773), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n346), .B2(new_n350), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n337), .A2(KEYINPUT112), .A3(new_n349), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n782), .B(new_n783), .C1(KEYINPUT32), .C2(new_n648), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n369), .A2(G472), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n765), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT42), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n636), .A2(new_n640), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n610), .A2(new_n616), .A3(KEYINPUT83), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT83), .B1(new_n610), .B2(new_n616), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n595), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n627), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n631), .B1(new_n792), .B2(new_n223), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n733), .B(new_n779), .C1(new_n788), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n773), .A2(new_n775), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n371), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(new_n276), .ZN(G33));
  OAI21_X1  g614(.A(new_n699), .B1(new_n714), .B2(new_n715), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n732), .B1(new_n801), .B2(new_n785), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n630), .A2(new_n641), .ZN(new_n803));
  INV_X1    g617(.A(new_n694), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n733), .A4(new_n779), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n802), .A2(new_n805), .A3(KEYINPUT113), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n690), .A2(new_n694), .A3(new_n592), .A4(new_n778), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n807), .B1(new_n371), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n269), .ZN(G36));
  INV_X1    g625(.A(new_n661), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n812), .A2(KEYINPUT43), .A3(new_n572), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n717), .B1(new_n766), .B2(new_n697), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT43), .B1(new_n812), .B2(new_n572), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n778), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n792), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n791), .A2(KEYINPUT45), .A3(new_n627), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(G469), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(G469), .A2(G902), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT46), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n788), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(KEYINPUT46), .A3(new_n824), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n592), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n705), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(new_n271), .ZN(G39));
  XNOR2_X1  g645(.A(new_n828), .B(KEYINPUT47), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n700), .A2(new_n732), .A3(new_n728), .A4(new_n778), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  NAND2_X1  g649(.A1(new_n641), .A2(new_n735), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT115), .Z(new_n838));
  INV_X1    g652(.A(new_n716), .ZN(new_n839));
  INV_X1    g653(.A(new_n722), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(KEYINPUT49), .B2(new_n836), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n592), .A2(new_n453), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n661), .A2(new_n765), .A3(new_n573), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT114), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n836), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n832), .B1(new_n592), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n813), .A2(new_n578), .A3(new_n815), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n767), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n779), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n768), .A2(new_n778), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n772), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n839), .A2(new_n578), .A3(new_n736), .A4(new_n779), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n661), .A2(new_n572), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n855), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n767), .A2(new_n768), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n840), .A2(new_n666), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT50), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n852), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n852), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n850), .A2(new_n750), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT120), .Z(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n870));
  INV_X1    g684(.A(new_n854), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n786), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n856), .A2(new_n662), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n874));
  INV_X1    g688(.A(new_n786), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n854), .A2(new_n874), .A3(KEYINPUT48), .A4(new_n875), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n574), .A2(new_n872), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n866), .A2(new_n867), .A3(new_n869), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n770), .B1(new_n737), .B2(new_n668), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n746), .A2(new_n755), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n810), .A2(new_n799), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n588), .A2(new_n883), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n571), .A2(new_n675), .A3(new_n684), .A4(new_n693), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n587), .A2(KEYINPUT116), .A3(new_n521), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n354), .B2(new_n370), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n690), .A2(new_n592), .A3(new_n778), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n796), .A2(new_n772), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n522), .A2(new_n523), .A3(new_n883), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT116), .B1(new_n587), .B2(new_n521), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT117), .B1(new_n893), .B2(new_n572), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n573), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n667), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n650), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n642), .A2(new_n668), .A3(new_n649), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n687), .ZN(new_n901));
  AND4_X1   g715(.A1(new_n643), .A2(new_n890), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n881), .A2(new_n882), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n683), .B(new_n693), .C1(new_n228), .C2(new_n230), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n588), .A2(new_n665), .A3(new_n718), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AND4_X1   g721(.A1(KEYINPUT118), .A2(new_n716), .A3(new_n642), .A4(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n690), .A2(new_n906), .A3(new_n592), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT118), .B1(new_n909), .B2(new_n716), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n702), .A2(new_n730), .A3(new_n776), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT52), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n716), .A2(new_n642), .A3(new_n907), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(KEYINPUT118), .A3(new_n716), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n454), .A2(new_n641), .A3(new_n733), .A4(new_n735), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n795), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n685), .B1(new_n354), .B2(new_n370), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n772), .A2(new_n920), .B1(new_n921), .B2(new_n695), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT52), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n918), .A2(new_n922), .A3(new_n923), .A4(new_n730), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n913), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n879), .B1(new_n903), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n746), .A2(new_n755), .A3(new_n880), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n787), .B(new_n798), .C1(new_n806), .C2(new_n809), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n890), .A2(new_n643), .A3(new_n899), .A4(new_n901), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n913), .A2(new_n924), .ZN(new_n931));
  INV_X1    g745(.A(new_n922), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT52), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n879), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT54), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n879), .B1(new_n932), .B2(KEYINPUT52), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n930), .A2(new_n931), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n926), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT119), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n937), .A2(new_n941), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT119), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n878), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(G952), .A2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n845), .B1(new_n946), .B2(new_n947), .ZN(G75));
  NOR2_X1   g762(.A1(new_n423), .A2(G952), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n223), .B1(new_n926), .B2(new_n940), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT56), .B1(new_n951), .B2(new_n447), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n417), .A2(new_n418), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(new_n425), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT55), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n950), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n952), .B2(new_n955), .ZN(G51));
  INV_X1    g771(.A(new_n823), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n824), .B(KEYINPUT57), .Z(new_n961));
  INV_X1    g775(.A(new_n941), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n938), .B1(new_n926), .B2(new_n940), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n639), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n949), .B1(new_n960), .B2(new_n965), .ZN(G54));
  NAND3_X1  g780(.A1(new_n951), .A2(KEYINPUT58), .A3(G475), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(new_n561), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n561), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(new_n949), .ZN(G60));
  XNOR2_X1  g784(.A(new_n658), .B(KEYINPUT123), .ZN(new_n971));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT59), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n971), .B(new_n973), .C1(new_n962), .C2(new_n963), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n950), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n945), .A2(new_n943), .A3(new_n973), .ZN(new_n976));
  INV_X1    g790(.A(new_n971), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(G63));
  NAND2_X1  g792(.A1(new_n926), .A2(new_n940), .ZN(new_n979));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT124), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n984), .B(new_n981), .C1(new_n926), .C2(new_n940), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n682), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n939), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n903), .A2(new_n925), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT53), .B1(new_n930), .B2(new_n931), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n984), .ZN(new_n991));
  INV_X1    g805(.A(new_n220), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n979), .A2(KEYINPUT124), .A3(new_n982), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n986), .A2(new_n994), .A3(new_n950), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n986), .A2(new_n994), .A3(KEYINPUT61), .A4(new_n950), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(G66));
  INV_X1    g813(.A(new_n579), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n423), .B1(new_n1000), .B2(G224), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n881), .A2(new_n643), .A3(new_n899), .A4(new_n901), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n1003), .B2(new_n423), .ZN(new_n1004));
  INV_X1    g818(.A(G898), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n953), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G69));
  OAI21_X1  g821(.A(new_n328), .B1(new_n330), .B2(KEYINPUT30), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT126), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n528), .A2(new_n529), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n912), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n724), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n802), .A2(new_n706), .A3(new_n778), .ZN(new_n1018));
  INV_X1    g832(.A(new_n662), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(new_n897), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1016), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1012), .B1(new_n1021), .B2(new_n423), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n423), .B1(G227), .B2(G900), .ZN(new_n1025));
  OR3_X1    g839(.A1(new_n829), .A2(new_n769), .A3(new_n786), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1017), .A2(new_n882), .A3(new_n1013), .A4(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1011), .A2(G953), .ZN(new_n1028));
  AOI22_X1  g842(.A1(new_n1027), .A2(new_n1028), .B1(new_n691), .B2(G953), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1025), .A2(new_n1024), .ZN(new_n1031));
  OR2_X1    g845(.A1(new_n1025), .A2(new_n1024), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1029), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1031), .B(new_n1032), .C1(new_n1022), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n1030), .A2(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  OAI21_X1  g851(.A(new_n1037), .B1(new_n1021), .B2(new_n1003), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n709), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1037), .B1(new_n1003), .B2(new_n1027), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1040), .A2(new_n239), .A3(new_n708), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n364), .A2(new_n333), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n936), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1043));
  AND4_X1   g857(.A1(new_n950), .A2(new_n1039), .A3(new_n1041), .A4(new_n1043), .ZN(G57));
endmodule


