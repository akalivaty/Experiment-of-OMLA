//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT28), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n204), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  OAI211_X1 g009(.A(KEYINPUT67), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(KEYINPUT26), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT67), .B1(new_n218), .B2(new_n207), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n205), .B(new_n206), .C1(new_n214), .C2(new_n219), .ZN(new_n220));
  OR3_X1    g019(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(new_n203), .ZN(new_n224));
  NAND3_X1  g023(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n221), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n212), .B(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT65), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(new_n217), .B2(new_n208), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n227), .B(new_n229), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT25), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  INV_X1    g034(.A(G134gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(G127gat), .ZN(new_n237));
  INV_X1    g036(.A(G127gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT68), .B(G134gat), .Z(new_n240));
  OAI211_X1 g039(.A(new_n237), .B(new_n239), .C1(new_n240), .C2(new_n238), .ZN(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT1), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n242), .B2(new_n243), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT70), .B(G120gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(new_n242), .ZN(new_n247));
  XNOR2_X1  g046(.A(G127gat), .B(G134gat), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n241), .A2(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n229), .A2(new_n251), .A3(new_n218), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n224), .B(new_n225), .C1(G183gat), .C2(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n220), .A2(new_n234), .A3(new_n250), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n220), .A2(new_n234), .A3(new_n254), .ZN(new_n257));
  INV_X1    g056(.A(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g058(.A1(KEYINPUT25), .A2(new_n233), .B1(new_n252), .B2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n250), .A4(new_n220), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G15gat), .B(G43gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT33), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(KEYINPUT32), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n266), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n269), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n266), .B2(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT33), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n277), .A2(KEYINPUT72), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT72), .B1(new_n277), .B2(new_n279), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n256), .A2(new_n259), .A3(new_n262), .A4(new_n264), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT34), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n283), .B2(KEYINPUT34), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(KEYINPUT34), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290));
  INV_X1    g089(.A(new_n288), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n291), .B(new_n275), .C1(new_n280), .C2(new_n281), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n280), .A2(new_n281), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(KEYINPUT76), .A3(new_n291), .A4(new_n275), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT77), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n257), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT77), .B1(new_n260), .B2(new_n220), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT22), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n305), .A3(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n300), .A2(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n257), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n304), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n257), .A2(new_n301), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n260), .A2(KEYINPUT77), .A3(new_n220), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n317), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n260), .A2(new_n220), .A3(new_n300), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n299), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n324), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n315), .ZN(new_n328));
  INV_X1    g127(.A(new_n299), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n319), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n326), .B1(new_n331), .B2(KEYINPUT30), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n328), .A2(new_n319), .A3(KEYINPUT30), .A4(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n333), .A2(new_n334), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n332), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  INV_X1    g138(.A(G85gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT0), .B(G57gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  INV_X1    g145(.A(G148gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(G141gat), .ZN(new_n348));
  INV_X1    g147(.A(G141gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(KEYINPUT81), .A3(G148gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(G141gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353));
  INV_X1    g152(.A(G155gat), .ZN(new_n354));
  INV_X1    g153(.A(G162gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n356), .B2(KEYINPUT2), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n357), .A3(KEYINPUT82), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n349), .A2(G148gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n351), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n351), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n356), .A2(new_n353), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n360), .A2(new_n361), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n250), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n370), .A2(new_n250), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n345), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT5), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(new_n369), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n258), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n344), .B1(new_n380), .B2(new_n371), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT5), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT85), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT83), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n386), .A3(KEYINPUT4), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n388), .A3(new_n250), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT84), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n370), .A2(new_n391), .A3(new_n388), .A4(new_n250), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n385), .A2(new_n387), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n250), .B1(new_n379), .B2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n370), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n345), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n376), .A2(new_n383), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n384), .A2(new_n389), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n394), .A2(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n344), .A2(new_n382), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n343), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n376), .A2(new_n383), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n393), .A2(new_n397), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n343), .ZN(new_n408));
  INV_X1    g207(.A(new_n403), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(KEYINPUT6), .B(new_n343), .C1(new_n398), .C2(new_n403), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n379), .B2(KEYINPUT3), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT29), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n315), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n379), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n315), .B1(new_n396), .B2(new_n417), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(KEYINPUT86), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT3), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n370), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n415), .B1(new_n427), .B2(new_n422), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(G22gat), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n423), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G78gat), .B(G106gat), .Z(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT31), .B(G50gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n423), .B2(new_n428), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT35), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n430), .A2(new_n432), .A3(new_n438), .A4(new_n436), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n338), .A2(new_n414), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n296), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n440), .A2(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n337), .A2(new_n335), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n329), .B1(new_n328), .B2(new_n319), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n330), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n414), .A2(new_n446), .A3(new_n447), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n282), .A2(KEYINPUT75), .A3(new_n288), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT75), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n289), .A2(new_n453), .A3(new_n292), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n445), .B1(new_n455), .B2(new_n441), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n412), .A2(new_n413), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n327), .B2(new_n316), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n304), .A2(new_n315), .A3(new_n318), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT38), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n328), .A2(new_n458), .A3(new_n319), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n299), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n331), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n461), .A2(KEYINPUT89), .A3(new_n299), .A4(new_n462), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n458), .B1(new_n328), .B2(new_n319), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n299), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT38), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n457), .A2(new_n465), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n335), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n450), .B1(new_n471), .B2(new_n336), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n408), .B1(new_n407), .B2(new_n409), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n344), .B1(new_n399), .B2(new_n400), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n372), .A2(new_n373), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n344), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n343), .B1(new_n474), .B2(new_n476), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT40), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT40), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n473), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n472), .A2(new_n483), .A3(KEYINPUT88), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT88), .B1(new_n472), .B2(new_n483), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n470), .B(new_n446), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n446), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n457), .B2(new_n472), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n296), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n454), .A2(KEYINPUT36), .A3(new_n452), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n456), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(G29gat), .A2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n505));
  INV_X1    g304(.A(G29gat), .ZN(new_n506));
  INV_X1    g305(.A(G36gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n497), .B1(new_n508), .B2(new_n499), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n496), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n503), .B(new_n497), .C1(new_n508), .C2(new_n499), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n495), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT17), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT16), .B1(new_n515), .B2(G1gat), .ZN(new_n516));
  INV_X1    g315(.A(G1gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(KEYINPUT90), .ZN(new_n518));
  NOR2_X1   g317(.A1(G15gat), .A2(G22gat), .ZN(new_n519));
  AND2_X1   g318(.A1(G15gat), .A2(G22gat), .ZN(new_n520));
  OAI22_X1  g319(.A1(new_n516), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(G15gat), .A2(G22gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n527), .A3(G8gat), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n521), .B(new_n526), .C1(new_n522), .C2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n495), .B1(new_n532), .B2(new_n512), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n510), .A2(new_n496), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n511), .A2(new_n513), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n528), .A2(new_n530), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT18), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n539), .B(new_n540), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n538), .B(KEYINPUT13), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT11), .B(G169gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  NAND4_X1  g354(.A1(new_n545), .A2(new_n547), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n544), .A2(KEYINPUT18), .B1(new_n548), .B2(new_n549), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(KEYINPUT93), .A3(new_n547), .A4(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n555), .B1(new_n559), .B2(new_n547), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n494), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G57gat), .B(G64gat), .Z(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n566), .A2(new_n572), .A3(new_n570), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n574), .A2(KEYINPUT21), .A3(new_n575), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n531), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n540), .B1(KEYINPUT21), .B2(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT96), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n584), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n583), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT8), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT7), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n340), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n599), .A2(new_n602), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G99gat), .B(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n340), .B2(new_n603), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT97), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n607), .A3(new_n613), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT17), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n539), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT41), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G134gat), .B(G162gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n624), .B(new_n630), .C1(new_n621), .C2(new_n626), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT98), .B1(new_n597), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n592), .A2(new_n596), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G230gat), .ZN(new_n639));
  INV_X1    g438(.A(G233gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n574), .A2(new_n575), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n615), .A2(new_n643), .A3(new_n618), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n574), .B(new_n575), .C1(new_n609), .C2(new_n614), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT10), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND4_X1   g445(.A1(KEYINPUT10), .A2(new_n576), .A3(new_n615), .A4(new_n618), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(new_n641), .A3(new_n645), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n648), .B2(new_n649), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n635), .A2(new_n638), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n565), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n457), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT99), .B(G1gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n472), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n664), .A2(KEYINPUT42), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n664), .B2(G8gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n667), .B2(new_n669), .ZN(G1325gat));
  AOI21_X1  g469(.A(G15gat), .B1(new_n660), .B2(new_n296), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n493), .A2(G15gat), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n660), .B2(new_n672), .ZN(G1326gat));
  NAND2_X1  g472(.A1(new_n660), .A2(new_n487), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(new_n597), .ZN(new_n677));
  INV_X1    g476(.A(new_n657), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n677), .A2(new_n637), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n565), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n506), .A3(new_n457), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n488), .A2(KEYINPUT100), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n338), .A2(new_n414), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n487), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n484), .A2(new_n485), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n446), .B1(new_n688), .B2(new_n414), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n683), .B(new_n686), .C1(new_n687), .C2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n456), .B1(new_n690), .B2(new_n493), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n634), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n494), .A2(KEYINPUT44), .A3(new_n634), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n562), .B1(new_n558), .B2(new_n560), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n677), .A2(new_n696), .A3(new_n678), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n414), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n699), .ZN(G1328gat));
  OAI21_X1  g499(.A(G36gat), .B1(new_n698), .B2(new_n338), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n565), .A2(new_n507), .A3(new_n472), .A4(new_n679), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n705));
  OAI221_X1 g504(.A(new_n701), .B1(KEYINPUT46), .B2(new_n702), .C1(new_n704), .C2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(new_n493), .ZN(new_n707));
  OAI21_X1  g506(.A(G43gat), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(G43gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n680), .A2(new_n709), .A3(new_n296), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n698), .B2(new_n446), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  INV_X1    g516(.A(G50gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n680), .A2(new_n718), .A3(new_n487), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n716), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(G1331gat));
  AND4_X1   g521(.A1(new_n696), .A2(new_n635), .A3(new_n638), .A4(new_n678), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n691), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n457), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g526(.A1(new_n724), .A2(new_n338), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  AND2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n728), .B2(new_n729), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n724), .B2(new_n707), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n296), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n568), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n724), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g537(.A1(new_n724), .A2(new_n446), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n569), .ZN(G1335gat));
  NOR3_X1   g539(.A1(new_n677), .A2(new_n564), .A3(new_n657), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n683), .A2(new_n686), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n742), .A2(new_n491), .A3(new_n492), .A4(new_n486), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n637), .B1(new_n743), .B2(new_n456), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n695), .B(new_n741), .C1(new_n744), .C2(KEYINPUT44), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n414), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n677), .A2(new_n564), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n691), .A2(new_n634), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n657), .B1(new_n748), .B2(KEYINPUT51), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n691), .A2(new_n750), .A3(new_n634), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n457), .A2(new_n340), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n746), .B1(new_n752), .B2(new_n753), .ZN(G1336gat));
  NAND2_X1  g553(.A1(new_n748), .A2(KEYINPUT51), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n338), .A2(G92gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(new_n678), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n749), .A2(KEYINPUT103), .A3(new_n751), .A4(new_n756), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n694), .A2(new_n472), .A3(new_n695), .A4(new_n741), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n766), .A3(new_n751), .A4(new_n756), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT104), .B1(new_n761), .B2(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(new_n757), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n765), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(new_n770), .ZN(G1337gat));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n772));
  OR3_X1    g571(.A1(new_n745), .A2(new_n772), .A3(new_n707), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n745), .B2(new_n707), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(G99gat), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(G99gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n296), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n752), .B2(new_n777), .ZN(G1338gat));
  OAI21_X1  g577(.A(G106gat), .B1(new_n745), .B2(new_n446), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n446), .A2(G106gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n752), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT106), .B(KEYINPUT53), .Z(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n782), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n779), .B(new_n784), .C1(new_n752), .C2(new_n780), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1339gat));
  OR2_X1    g585(.A1(new_n548), .A2(new_n549), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n537), .A2(new_n541), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(G229gat), .A3(G233gat), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n554), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n561), .A2(KEYINPUT109), .A3(new_n678), .A4(new_n791), .ZN(new_n792));
  OR3_X1    g591(.A1(new_n646), .A2(new_n647), .A3(new_n642), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(KEYINPUT54), .A3(new_n648), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n642), .C1(new_n646), .C2(new_n647), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n796), .A2(KEYINPUT107), .A3(new_n652), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT107), .B1(new_n796), .B2(new_n652), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT55), .B(new_n794), .C1(new_n797), .C2(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n654), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n792), .B1(new_n696), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n657), .B(new_n790), .C1(new_n558), .C2(new_n560), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(KEYINPUT109), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT110), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n790), .B1(new_n558), .B2(new_n560), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n678), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n801), .A2(new_n654), .A3(new_n802), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n564), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .A4(new_n792), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n807), .A2(new_n637), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n634), .A2(new_n808), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT108), .B1(new_n817), .B2(new_n803), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n812), .A2(new_n819), .A3(new_n634), .A4(new_n808), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n677), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n658), .A2(new_n564), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n472), .A2(new_n414), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n824), .A2(new_n446), .A3(new_n296), .A4(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n696), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n454), .A2(new_n452), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n824), .A2(new_n828), .A3(new_n446), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n564), .A2(new_n242), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n826), .B2(new_n657), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n678), .A2(new_n246), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n829), .B2(new_n833), .ZN(G1341gat));
  NOR3_X1   g633(.A1(new_n826), .A2(new_n238), .A3(new_n597), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n238), .B1(new_n829), .B2(new_n597), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n836), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(G1342gat));
  OR2_X1    g639(.A1(new_n637), .A2(new_n240), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n829), .A2(KEYINPUT56), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n826), .B2(new_n637), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT56), .B1(new_n829), .B2(new_n841), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n843), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1343gat));
  NOR3_X1   g648(.A1(new_n493), .A2(new_n414), .A3(new_n472), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n851), .B(new_n487), .C1(new_n822), .C2(new_n823), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n803), .A2(new_n696), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n805), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n809), .B(KEYINPUT113), .C1(new_n696), .C2(new_n803), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n637), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n677), .B1(new_n857), .B2(new_n821), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n823), .B1(new_n858), .B2(KEYINPUT114), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n812), .A2(new_n564), .B1(new_n678), .B2(new_n808), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n634), .B1(new_n861), .B2(KEYINPUT113), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n862), .A2(new_n855), .B1(new_n818), .B2(new_n820), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n860), .B1(new_n863), .B2(new_n677), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n446), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n850), .B(new_n852), .C1(new_n865), .C2(new_n851), .ZN(new_n866));
  OAI21_X1  g665(.A(G141gat), .B1(new_n866), .B2(new_n696), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT115), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n487), .B1(new_n822), .B2(new_n823), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(new_n349), .A3(new_n564), .A4(new_n850), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n859), .A2(new_n864), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n851), .B1(new_n872), .B2(new_n487), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n852), .A2(new_n850), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n873), .A2(new_n874), .A3(new_n696), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n875), .B2(new_n349), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n876), .A3(KEYINPUT58), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n867), .B(new_n871), .C1(KEYINPUT115), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n870), .A2(new_n850), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n347), .A3(new_n678), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n817), .A2(new_n803), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n677), .B1(new_n857), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n851), .B(new_n487), .C1(new_n888), .C2(new_n823), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n678), .A3(new_n850), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n884), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n866), .A2(new_n657), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(KEYINPUT59), .A3(new_n347), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n883), .B1(new_n892), .B2(new_n894), .ZN(G1345gat));
  NOR3_X1   g694(.A1(new_n866), .A2(new_n354), .A3(new_n597), .ZN(new_n896));
  AOI21_X1  g695(.A(G155gat), .B1(new_n882), .B2(new_n677), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  NOR3_X1   g697(.A1(new_n866), .A2(new_n355), .A3(new_n637), .ZN(new_n899));
  AOI21_X1  g698(.A(G162gat), .B1(new_n882), .B2(new_n634), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n457), .A2(new_n338), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n735), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n903), .B(new_n446), .C1(new_n822), .C2(new_n823), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n696), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n824), .A2(new_n828), .A3(new_n446), .A4(new_n902), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n696), .A2(G169gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(G1348gat));
  INV_X1    g709(.A(new_n904), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(G176gat), .A3(new_n678), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n906), .A2(new_n657), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(G176gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(G1349gat));
  NAND4_X1  g716(.A1(new_n824), .A2(new_n446), .A3(new_n677), .A4(new_n903), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(KEYINPUT118), .ZN(new_n919));
  OAI21_X1  g718(.A(G183gat), .B1(new_n918), .B2(KEYINPUT118), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n677), .A2(new_n202), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n919), .A2(new_n920), .B1(new_n906), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(KEYINPUT119), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n924), .ZN(new_n926));
  OAI221_X1 g725(.A(new_n926), .B1(new_n906), .B2(new_n921), .C1(new_n919), .C2(new_n920), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n904), .B2(new_n637), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT61), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(KEYINPUT61), .B2(new_n929), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n929), .B2(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n634), .A2(new_n203), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(new_n906), .B2(new_n934), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n493), .A2(new_n457), .A3(new_n338), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n890), .A2(new_n564), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g738(.A(KEYINPUT121), .B(G197gat), .Z(new_n940));
  NAND4_X1  g739(.A1(new_n890), .A2(KEYINPUT122), .A3(new_n564), .A4(new_n936), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n824), .A2(new_n487), .A3(new_n936), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n943), .A2(new_n696), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1352gat));
  OR2_X1    g744(.A1(new_n657), .A2(G204gat), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT62), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT123), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n943), .A2(KEYINPUT62), .A3(new_n946), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n890), .A2(new_n678), .A3(new_n936), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(G204gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n948), .A2(new_n951), .ZN(G1353gat));
  NAND4_X1  g751(.A1(new_n885), .A2(new_n677), .A3(new_n889), .A4(new_n936), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(G211gat), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n953), .A2(new_n959), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n677), .A2(new_n307), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n943), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT124), .Z(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n964), .ZN(G1354gat));
  INV_X1    g764(.A(new_n943), .ZN(new_n966));
  AOI21_X1  g765(.A(G218gat), .B1(new_n966), .B2(new_n634), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n890), .A2(new_n936), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n634), .A2(G218gat), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT127), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n968), .B2(KEYINPUT126), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n967), .B1(new_n969), .B2(new_n972), .ZN(G1355gat));
endmodule


