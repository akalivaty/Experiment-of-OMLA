//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G2106), .B2(new_n453), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT68), .Z(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n470), .A2(new_n473), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n467), .A2(new_n471), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n474), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n471), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .A3(G138), .A4(new_n471), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n463), .A2(G2105), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n496), .A2(G2105), .B1(G102), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n502), .B(new_n504), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G88), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n505), .A2(new_n506), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n502), .A2(new_n504), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n513), .A2(new_n518), .ZN(G166));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n510), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n511), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT70), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n523), .A2(new_n524), .A3(new_n529), .A4(new_n526), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(G168));
  XNOR2_X1  g106(.A(KEYINPUT71), .B(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n511), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n533), .B1(new_n534), .B2(new_n507), .C1(new_n535), .C2(new_n514), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  OR2_X1    g112(.A1(new_n505), .A2(new_n506), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n507), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n515), .A2(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n514), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(KEYINPUT8), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n502), .A2(new_n504), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n508), .B2(G91), .ZN(new_n559));
  OAI211_X1 g134(.A(G53), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(new_n518), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n564), .A2(new_n565), .A3(new_n509), .A4(new_n512), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n509), .B(new_n512), .C1(new_n567), .C2(new_n514), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G303));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n507), .A2(KEYINPUT75), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n511), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT75), .B1(new_n507), .B2(new_n571), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(G288));
  AND3_X1   g151(.A1(new_n502), .A2(new_n504), .A3(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n515), .A2(new_n538), .A3(G86), .ZN(new_n584));
  OAI211_X1 g159(.A(G48), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n583), .A2(KEYINPUT77), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n585), .B1(new_n507), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g164(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT76), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n502), .A2(new_n504), .A3(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n514), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n556), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n508), .A2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n511), .A2(G47), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n556), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(new_n511), .B2(G54), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT10), .B1(new_n507), .B2(new_n610), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n507), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n605), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(G299), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G168), .B2(new_n617), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(G168), .B2(new_n617), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NOR2_X1   g197(.A1(new_n546), .A2(G868), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n613), .A2(G559), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT78), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n623), .B1(new_n625), .B2(G868), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g203(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n474), .A2(G135), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n632), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2435), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2438), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n648), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n641), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n640), .A3(new_n653), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n658), .A3(G14), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT81), .Z(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(KEYINPUT82), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT17), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n661), .B2(new_n663), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  MUX2_X1   g244(.A(new_n669), .B(new_n663), .S(new_n661), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n665), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2096), .ZN(new_n673));
  INV_X1    g248(.A(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n686), .C2(new_n685), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1976), .ZN(new_n704));
  NOR2_X1   g279(.A1(G6), .A2(G16), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n596), .B2(G16), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n698), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n698), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(KEYINPUT34), .B1(new_n704), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n703), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n716), .A2(new_n717), .A3(new_n708), .A4(new_n712), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n474), .A2(G131), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n481), .A2(G119), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n723));
  OR3_X1    g298(.A1(new_n723), .A2(G95), .A3(G2105), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(G95), .B2(G2105), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n471), .A2(G107), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n724), .A2(new_n725), .A3(G2104), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n721), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n720), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT35), .B(G1991), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n730), .B(new_n731), .Z(new_n732));
  NAND4_X1  g307(.A1(new_n714), .A2(new_n718), .A3(KEYINPUT86), .A4(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G24), .ZN(new_n735));
  AND3_X1   g310(.A1(new_n601), .A2(new_n603), .A3(new_n602), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1986), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n734), .A2(KEYINPUT36), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n733), .B2(new_n738), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n481), .A2(G129), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n474), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n497), .A2(G105), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT89), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT26), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT27), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1996), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n719), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n719), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(KEYINPUT96), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(KEYINPUT96), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n759));
  OR3_X1    g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT97), .B(KEYINPUT23), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n698), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G299), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT24), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n719), .B1(new_n770), .B2(G34), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n770), .A2(G34), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G160), .B2(G29), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n776), .A2(new_n777), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT93), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(KEYINPUT93), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n497), .A2(G103), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT25), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(G115), .A2(G2104), .ZN(new_n792));
  INV_X1    g367(.A(G127), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n467), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G2105), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n474), .A2(G139), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n791), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G33), .B(new_n797), .S(G29), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2072), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT31), .B(G11), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT90), .B(G28), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT30), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(new_n719), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n803), .C1(new_n637), .C2(new_n719), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n698), .A2(G19), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n546), .B2(new_n698), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1341), .Z(new_n808));
  NAND4_X1  g383(.A1(new_n769), .A2(new_n788), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G21), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G168), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1966), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n719), .A2(G26), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n481), .A2(G128), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n474), .A2(G140), .ZN(new_n815));
  OR2_X1    g390(.A1(G104), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n719), .ZN(new_n820));
  MUX2_X1   g395(.A(new_n813), .B(new_n820), .S(KEYINPUT28), .Z(new_n821));
  INV_X1    g396(.A(G2067), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n719), .A2(G27), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G164), .B2(new_n719), .ZN(new_n826));
  MUX2_X1   g401(.A(new_n825), .B(new_n826), .S(KEYINPUT94), .Z(new_n827));
  XOR2_X1   g402(.A(KEYINPUT95), .B(G2078), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR4_X1   g404(.A1(new_n809), .A2(new_n812), .A3(new_n824), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n740), .A2(new_n742), .A3(new_n754), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n760), .A2(new_n762), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G2090), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n698), .A2(G4), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n614), .B2(new_n698), .ZN(new_n836));
  INV_X1    g411(.A(G1348), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT91), .B1(G5), .B2(G16), .ZN(new_n840));
  OR3_X1    g415(.A1(KEYINPUT91), .A2(G5), .A3(G16), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n840), .B(new_n841), .C1(G301), .C2(new_n698), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT92), .B(G1961), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR4_X1   g419(.A1(new_n831), .A2(new_n834), .A3(new_n839), .A4(new_n844), .ZN(G311));
  INV_X1    g420(.A(new_n831), .ZN(new_n846));
  INV_X1    g421(.A(new_n844), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n846), .A2(new_n833), .A3(new_n838), .A4(new_n847), .ZN(G150));
  OAI211_X1 g423(.A(G55), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n849));
  INV_X1    g424(.A(G93), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n507), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n502), .A2(new_n504), .A3(G67), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n514), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT99), .B(G860), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NOR2_X1   g434(.A1(new_n613), .A2(new_n621), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT39), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n546), .A2(new_n856), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n855), .B1(new_n542), .B2(new_n545), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n863), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n859), .B1(new_n867), .B2(new_n857), .ZN(G145));
  XNOR2_X1  g443(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n629), .B(KEYINPUT12), .Z(new_n871));
  NAND3_X1  g446(.A1(new_n491), .A2(G130), .A3(G2105), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n491), .A2(G142), .A3(new_n471), .ZN(new_n873));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n874), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n630), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n876), .A2(new_n728), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n728), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n870), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n729), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n876), .A2(new_n728), .A3(new_n878), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n869), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT104), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n497), .A2(G102), .ZN(new_n891));
  INV_X1    g466(.A(new_n495), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n491), .B2(G126), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n893), .B2(new_n471), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n490), .A2(new_n492), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n493), .A2(new_n498), .A3(KEYINPUT100), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n751), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n747), .A2(new_n750), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n896), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n819), .B1(new_n797), .B2(KEYINPUT101), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n795), .A2(new_n796), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n818), .A4(new_n791), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n899), .A3(new_n901), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n888), .A2(new_n889), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n909), .A2(new_n889), .A3(new_n910), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n637), .B1(new_n477), .B2(new_n479), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n477), .A2(new_n479), .A3(new_n637), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n914), .A2(G162), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(G162), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  OAI22_X1  g492(.A1(new_n911), .A2(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n909), .A2(new_n889), .A3(new_n910), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n909), .A2(new_n910), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT104), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT104), .B1(new_n881), .B2(new_n885), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n919), .B(new_n920), .C1(new_n921), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n918), .A2(new_n925), .A3(KEYINPUT105), .A4(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n931), .A2(KEYINPUT106), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(KEYINPUT106), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n932), .B2(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G395));
  NAND2_X1  g512(.A1(new_n856), .A2(new_n617), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n866), .B(KEYINPUT107), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(new_n625), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n558), .A2(G651), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n508), .A2(G91), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT9), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n560), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n941), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n559), .A2(KEYINPUT108), .A3(new_n561), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n614), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n613), .A2(G299), .A3(new_n941), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT41), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n940), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n951), .B(KEYINPUT109), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n940), .A2(new_n957), .ZN(new_n958));
  MUX2_X1   g533(.A(KEYINPUT110), .B(new_n956), .S(new_n958), .Z(new_n959));
  NAND2_X1  g534(.A1(G166), .A2(G290), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n568), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n960), .A2(new_n596), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n596), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g538(.A(G288), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G305), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(new_n596), .A3(new_n961), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n700), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n969), .B1(KEYINPUT111), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n959), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n938), .B1(new_n974), .B2(new_n617), .ZN(G295));
  OAI21_X1  g550(.A(new_n938), .B1(new_n974), .B2(new_n617), .ZN(G331));
  AND3_X1   g551(.A1(new_n528), .A2(new_n530), .A3(G301), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n864), .A2(new_n865), .ZN(new_n978));
  AOI21_X1  g553(.A(G301), .B1(new_n528), .B2(new_n530), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(G168), .A2(G171), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n528), .A2(new_n530), .A3(G301), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n981), .A2(new_n982), .B1(new_n864), .B2(new_n865), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n951), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n866), .A2(new_n982), .A3(new_n981), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n952), .A2(new_n985), .A3(new_n954), .A4(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n984), .A2(new_n987), .A3(new_n969), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n969), .B1(new_n984), .B2(new_n987), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n988), .A2(new_n989), .A3(G37), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT112), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n952), .A2(KEYINPUT113), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n954), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n949), .A2(KEYINPUT113), .A3(new_n953), .A4(new_n950), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n994), .A2(new_n985), .A3(new_n986), .A4(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n980), .A2(new_n983), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n996), .B(new_n969), .C1(new_n957), .C2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n989), .A2(G37), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n991), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n989), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n984), .A2(new_n987), .A3(new_n969), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n926), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT43), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n992), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n998), .A2(KEYINPUT43), .A3(new_n999), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(KEYINPUT43), .B2(new_n990), .ZN(new_n1008));
  MUX2_X1   g583(.A(new_n1006), .B(new_n1008), .S(KEYINPUT44), .Z(G397));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n898), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n470), .A2(new_n473), .A3(new_n475), .A4(G40), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(KEYINPUT114), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(KEYINPUT114), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1996), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n900), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n728), .A2(new_n731), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n728), .A2(new_n731), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n819), .A2(new_n822), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n818), .A2(G2067), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G290), .A2(G1986), .ZN(new_n1027));
  AND2_X1   g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1018), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1014), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n493), .B2(new_n498), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n583), .A2(new_n1036), .A3(new_n584), .A4(new_n585), .ZN(new_n1037));
  OAI21_X1  g612(.A(G1981), .B1(new_n589), .B2(new_n594), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT117), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(G1981), .C1(new_n589), .C2(new_n594), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1039), .A2(KEYINPUT118), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1010), .B1(new_n894), .B2(new_n895), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n1014), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1040), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(KEYINPUT119), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1055), .B(new_n1040), .C1(new_n1039), .C2(new_n1042), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n715), .B(new_n700), .C1(new_n1052), .C2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(new_n1037), .B(KEYINPUT120), .Z(new_n1059));
  AOI21_X1  g634(.A(new_n1035), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n700), .A2(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1061), .B1(new_n1051), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n715), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1051), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1064), .B(new_n1066), .C1(new_n1052), .C2(new_n1057), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(G303), .B2(G8), .ZN(new_n1069));
  OR2_X1    g644(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n1050), .B(new_n1070), .C1(new_n566), .C2(new_n569), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1384), .B1(new_n896), .B2(new_n897), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1014), .B1(new_n1073), .B2(KEYINPUT45), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1048), .A2(new_n1012), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1971), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT115), .B1(new_n1033), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1014), .B1(new_n1033), .B2(new_n1077), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1048), .A2(new_n1080), .A3(KEYINPUT50), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n761), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(G8), .B(new_n1072), .C1(new_n1076), .C2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1067), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1031), .B1(new_n1060), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1053), .B(KEYINPUT119), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1035), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1063), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT100), .B1(new_n493), .B2(new_n498), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n894), .A2(new_n895), .A3(new_n890), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT45), .B(new_n1010), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(new_n1032), .A3(new_n1075), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n711), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1050), .B1(new_n1094), .B2(new_n1082), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1089), .A2(new_n1095), .A3(new_n1072), .A4(new_n1066), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1059), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1976), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n700), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT121), .B(new_n1096), .C1(new_n1099), .C2(new_n1035), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1086), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1077), .B(new_n1010), .C1(new_n894), .C2(new_n895), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1032), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1077), .B1(new_n499), .B2(new_n1010), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1105), .A2(new_n1106), .A3(G2090), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1093), .B2(new_n711), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1103), .B1(new_n1108), .B2(new_n1050), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1109), .A2(new_n1084), .A3(new_n1089), .A4(new_n1066), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1033), .A2(KEYINPUT45), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(new_n1075), .A3(new_n1032), .ZN(new_n1112));
  INV_X1    g687(.A(G1966), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1078), .A2(new_n1079), .A3(new_n783), .A4(new_n1081), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1050), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G168), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1102), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1102), .B1(new_n1119), .B2(new_n1103), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1067), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1117), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1084), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1101), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT122), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1101), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1114), .A2(new_n1115), .A3(G168), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G8), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(KEYINPUT125), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1116), .A2(G286), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1137), .A3(new_n1132), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT62), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1093), .A2(G2078), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(KEYINPUT53), .ZN(new_n1142));
  INV_X1    g717(.A(G1961), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G2078), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT53), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1147), .B2(new_n1112), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1135), .A2(new_n1149), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1140), .A2(G171), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1092), .A2(new_n1032), .A3(new_n1075), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G1956), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT123), .ZN(new_n1157));
  XNOR2_X1  g732(.A(G299), .B(KEYINPUT57), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1144), .A2(new_n837), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1034), .A2(G2067), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n613), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n1157), .A2(new_n1158), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n614), .B(new_n1162), .C1(new_n1144), .C2(new_n837), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT60), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT124), .B(G1996), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT58), .B(G1341), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1093), .A2(new_n1168), .B1(new_n1049), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n546), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(KEYINPUT59), .A3(new_n546), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1161), .A2(new_n1175), .A3(new_n614), .A4(new_n1163), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1167), .A2(new_n1173), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  OR3_X1    g752(.A1(new_n1156), .A2(KEYINPUT61), .A3(new_n1158), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1159), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1160), .B1(new_n1179), .B2(KEYINPUT61), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1165), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G301), .B(KEYINPUT54), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1148), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1183), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1074), .A2(new_n1013), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1145), .B(new_n1185), .C1(new_n1147), .C2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1182), .A2(new_n1184), .A3(new_n1139), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1110), .B1(new_n1151), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1030), .B1(new_n1129), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1018), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(KEYINPUT48), .A3(new_n1027), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1026), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT48), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1027), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1194), .B1(new_n1018), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1192), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1023), .B1(new_n1198), .B2(new_n1022), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1191), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1025), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1191), .B1(new_n900), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1191), .A2(KEYINPUT46), .A3(new_n1019), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT46), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(new_n1018), .B2(G1996), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(KEYINPUT126), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1203), .A2(new_n1204), .A3(new_n1209), .A4(new_n1206), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(KEYINPUT47), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT47), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1208), .A2(new_n1213), .A3(new_n1210), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1201), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1190), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g791(.A1(new_n659), .A2(new_n675), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n1218), .B1(new_n929), .B2(new_n930), .ZN(new_n1219));
  INV_X1    g793(.A(G229), .ZN(new_n1220));
  NAND4_X1  g794(.A1(new_n1006), .A2(new_n1219), .A3(G319), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n1222));
  XNOR2_X1  g796(.A(new_n1221), .B(new_n1222), .ZN(G308));
  XNOR2_X1  g797(.A(new_n1221), .B(KEYINPUT127), .ZN(G225));
endmodule


