//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1198;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT68), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n455), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n468), .B2(G2104), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n479), .A2(G137), .A3(new_n465), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n479), .A2(G2105), .A3(new_n480), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT70), .Z(new_n490));
  NAND4_X1  g065(.A1(new_n480), .A2(new_n478), .A3(new_n465), .A4(new_n469), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI211_X1 g067(.A(new_n486), .B(new_n490), .C1(G136), .C2(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n480), .A2(new_n478), .A3(new_n469), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n467), .A2(new_n469), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n480), .A2(new_n478), .A3(new_n469), .A4(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n506), .A3(new_n503), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n499), .B1(new_n505), .B2(new_n507), .ZN(G164));
  OR2_X1    g083(.A1(KEYINPUT72), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT72), .A2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(KEYINPUT6), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT73), .A3(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n511), .A2(G543), .A3(new_n513), .A4(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  AND4_X1   g095(.A1(new_n511), .A2(new_n513), .A3(new_n520), .A4(new_n516), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n509), .A2(new_n510), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n520), .A2(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT74), .Z(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n519), .A2(new_n522), .A3(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n511), .A2(new_n520), .A3(new_n513), .A4(new_n516), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(G51), .B2(new_n518), .ZN(G168));
  NAND2_X1  g113(.A1(new_n518), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n521), .A2(G90), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n523), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n518), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n521), .A2(G81), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n542), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n517), .A2(KEYINPUT9), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n517), .B2(new_n558), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT76), .B(G65), .Z(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n520), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n515), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(G91), .B2(new_n521), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  NAND3_X1  g143(.A1(new_n521), .A2(KEYINPUT77), .A3(G87), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n535), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g148(.A(KEYINPUT5), .B(G543), .Z(new_n574));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n515), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n518), .B2(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n521), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(new_n523), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n516), .A2(new_n513), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n584), .A2(G48), .A3(G543), .A4(new_n511), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n579), .A2(new_n583), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n542), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT78), .Z(new_n589));
  AOI22_X1  g164(.A1(G47), .A2(new_n518), .B1(new_n521), .B2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n535), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n515), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n598));
  INV_X1    g173(.A(G54), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(new_n517), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n597), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n592), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n592), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n550), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n603), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n497), .A2(new_n473), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(G2100), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n621), .B2(new_n620), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n622), .A2(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n492), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n465), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n487), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n626), .A2(new_n636), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(G2072), .A2(G2078), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n442), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n659), .A2(KEYINPUT85), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(KEYINPUT85), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(new_n661), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n659), .B(KEYINPUT17), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n666), .B(new_n657), .C1(new_n667), .C2(new_n661), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n661), .A3(new_n656), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  NOR3_X1   g258(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  NAND2_X1  g267(.A1(G162), .A2(G29), .ZN(new_n693));
  OR2_X1    g268(.A1(G29), .A2(G35), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G27), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G164), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G2078), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n698), .A2(G2090), .B1(KEYINPUT98), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G2090), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n696), .B2(new_n697), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G34), .ZN(new_n709));
  AOI21_X1  g284(.A(G29), .B1(new_n709), .B2(KEYINPUT24), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(KEYINPUT24), .B2(new_n709), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n482), .B2(new_n699), .ZN(new_n712));
  INV_X1    g287(.A(G2084), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G5), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G171), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n492), .A2(G141), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT93), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n488), .A2(G129), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT26), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n723), .A2(new_n724), .B1(G105), .B2(new_n473), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n719), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(new_n699), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n699), .B2(G32), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n714), .B1(G1961), .B2(new_n717), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT97), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT95), .Z(new_n737));
  INV_X1    g312(.A(new_n635), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n715), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n715), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(G29), .B1(G1966), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(KEYINPUT30), .A2(G28), .ZN(new_n742));
  NAND2_X1  g317(.A1(KEYINPUT30), .A2(G28), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  AOI211_X1 g320(.A(new_n744), .B(new_n745), .C1(new_n717), .C2(G1961), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n741), .B(new_n746), .C1(G1966), .C2(new_n740), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT96), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n699), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n492), .A2(G140), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT92), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G116), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n488), .B2(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2067), .ZN(new_n760));
  INV_X1    g335(.A(G1348), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n604), .A2(new_n715), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G4), .B2(new_n715), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n704), .A2(KEYINPUT98), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n699), .A2(G33), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n497), .A2(G127), .ZN(new_n767));
  INV_X1    g342(.A(G115), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n466), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n770));
  NAND2_X1  g345(.A1(G103), .A2(G2104), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n769), .A2(G2105), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n492), .A2(G139), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n766), .B1(new_n776), .B2(new_n699), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n777), .A2(G2072), .B1(new_n713), .B2(new_n712), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G2072), .B2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n715), .A2(G20), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT23), .Z(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G299), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n715), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n551), .B2(new_n715), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n765), .A2(new_n779), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n764), .B(new_n787), .C1(new_n761), .C2(new_n763), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n708), .A2(new_n735), .A3(new_n749), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G22), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G166), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT90), .B(G1971), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G23), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT89), .ZN(new_n795));
  INV_X1    g370(.A(G288), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(G16), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT33), .B(G1976), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n793), .A2(new_n799), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n806));
  MUX2_X1   g381(.A(G24), .B(G290), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1986), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n699), .A2(G25), .ZN(new_n809));
  INV_X1    g384(.A(G119), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n465), .A2(G107), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n487), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n492), .A2(G131), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n809), .B1(new_n815), .B2(new_n699), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT88), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  OR4_X1    g394(.A1(new_n805), .A2(new_n806), .A3(new_n808), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n821));
  OR2_X1    g396(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n821), .B2(new_n820), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n789), .A2(new_n824), .ZN(G311));
  OR2_X1    g400(.A1(new_n789), .A2(new_n824), .ZN(G150));
  NAND2_X1  g401(.A1(new_n604), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT99), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n518), .A2(G55), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n521), .A2(G93), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n830), .B(new_n831), .C1(new_n542), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n550), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n829), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n835), .A2(KEYINPUT100), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT100), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n833), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(KEYINPUT105), .B(G37), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n776), .A2(KEYINPUT102), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n758), .B1(new_n728), .B2(new_n729), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n726), .A2(new_n727), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n726), .A2(new_n727), .ZN(new_n852));
  INV_X1    g427(.A(new_n758), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n499), .A2(new_n504), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n850), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n850), .B2(new_n854), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n850), .A2(new_n854), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n855), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n850), .A2(new_n854), .A3(new_n856), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n848), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n866));
  INV_X1    g441(.A(G130), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n487), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G142), .B2(new_n492), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n620), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n620), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n815), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n864), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n635), .B(new_n482), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(G162), .Z(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n864), .B2(new_n877), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n846), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n864), .A2(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT104), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n864), .A2(new_n889), .A3(new_n880), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n881), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n884), .ZN(new_n892));
  OAI211_X1 g467(.A(KEYINPUT40), .B(new_n886), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n864), .A2(new_n889), .A3(new_n880), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n889), .B1(new_n864), .B2(new_n880), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n882), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n884), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n898), .B2(new_n886), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n894), .A2(new_n899), .ZN(G395));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n603), .B1(new_n608), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n901), .B2(new_n608), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n603), .A2(KEYINPUT107), .A3(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT108), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n834), .B(KEYINPUT106), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n615), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n905), .B(KEYINPUT41), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  XNOR2_X1  g489(.A(G288), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(G290), .ZN(new_n916));
  XNOR2_X1  g491(.A(G303), .B(G305), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(KEYINPUT110), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n907), .A2(new_n909), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n922), .B(new_n923), .C1(new_n909), .C2(new_n911), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n913), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n921), .B1(new_n913), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n833), .A2(new_n613), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n920), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n918), .A2(KEYINPUT111), .A3(new_n919), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n905), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT41), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n905), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n834), .A2(G171), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n834), .A2(G171), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G168), .ZN(new_n942));
  OAI21_X1  g517(.A(G286), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n936), .A2(new_n938), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n946), .B2(new_n905), .ZN(new_n947));
  AOI21_X1  g522(.A(G37), .B1(new_n934), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n944), .B(new_n920), .C1(new_n946), .C2(new_n905), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT43), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n845), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n906), .A2(new_n945), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n933), .A2(new_n932), .B1(new_n952), .B2(new_n944), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n948), .B2(new_n949), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n951), .A2(new_n953), .A3(KEYINPUT43), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT112), .B(G1384), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n855), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n470), .A2(new_n471), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G2105), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n481), .A2(new_n966), .A3(G40), .A4(new_n474), .ZN(new_n967));
  OR3_X1    g542(.A1(new_n964), .A2(KEYINPUT113), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT113), .B1(new_n964), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(G290), .A2(G1986), .ZN(new_n972));
  AND2_X1   g547(.A1(G290), .A2(G1986), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n851), .A2(new_n852), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n971), .A3(G1996), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT114), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n873), .A2(new_n818), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n873), .A2(new_n818), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n975), .A2(G1996), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n758), .A2(G2067), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n758), .A2(G2067), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n971), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  AND4_X1   g560(.A1(new_n974), .A2(new_n977), .A3(new_n980), .A4(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n499), .B2(new_n504), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n967), .B1(new_n988), .B2(new_n961), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n497), .A2(new_n498), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n501), .A2(new_n506), .A3(new_n503), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n506), .B1(new_n501), .B2(new_n503), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n989), .A2(new_n996), .A3(KEYINPUT53), .A4(new_n702), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n995), .B2(new_n987), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n998), .B(new_n987), .C1(new_n499), .C2(new_n504), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n999), .A2(new_n967), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT124), .B(G1961), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n997), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT45), .B1(new_n995), .B2(new_n987), .ZN(new_n1005));
  INV_X1    g580(.A(G137), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n491), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G40), .ZN(new_n1008));
  NOR4_X1   g583(.A1(new_n1007), .A2(new_n472), .A3(new_n1008), .A4(new_n475), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT45), .B(new_n962), .C1(new_n499), .C2(new_n504), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT53), .B1(new_n1012), .B2(new_n702), .ZN(new_n1013));
  OAI21_X1  g588(.A(G171), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n476), .A2(G40), .A3(new_n713), .A4(new_n481), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n999), .A2(new_n1001), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1966), .B1(new_n989), .B2(new_n996), .ZN(new_n1017));
  OAI21_X1  g592(.A(G286), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1966), .ZN(new_n1019));
  NOR3_X1   g594(.A1(G164), .A2(new_n961), .A3(G1384), .ZN(new_n1020));
  INV_X1    g595(.A(new_n504), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n992), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1009), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1019), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1015), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G164), .A2(G1384), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1000), .B(new_n1025), .C1(new_n1026), .C2(new_n998), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(G168), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1018), .A2(new_n1028), .A3(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT51), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1031), .A3(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1014), .B1(new_n1033), .B2(KEYINPUT62), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT126), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(G166), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1009), .B1(new_n1022), .B2(new_n998), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n995), .A2(new_n998), .A3(new_n987), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT118), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n995), .A2(new_n1044), .A3(new_n998), .A4(new_n987), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n706), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1012), .A2(G1971), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1040), .B1(new_n1050), .B2(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n988), .A2(new_n967), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n1037), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT115), .B(G86), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n583), .B(new_n585), .C1(new_n535), .C2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n579), .A2(new_n583), .A3(new_n1057), .A4(new_n585), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(KEYINPUT117), .B2(KEYINPUT49), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(KEYINPUT116), .A3(new_n1058), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT49), .B1(new_n1063), .B2(KEYINPUT117), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1053), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NOR4_X1   g640(.A1(new_n999), .A2(new_n1001), .A3(G2090), .A4(new_n967), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1040), .B(G8), .C1(new_n1048), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n573), .A2(G1976), .A3(new_n577), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1053), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1053), .A2(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1070), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1065), .A2(new_n1067), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1035), .B1(new_n1051), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1069), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1022), .A2(new_n1009), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G8), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT52), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1074), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1071), .B2(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1063), .A2(KEYINPUT117), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1084), .A2(KEYINPUT49), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n1085), .B2(new_n1053), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1040), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1048), .B1(new_n706), .B2(new_n1046), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1037), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n1089), .A3(KEYINPUT126), .A4(new_n1067), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1030), .A2(new_n1091), .A3(new_n1032), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1034), .A2(new_n1077), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n796), .A2(new_n1073), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1058), .B1(new_n1085), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1067), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1053), .A2(new_n1095), .B1(new_n1086), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1098), .B(new_n1099), .C1(new_n561), .C2(new_n566), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g676(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1102));
  AND4_X1   g677(.A1(new_n561), .A2(new_n566), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1012), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1104), .B(new_n1106), .C1(G1956), .C2(new_n1046), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1079), .A2(G2067), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1009), .B(new_n1000), .C1(new_n1026), .C2(new_n998), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n761), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT121), .B1(new_n1111), .B2(new_n603), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n999), .A2(new_n1001), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1348), .B1(new_n1114), .B2(new_n1009), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1113), .B(new_n604), .C1(new_n1115), .C2(new_n1109), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1106), .B1(new_n1046), .B2(G1956), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1104), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1108), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT61), .B1(new_n1120), .B2(new_n1107), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1109), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(KEYINPUT60), .C1(new_n1002), .C2(G1348), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n604), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n988), .B2(new_n967), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT122), .B(new_n1128), .C1(new_n988), .C2(new_n967), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1005), .A2(new_n1011), .A3(G1996), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n551), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT123), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1110), .A2(new_n761), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n603), .A4(new_n1123), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n551), .B(new_n1137), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1122), .A2(new_n1127), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1120), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1121), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1012), .A2(new_n702), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1003), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1110), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1149), .B(G2078), .C1(new_n967), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1154), .A2(new_n964), .A3(new_n1010), .A4(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1150), .A2(G301), .A3(new_n1152), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1014), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1147), .A2(new_n1158), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1150), .A2(G301), .A3(new_n1152), .A4(new_n997), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1150), .A2(new_n1152), .A3(new_n1156), .ZN(new_n1161));
  OAI211_X1 g736(.A(KEYINPUT54), .B(new_n1160), .C1(new_n1161), .C2(G301), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1159), .A2(new_n1090), .A3(new_n1077), .A4(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1093), .B(new_n1097), .C1(new_n1146), .C2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(G8), .B(G168), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1051), .A2(new_n1076), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n1166), .B2(KEYINPUT119), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1076), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1089), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1170), .B2(new_n1165), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n1172));
  OAI21_X1  g747(.A(G8), .B1(new_n1048), .B2(new_n1066), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1172), .B(new_n1165), .C1(new_n1173), .C2(new_n1087), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1167), .A2(new_n1171), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n986), .B1(new_n1164), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n977), .A2(new_n979), .A3(new_n985), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n970), .B1(new_n1177), .B2(new_n982), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT46), .B1(new_n970), .B2(G1996), .ZN(new_n1179));
  OR3_X1    g754(.A1(new_n970), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n730), .A2(new_n983), .A3(new_n982), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1179), .A2(new_n1180), .B1(new_n1181), .B2(new_n971), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT47), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n971), .A2(new_n972), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  AND4_X1   g760(.A1(new_n980), .A2(new_n977), .A3(new_n985), .A4(new_n1185), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1178), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1176), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1176), .A2(new_n1187), .A3(KEYINPUT127), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g767(.A1(G229), .A2(new_n463), .A3(new_n654), .A4(G227), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n1194), .B1(new_n957), .B2(new_n958), .ZN(new_n1195));
  AND2_X1   g769(.A1(new_n898), .A2(new_n886), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1195), .A2(new_n1196), .ZN(G308));
  NAND2_X1  g771(.A1(new_n898), .A2(new_n886), .ZN(new_n1198));
  OAI211_X1 g772(.A(new_n1198), .B(new_n1194), .C1(new_n957), .C2(new_n958), .ZN(G225));
endmodule


