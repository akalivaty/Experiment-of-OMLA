//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n202), .B(new_n205), .C1(new_n206), .C2(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n202), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n221), .A2(KEYINPUT68), .A3(G120gat), .A4(new_n222), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n221), .A2(G120gat), .A3(new_n222), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G120gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n220), .B(new_n223), .C1(new_n224), .C2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n218), .ZN(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n217), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT67), .B(G113gat), .Z(new_n233));
  AOI21_X1  g032(.A(new_n227), .B1(new_n233), .B2(G120gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n223), .A2(new_n219), .A3(new_n218), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n216), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n237), .A3(KEYINPUT84), .ZN(new_n238));
  NAND2_X1  g037(.A1(G225gat), .A2(G233gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT82), .Z(new_n240));
  INV_X1    g039(.A(KEYINPUT84), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n241), .A3(new_n216), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n216), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n207), .A2(new_n251), .A3(new_n215), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n240), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n236), .B2(new_n216), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n217), .A2(new_n228), .A3(KEYINPUT4), .A4(new_n231), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT83), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n240), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT81), .B1(new_n216), .B2(KEYINPUT3), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n247), .B(new_n251), .C1(new_n207), .C2(new_n215), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(new_n265), .B2(new_n253), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT83), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n266), .A2(new_n267), .A3(new_n259), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n245), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT0), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(KEYINPUT85), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n259), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n255), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n269), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n273), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n267), .B1(new_n266), .B2(new_n259), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n255), .A2(KEYINPUT83), .A3(new_n260), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n244), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n259), .B(KEYINPUT85), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n255), .A2(new_n276), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n279), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n278), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT6), .B(new_n279), .C1(new_n282), .C2(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(G211gat), .A2(G218gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT72), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G211gat), .B(G218gat), .Z(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(KEYINPUT73), .ZN(new_n294));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G204gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(G197gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n290), .A2(KEYINPUT72), .A3(new_n291), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(G197gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n296), .B(new_n295), .C1(new_n302), .C2(new_n292), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n304), .A2(KEYINPUT74), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT74), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n310), .A2(KEYINPUT26), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT27), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT66), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  AOI21_X1  g122(.A(G190gat), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT28), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n321), .A2(new_n326), .A3(G190gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n316), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G169gat), .ZN(new_n329));
  INV_X1    g128(.A(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT25), .A4(new_n314), .ZN(new_n334));
  NOR2_X1   g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n309), .A2(KEYINPUT24), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(G183gat), .A3(G190gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT65), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n331), .A2(new_n333), .A3(new_n314), .ZN(new_n341));
  INV_X1    g140(.A(G190gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n319), .A2(new_n342), .A3(KEYINPUT64), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(G183gat), .B2(G190gat), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n336), .A2(new_n338), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n341), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n340), .B1(new_n348), .B2(KEYINPUT25), .ZN(new_n349));
  INV_X1    g148(.A(new_n335), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n331), .A2(new_n314), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n333), .A2(KEYINPUT25), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n328), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(KEYINPUT76), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n355), .B(new_n340), .C1(KEYINPUT25), .C2(new_n348), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n365), .B2(new_n328), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n366), .B2(new_n361), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  INV_X1    g168(.A(new_n360), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n357), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(KEYINPUT77), .B(new_n360), .C1(new_n365), .C2(new_n328), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n308), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n366), .A2(new_n370), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n377), .A2(new_n378), .B1(new_n357), .B2(new_n361), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n304), .A2(new_n305), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n366), .B2(new_n370), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(KEYINPUT78), .B(new_n308), .C1(new_n368), .C2(new_n373), .ZN(new_n384));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  NAND4_X1  g186(.A1(new_n376), .A2(new_n383), .A3(new_n384), .A4(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n288), .A2(new_n289), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(new_n383), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n363), .B(new_n367), .C1(new_n371), .C2(new_n372), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT78), .B1(new_n392), .B2(new_n308), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n387), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n387), .A2(KEYINPUT30), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n376), .A2(new_n383), .A3(new_n384), .A4(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n394), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n390), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT86), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT86), .B(new_n390), .C1(new_n398), .C2(new_n399), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  INV_X1    g203(.A(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n304), .A2(new_n305), .A3(new_n358), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n251), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n216), .ZN(new_n410));
  INV_X1    g209(.A(G228gat), .ZN(new_n411));
  INV_X1    g210(.A(G233gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n252), .A2(new_n358), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n308), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n308), .A2(KEYINPUT88), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT3), .B1(new_n408), .B2(KEYINPUT87), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n304), .A2(new_n305), .A3(new_n422), .A4(new_n358), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n216), .ZN(new_n425));
  INV_X1    g224(.A(new_n415), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n381), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n413), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(G22gat), .B1(new_n420), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G78gat), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT88), .B1(new_n308), .B2(new_n415), .ZN(new_n432));
  NOR4_X1   g231(.A1(new_n306), .A2(new_n426), .A3(new_n307), .A4(new_n417), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n413), .B(new_n410), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G22gat), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n217), .B1(new_n421), .B2(new_n423), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n436), .A2(new_n427), .B1(new_n411), .B2(new_n412), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n431), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n431), .B1(new_n430), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n407), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n420), .A2(new_n429), .A3(G22gat), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n435), .B1(new_n434), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g243(.A(G78gat), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n439), .A3(new_n406), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n236), .A2(KEYINPUT69), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n236), .A2(KEYINPUT69), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n357), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n365), .A2(KEYINPUT69), .A3(new_n236), .A4(new_n328), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n450), .A2(G227gat), .A3(G233gat), .A4(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(G71gat), .B(G99gat), .Z(new_n453));
  XNOR2_X1  g252(.A(G15gat), .B(G43gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT33), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(KEYINPUT32), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT70), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT70), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n452), .A2(new_n459), .A3(KEYINPUT32), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n450), .A2(new_n451), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n463));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n462), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT32), .ZN(new_n468));
  INV_X1    g267(.A(new_n452), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n468), .B(new_n455), .C1(new_n469), .C2(KEYINPUT33), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n461), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n467), .B1(new_n461), .B2(new_n470), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n447), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n402), .A2(new_n403), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT35), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n394), .A2(new_n397), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n388), .A2(new_n389), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n288), .A2(new_n289), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT35), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n442), .A2(new_n446), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT71), .B1(new_n471), .B2(new_n472), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n461), .A2(new_n467), .A3(new_n470), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n481), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n476), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n402), .A2(new_n403), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n447), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n394), .A2(new_n397), .B1(new_n388), .B2(new_n389), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n265), .A2(new_n253), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n240), .B1(new_n283), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT39), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n238), .A2(new_n242), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(new_n262), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n496), .B(new_n240), .C1(new_n283), .C2(new_n494), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n273), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(KEYINPUT40), .A3(new_n273), .A4(new_n500), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n286), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n446), .B(new_n442), .C1(new_n493), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n288), .A2(new_n289), .A3(new_n388), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n376), .A2(new_n508), .A3(new_n383), .A4(new_n384), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n392), .A2(new_n308), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n381), .B1(new_n379), .B2(new_n382), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT37), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n387), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT38), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT37), .B1(new_n391), .B2(new_n393), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(new_n509), .A3(KEYINPUT38), .A4(new_n513), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n507), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT36), .B1(new_n483), .B2(new_n486), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n473), .A2(new_n521), .ZN(new_n522));
  OAI22_X1  g321(.A1(new_n506), .A2(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n492), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n490), .A2(new_n525), .A3(KEYINPUT89), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n488), .B1(KEYINPUT35), .B2(new_n475), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n482), .B1(new_n402), .B2(new_n403), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n523), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G57gat), .B(G64gat), .Z(new_n533));
  INV_X1    g332(.A(KEYINPUT9), .ZN(new_n534));
  INV_X1    g333(.A(G71gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n431), .ZN(new_n536));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n533), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT94), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n540), .A2(new_n533), .A3(KEYINPUT94), .A4(new_n536), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT95), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT97), .ZN(new_n550));
  XOR2_X1   g349(.A(G127gat), .B(G155gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT98), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n550), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT16), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(G1gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(G1gat), .B2(new_n558), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(G8gat), .Z(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n545), .B2(new_n546), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n563), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n557), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n555), .A2(new_n567), .A3(new_n556), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR3_X1   g370(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(KEYINPUT91), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(KEYINPUT91), .B2(new_n573), .ZN(new_n575));
  INV_X1    g374(.A(G29gat), .ZN(new_n576));
  INV_X1    g375(.A(G36gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G50gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G43gat), .ZN(new_n580));
  INV_X1    g379(.A(G43gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G50gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n582), .A3(KEYINPUT15), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT92), .B1(new_n581), .B2(G50gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(G43gat), .B2(new_n579), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n581), .A2(KEYINPUT92), .A3(G50gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT15), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n573), .ZN(new_n590));
  OAI221_X1 g389(.A(new_n583), .B1(new_n576), .B2(new_n577), .C1(new_n590), .C2(new_n572), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n594), .A2(KEYINPUT17), .ZN(new_n595));
  INV_X1    g394(.A(G99gat), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT8), .B1(new_n596), .B2(new_n405), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT101), .ZN(new_n599));
  OAI221_X1 g398(.A(new_n597), .B1(G85gat), .B2(G92gat), .C1(KEYINPUT7), .C2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT7), .B1(new_n598), .B2(KEYINPUT101), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(KEYINPUT101), .B2(new_n598), .ZN(new_n602));
  XOR2_X1   g401(.A(G99gat), .B(G106gat), .Z(new_n603));
  OR3_X1    g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n600), .B2(new_n602), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n594), .A2(KEYINPUT17), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n595), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n606), .ZN(new_n609));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n609), .A2(new_n593), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT100), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n571), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n545), .A2(new_n625), .A3(new_n606), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n606), .A2(new_n544), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n545), .B2(new_n609), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT102), .B(KEYINPUT10), .Z(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n627), .B(new_n631), .C1(new_n545), .C2(new_n609), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n562), .B(new_n593), .Z(new_n643));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT13), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n594), .A2(new_n562), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n607), .A2(new_n562), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n595), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n644), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT18), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G169gat), .B(G197gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT12), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n652), .B2(KEYINPUT93), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n653), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n624), .A2(new_n642), .A3(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n532), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n480), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n479), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT103), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  MUX2_X1   g472(.A(KEYINPUT103), .B(new_n672), .S(new_n673), .Z(new_n674));
  NOR2_X1   g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n670), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(G8gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(new_n667), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n520), .A2(new_n522), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n487), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n680), .B2(new_n685), .ZN(G1326gat));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n687), .A3(new_n447), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n667), .B2(new_n447), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT105), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n690), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n688), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n695), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n623), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n526), .A2(new_n531), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n571), .A2(new_n642), .A3(new_n665), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n576), .A3(new_n480), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n524), .B1(new_n529), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n492), .A2(KEYINPUT107), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n490), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n699), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n700), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT106), .B1(new_n700), .B2(KEYINPUT44), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(new_n702), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(new_n480), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n706), .B1(new_n717), .B2(new_n576), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n704), .A2(new_n577), .A3(new_n479), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n716), .A2(new_n479), .ZN(new_n724));
  OAI221_X1 g523(.A(new_n723), .B1(new_n721), .B2(new_n719), .C1(new_n724), .C2(new_n577), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n715), .A2(new_n681), .A3(new_n702), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G43gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n704), .A2(new_n581), .A3(new_n487), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT47), .B1(new_n729), .B2(KEYINPUT110), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n731), .B(new_n732), .C1(new_n727), .C2(new_n728), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n733), .ZN(G1330gat));
  NAND3_X1  g533(.A1(new_n716), .A2(G50gat), .A3(new_n447), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n704), .A2(KEYINPUT111), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n447), .B1(new_n703), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n579), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT48), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n735), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1331gat));
  NOR3_X1   g543(.A1(new_n624), .A2(new_n641), .A3(new_n664), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(new_n710), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n480), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT112), .B(G57gat), .Z(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n479), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT49), .B(G64gat), .Z(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(G1333gat));
  AOI21_X1  g552(.A(new_n535), .B1(new_n746), .B2(new_n681), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n684), .A2(G71gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n746), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n746), .A2(new_n447), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n571), .A2(new_n664), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n642), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n700), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n767), .B2(new_n712), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n480), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n760), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(KEYINPUT113), .A3(new_n480), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n772), .A3(G85gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n710), .A2(new_n699), .A3(new_n761), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT51), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n710), .A2(new_n776), .A3(new_n699), .A4(new_n761), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(new_n642), .ZN(new_n779));
  INV_X1    g578(.A(G85gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n480), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n773), .A2(new_n781), .ZN(G1336gat));
  OR3_X1    g581(.A1(new_n641), .A2(G92gat), .A3(new_n493), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT114), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(new_n778), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n762), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n715), .A2(new_n479), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(G92gat), .ZN(new_n794));
  NOR2_X1   g593(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n774), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n774), .A2(new_n795), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n784), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n793), .A2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n769), .B2(new_n682), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n779), .A2(new_n596), .A3(new_n487), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1338gat));
  AOI21_X1  g603(.A(new_n405), .B1(new_n768), .B2(new_n447), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n482), .A2(G106gat), .A3(new_n641), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n796), .B2(new_n797), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT117), .B(KEYINPUT53), .C1(new_n805), .C2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n715), .A2(new_n447), .A3(new_n787), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(G106gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(G106gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n775), .A2(new_n777), .A3(new_n806), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  AOI211_X1 g619(.A(new_n820), .B(new_n817), .C1(new_n811), .C2(G106gat), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n809), .B(new_n814), .C1(new_n819), .C2(new_n821), .ZN(G1339gat));
  AND2_X1   g621(.A1(new_n569), .A2(new_n570), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n632), .A2(KEYINPUT54), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n630), .A2(new_n631), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n632), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n638), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n640), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n638), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n664), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n649), .A2(new_n644), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n643), .A2(new_n645), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n658), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n653), .A2(new_n659), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n642), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n699), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  AND4_X1   g637(.A1(new_n699), .A2(new_n831), .A3(new_n835), .A4(new_n836), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n823), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n571), .A2(new_n623), .A3(new_n641), .A4(new_n665), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n770), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(new_n493), .A3(new_n474), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n664), .A2(new_n233), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT119), .Z(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n770), .A2(new_n479), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(new_n684), .A3(new_n447), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n665), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n854), .ZN(G1340gat));
  INV_X1    g654(.A(G120gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n852), .B2(new_n642), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT120), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n845), .A2(new_n856), .A3(new_n642), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n861), .A3(new_n571), .ZN(new_n862));
  OAI21_X1  g661(.A(G127gat), .B1(new_n853), .B2(new_n823), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1342gat));
  INV_X1    g663(.A(G134gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n845), .A2(new_n865), .A3(new_n699), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n853), .B2(new_n623), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G1343gat));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n842), .B2(new_n447), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n872), .B(new_n482), .C1(new_n840), .C2(new_n841), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n681), .A2(new_n850), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n842), .A2(KEYINPUT57), .A3(new_n447), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n875), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n880), .A3(new_n664), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n879), .B1(new_n875), .B2(new_n874), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(KEYINPUT122), .A3(new_n664), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(G141gat), .A3(new_n885), .ZN(new_n886));
  AND4_X1   g685(.A1(new_n447), .A2(new_n844), .A3(new_n682), .A4(new_n493), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(new_n208), .A3(new_n664), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n208), .B1(new_n884), .B2(new_n664), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT58), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1344gat));
  NAND3_X1  g692(.A1(new_n887), .A2(new_n210), .A3(new_n642), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT123), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT59), .B(new_n210), .C1(new_n884), .C2(new_n642), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n871), .A2(new_n873), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n642), .A3(new_n877), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n895), .B1(new_n896), .B2(new_n900), .ZN(G1345gat));
  INV_X1    g700(.A(new_n884), .ZN(new_n902));
  OAI21_X1  g701(.A(G155gat), .B1(new_n902), .B2(new_n823), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n203), .A3(new_n571), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1346gat));
  OAI21_X1  g704(.A(G162gat), .B1(new_n902), .B2(new_n623), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n204), .A3(new_n699), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n493), .A2(new_n480), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n842), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n474), .ZN(new_n911));
  AOI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n664), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n684), .A2(new_n447), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(new_n329), .A3(new_n665), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n915), .ZN(G1348gat));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n330), .A3(new_n642), .ZN(new_n917));
  OAI21_X1  g716(.A(G176gat), .B1(new_n914), .B2(new_n641), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1349gat));
  NAND4_X1  g718(.A1(new_n911), .A2(new_n318), .A3(new_n320), .A4(new_n571), .ZN(new_n920));
  OAI21_X1  g719(.A(G183gat), .B1(new_n914), .B2(new_n823), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g721(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n911), .A2(new_n342), .A3(new_n699), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n913), .A3(new_n699), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(G190gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n926), .B2(G190gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT125), .Z(G1351gat));
  XNOR2_X1  g730(.A(KEYINPUT126), .B(G197gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n682), .A2(new_n909), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n898), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n936), .B2(new_n665), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n843), .A2(new_n482), .A3(new_n934), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n664), .A3(new_n932), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1352gat));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n298), .A3(new_n642), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT62), .Z(new_n942));
  OAI21_X1  g741(.A(G204gat), .B1(new_n936), .B2(new_n641), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1353gat));
  INV_X1    g743(.A(G211gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n938), .A2(new_n945), .A3(new_n571), .ZN(new_n946));
  INV_X1    g745(.A(new_n936), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n571), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  NAND2_X1  g750(.A1(new_n938), .A2(new_n699), .ZN(new_n952));
  INV_X1    g751(.A(G218gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n623), .A2(new_n953), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n955), .A2(new_n956), .B1(new_n947), .B2(new_n957), .ZN(G1355gat));
endmodule


