//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n187));
  INV_X1    g001(.A(G478), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT15), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT9), .B(G234), .ZN(new_n191));
  INV_X1    g005(.A(G217), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n191), .A2(new_n192), .A3(G953), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT93), .B1(new_n195), .B2(G128), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT93), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT94), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n196), .A2(new_n199), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT13), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n195), .A2(KEYINPUT13), .A3(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(G134), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT94), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n200), .A2(new_n211), .A3(new_n201), .A4(new_n202), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G122), .ZN(new_n216));
  INV_X1    g030(.A(G122), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G116), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT91), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT91), .B1(new_n216), .B2(new_n218), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n218), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT91), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT91), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G107), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT92), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n221), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n213), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(KEYINPUT14), .A3(G122), .ZN(new_n232));
  OAI211_X1 g046(.A(G107), .B(new_n232), .C1(new_n222), .C2(KEYINPUT14), .ZN(new_n233));
  INV_X1    g047(.A(new_n203), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n201), .B1(new_n200), .B2(new_n202), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n221), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n194), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n204), .A2(new_n210), .A3(new_n212), .ZN(new_n239));
  INV_X1    g053(.A(new_n230), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n229), .B1(new_n221), .B2(new_n226), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n236), .A3(new_n193), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G902), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n190), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI211_X1 g060(.A(G902), .B(new_n189), .C1(new_n238), .C2(new_n243), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G140), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G125), .ZN(new_n250));
  INV_X1    g064(.A(G125), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G140), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT81), .A4(KEYINPUT16), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT16), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT81), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n250), .B2(KEYINPUT16), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G214), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n195), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT17), .A3(G131), .ZN(new_n266));
  INV_X1    g080(.A(G146), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n253), .C1(new_n254), .C2(new_n256), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT90), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n262), .A2(new_n271), .A3(new_n264), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT88), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n265), .A2(G131), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n262), .A2(KEYINPUT88), .A3(new_n271), .A4(new_n264), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT90), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n258), .A2(new_n266), .A3(new_n280), .A4(new_n268), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n270), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G113), .B(G122), .ZN(new_n283));
  INV_X1    g097(.A(G104), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n250), .A2(new_n252), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(new_n267), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT18), .A2(G131), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n262), .A2(new_n264), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n265), .A2(KEYINPUT18), .A3(G131), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n282), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n285), .B1(new_n282), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n245), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G475), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n282), .A2(new_n285), .A3(new_n291), .ZN(new_n297));
  AND2_X1   g111(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n286), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n258), .B1(new_n301), .B2(G146), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n291), .B1(new_n302), .B2(new_n277), .ZN(new_n303));
  INV_X1    g117(.A(new_n285), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G475), .A2(G902), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n296), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n307), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT20), .B(new_n309), .C1(new_n297), .C2(new_n305), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n248), .B(new_n295), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G952), .ZN(new_n312));
  AOI211_X1 g126(.A(G953), .B(new_n312), .C1(G234), .C2(G237), .ZN(new_n313));
  AOI211_X1 g127(.A(new_n245), .B(new_n260), .C1(G234), .C2(G237), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT21), .B(G898), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n187), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n297), .A2(new_n305), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT20), .B1(new_n318), .B2(new_n309), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n306), .A2(new_n296), .A3(new_n307), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n319), .A2(new_n320), .B1(G475), .B2(new_n294), .ZN(new_n321));
  INV_X1    g135(.A(new_n316), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(KEYINPUT95), .A3(new_n322), .A4(new_n248), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G122), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT2), .B(G113), .Z(new_n329));
  XNOR2_X1  g143(.A(G116), .B(G119), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n329), .A2(new_n330), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(new_n284), .B2(G107), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n214), .A3(G104), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n284), .A2(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n340));
  INV_X1    g154(.A(G101), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n334), .A2(new_n336), .A3(new_n341), .A4(new_n337), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT83), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n342), .A2(KEYINPUT4), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n339), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n333), .B(new_n340), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n330), .A2(KEYINPUT5), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n215), .A2(KEYINPUT5), .A3(G119), .ZN(new_n350));
  INV_X1    g164(.A(G113), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n349), .A2(new_n352), .B1(new_n329), .B2(new_n330), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n284), .A2(G107), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n214), .A2(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(G101), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n342), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n328), .B1(new_n348), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n361));
  INV_X1    g175(.A(new_n333), .ZN(new_n362));
  INV_X1    g176(.A(new_n340), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n346), .B1(new_n345), .B2(new_n339), .ZN(new_n364));
  AND4_X1   g178(.A1(new_n346), .A2(new_n339), .A3(KEYINPUT4), .A4(new_n342), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n359), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n327), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT6), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(KEYINPUT6), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n327), .B1(new_n366), .B2(new_n367), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT6), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n373), .B(new_n328), .C1(new_n348), .C2(new_n359), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT84), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n369), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n267), .A2(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n195), .A2(G146), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n195), .A2(G146), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n267), .B2(G143), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n195), .A2(KEYINPUT65), .A3(G146), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n198), .B1(new_n378), .B2(KEYINPUT1), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n380), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n387), .A2(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n378), .A2(new_n379), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT0), .A2(G128), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(KEYINPUT64), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT64), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT0), .A3(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT0), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n198), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n392), .B1(new_n399), .B2(new_n385), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n393), .A2(new_n395), .B1(new_n397), .B2(new_n198), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n383), .A2(new_n384), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT66), .B(new_n401), .C1(new_n402), .C2(new_n381), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n391), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n388), .B1(new_n404), .B2(new_n251), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n260), .A2(G224), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n376), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n388), .B(new_n406), .C1(new_n404), .C2(new_n251), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT7), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n411), .A2(KEYINPUT87), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n342), .A2(new_n357), .A3(KEYINPUT85), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n353), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n353), .A2(new_n414), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n327), .B(KEYINPUT8), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT86), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(new_n420), .A3(new_n416), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n406), .A2(KEYINPUT7), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n419), .A2(new_n421), .B1(new_n405), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT87), .B1(new_n411), .B2(new_n412), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n413), .A2(new_n423), .A3(new_n368), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n245), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n409), .A2(new_n410), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n410), .ZN(new_n429));
  OAI211_X1 g243(.A(KEYINPUT84), .B(new_n374), .C1(new_n370), .C2(new_n371), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n407), .B1(new_n430), .B2(new_n369), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n429), .B1(new_n431), .B2(new_n426), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n326), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G221), .ZN(new_n434));
  INV_X1    g248(.A(new_n191), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n245), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G469), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n378), .A2(KEYINPUT1), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n389), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n380), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n342), .A2(new_n357), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n387), .B2(new_n443), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT67), .B1(new_n201), .B2(G137), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT11), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G134), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(KEYINPUT67), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n201), .A2(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT69), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n446), .A2(KEYINPUT11), .B1(new_n201), .B2(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT69), .A3(new_n451), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n455), .A2(KEYINPUT70), .A3(G131), .A4(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n447), .A2(new_n451), .A3(new_n271), .A4(new_n452), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n456), .A2(new_n461), .A3(new_n271), .A4(new_n451), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n271), .B1(new_n453), .B2(new_n454), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT70), .B1(new_n465), .B2(new_n457), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n445), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n455), .A2(G131), .A3(new_n457), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n463), .A3(new_n458), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT12), .A3(new_n445), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G110), .B(G140), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n260), .A2(G227), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n443), .A2(new_n387), .A3(KEYINPUT10), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n358), .B1(new_n380), .B2(new_n441), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(KEYINPUT10), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n340), .B1(new_n344), .B2(new_n347), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n404), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n464), .A2(new_n466), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n478), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n478), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n404), .B(new_n363), .C1(new_n364), .C2(new_n365), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n387), .A2(KEYINPUT10), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n489), .A2(new_n443), .B1(new_n444), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n473), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n488), .A3(new_n491), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n438), .B(new_n245), .C1(new_n486), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n485), .A2(new_n493), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n469), .A2(new_n474), .B1(new_n484), .B2(new_n483), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(new_n487), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n438), .B1(new_n500), .B2(new_n245), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n437), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n324), .A2(new_n433), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT32), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n271), .B1(new_n449), .B2(new_n452), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n508), .B(KEYINPUT72), .Z(new_n509));
  NAND3_X1  g323(.A1(new_n463), .A2(new_n509), .A3(new_n387), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n473), .B2(new_n404), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n404), .B1(new_n464), .B2(new_n466), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n473), .A2(KEYINPUT71), .A3(new_n404), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n362), .B(new_n513), .C1(new_n518), .C2(KEYINPUT30), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n514), .A2(new_n333), .A3(new_n510), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n263), .A2(G210), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n521), .B(KEYINPUT27), .Z(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT26), .B(G101), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n522), .B(new_n523), .Z(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n519), .A2(KEYINPUT31), .A3(new_n520), .A4(new_n524), .ZN(new_n528));
  INV_X1    g342(.A(new_n524), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n516), .A2(new_n517), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n333), .B1(new_n530), .B2(new_n510), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n520), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n514), .A2(KEYINPUT28), .A3(new_n333), .A4(new_n510), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n529), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n534), .B(new_n533), .C1(new_n518), .C2(new_n333), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n529), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n527), .A2(new_n528), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n507), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n527), .A2(new_n528), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n537), .A2(new_n540), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n543), .A2(new_n507), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n520), .B(KEYINPUT74), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT75), .B1(new_n512), .B2(new_n333), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n514), .A2(new_n510), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n362), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT28), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n533), .B(KEYINPUT76), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT29), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n529), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n245), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n558), .B1(new_n538), .B2(new_n529), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n524), .B1(new_n519), .B2(new_n520), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G472), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n544), .A2(new_n549), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n198), .A2(G119), .ZN(new_n567));
  INV_X1    g381(.A(G119), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT24), .B(G110), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT79), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n258), .A2(new_n268), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT80), .B1(new_n198), .B2(G119), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT23), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n569), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G110), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n570), .A2(new_n571), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n579), .B2(G110), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n286), .A2(new_n267), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n258), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n581), .A2(new_n585), .A3(new_n589), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n245), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n594));
  NAND2_X1  g408(.A1(G217), .A2(G902), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n192), .B2(G234), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT77), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT78), .Z(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT25), .B1(new_n593), .B2(KEYINPUT82), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n591), .A2(new_n592), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n597), .A2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n324), .A2(KEYINPUT96), .A3(new_n503), .A4(new_n433), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n506), .A2(new_n566), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  AOI21_X1  g422(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n547), .A2(new_n245), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(G472), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n503), .A2(new_n605), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n231), .A2(new_n237), .A3(new_n194), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n193), .B1(new_n242), .B2(new_n236), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n245), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n188), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT33), .B1(new_n238), .B2(new_n243), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n231), .B2(new_n237), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n242), .A2(KEYINPUT97), .A3(new_n236), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n194), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n621), .A2(new_n622), .A3(KEYINPUT98), .A4(new_n194), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n243), .A2(KEYINPUT33), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n188), .A2(G902), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n618), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n321), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n433), .A3(new_n322), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n613), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n616), .A2(new_n189), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n244), .A2(new_n245), .A3(new_n190), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n640), .B(new_n295), .C1(new_n308), .C2(new_n310), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT99), .B1(new_n641), .B2(new_n316), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n321), .A2(new_n643), .A3(new_n322), .A4(new_n640), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n433), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n613), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n586), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n604), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(new_n599), .B2(new_n600), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n506), .A2(new_n611), .A3(new_n606), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n313), .B1(new_n314), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n641), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n428), .A2(new_n432), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n325), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n653), .B(new_n437), .C1(new_n497), .C2(new_n501), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n566), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XOR2_X1   g479(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n660), .B(new_n666), .ZN(new_n667));
  NOR4_X1   g481(.A1(new_n667), .A2(new_n326), .A3(new_n248), .A4(new_n321), .ZN(new_n668));
  OR3_X1    g482(.A1(new_n550), .A2(new_n555), .A3(new_n524), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n245), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n529), .B1(new_n519), .B2(new_n520), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n548), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n672), .B1(new_n541), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n544), .ZN(new_n676));
  INV_X1    g490(.A(new_n653), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n668), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(KEYINPUT101), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n658), .B(new_n681), .Z(new_n682));
  OR2_X1    g496(.A1(new_n502), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT40), .Z(new_n684));
  NAND3_X1  g498(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT103), .B(G143), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G45));
  OAI21_X1  g501(.A(new_n295), .B1(new_n308), .B2(new_n310), .ZN(new_n688));
  INV_X1    g502(.A(new_n658), .ZN(new_n689));
  INV_X1    g503(.A(new_n630), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n690), .B(new_n619), .C1(new_n627), .C2(new_n628), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n688), .B(new_n689), .C1(new_n691), .C2(new_n618), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n566), .A2(new_n663), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND2_X1  g509(.A1(new_n493), .A2(new_n494), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(new_n478), .B1(new_n475), .B2(new_n485), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n496), .ZN(new_n700));
  OAI211_X1 g514(.A(KEYINPUT104), .B(G469), .C1(new_n697), .C2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n605), .A3(new_n437), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n633), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n566), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT41), .B(G113), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT105), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G15));
  NOR2_X1   g522(.A1(new_n645), .A2(new_n703), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n566), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT106), .B(G116), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G18));
  AOI21_X1  g526(.A(new_n677), .B1(new_n317), .B2(new_n323), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n702), .A2(new_n437), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n661), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n566), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NAND2_X1  g531(.A1(new_n556), .A2(new_n557), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n529), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n545), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n610), .A2(G472), .B1(new_n542), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n436), .B1(new_n700), .B2(new_n701), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n321), .A2(new_n248), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n433), .A3(new_n322), .A4(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n721), .A2(KEYINPUT107), .A3(new_n605), .A4(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  OAI21_X1  g541(.A(G472), .B1(new_n541), .B2(G902), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n720), .A2(new_n542), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n605), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n727), .B1(new_n730), .B2(new_n724), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NOR3_X1   g547(.A1(new_n714), .A2(new_n661), .A3(new_n692), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n728), .A3(new_n653), .A4(new_n729), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  NAND3_X1  g550(.A1(new_n428), .A2(new_n325), .A3(new_n432), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n692), .A2(new_n737), .A3(new_n502), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n547), .A2(new_n740), .A3(new_n548), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT108), .B1(new_n541), .B2(new_n673), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n565), .B1(new_n609), .B2(KEYINPUT32), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n605), .B(new_n739), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n741), .A2(new_n544), .A3(new_n742), .A4(new_n565), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n605), .A4(new_n739), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n737), .A2(new_n502), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n566), .A2(new_n605), .A3(new_n693), .A4(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n746), .A2(new_n749), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT110), .B(G131), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G33));
  NAND4_X1  g568(.A1(new_n566), .A2(new_n605), .A3(new_n659), .A4(new_n750), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  NOR2_X1   g570(.A1(new_n631), .A2(new_n688), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n611), .A2(new_n759), .A3(new_n677), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n761));
  INV_X1    g575(.A(new_n737), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n438), .B1(new_n500), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n764), .B2(new_n500), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n438), .A2(new_n245), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(KEYINPUT46), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n496), .B1(new_n769), .B2(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n437), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n682), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  XOR2_X1   g589(.A(new_n772), .B(KEYINPUT47), .Z(new_n776));
  INV_X1    g590(.A(new_n566), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n692), .A2(new_n737), .A3(new_n605), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n566), .B1(new_n704), .B2(new_n709), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n716), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n728), .A2(new_n729), .A3(new_n653), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n692), .A2(new_n737), .A3(new_n502), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n428), .A2(new_n432), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n311), .A2(new_n658), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(KEYINPUT113), .A3(new_n325), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n662), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n321), .A2(new_n248), .A3(new_n689), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n790), .B1(new_n737), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n788), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n784), .A2(new_n785), .B1(new_n793), .B2(new_n566), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n783), .A2(new_n732), .A3(new_n755), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n752), .ZN(new_n796));
  INV_X1    g610(.A(new_n723), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n437), .B(new_n689), .C1(new_n497), .C2(new_n501), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n661), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n609), .A2(KEYINPUT32), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n799), .B(new_n677), .C1(new_n800), .C2(new_n674), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n664), .A2(new_n694), .A3(new_n735), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n633), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n632), .A2(new_n433), .A3(KEYINPUT111), .A4(new_n322), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n611), .A2(new_n612), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n607), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n607), .A2(new_n808), .A3(KEYINPUT112), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n661), .A2(new_n316), .A3(new_n641), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n611), .A2(new_n612), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n654), .A2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n811), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n796), .A2(new_n804), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n811), .A2(new_n812), .A3(new_n815), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n752), .A3(new_n795), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n664), .A2(new_n735), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT52), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n818), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n804), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n781), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n818), .B1(new_n822), .B2(KEYINPUT52), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n796), .A2(new_n804), .A3(new_n816), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n819), .A2(new_n781), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n831), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT114), .B1(new_n833), .B2(new_n826), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n667), .A2(new_n326), .A3(new_n722), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT115), .ZN(new_n837));
  INV_X1    g651(.A(new_n313), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n759), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n730), .ZN(new_n840));
  OR2_X1    g654(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n843));
  NAND2_X1  g657(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n837), .A2(new_n840), .A3(new_n844), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n762), .A2(new_n722), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n605), .A2(new_n313), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n676), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n691), .A2(new_n688), .A3(new_n618), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n847), .A2(new_n784), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n843), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT117), .A4(new_n851), .ZN(new_n855));
  INV_X1    g669(.A(new_n702), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n437), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n762), .B(new_n840), .C1(new_n776), .C2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n854), .A2(KEYINPUT51), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n747), .A2(new_n605), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n847), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT48), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n312), .B(G953), .C1(new_n849), .C2(new_n632), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n847), .A2(KEYINPUT48), .A3(new_n860), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n840), .A2(new_n715), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n858), .A2(new_n843), .A3(new_n845), .A4(new_n851), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n859), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n859), .A2(KEYINPUT118), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n835), .A2(new_n875), .B1(G952), .B2(G953), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n856), .A2(KEYINPUT49), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n856), .A2(KEYINPUT49), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n757), .A2(new_n605), .A3(new_n325), .A4(new_n437), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n667), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n876), .B1(new_n676), .B2(new_n881), .ZN(G75));
  AOI21_X1  g696(.A(new_n245), .B1(new_n819), .B2(new_n830), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(G210), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n376), .A2(new_n408), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n431), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n884), .B1(new_n883), .B2(G210), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n260), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n883), .B2(G210), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n889), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n892), .A2(new_n896), .ZN(G51));
  XNOR2_X1  g711(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n767), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n781), .B1(new_n819), .B2(new_n830), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n833), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n495), .B2(new_n486), .ZN(new_n902));
  INV_X1    g716(.A(new_n883), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(new_n766), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n893), .B1(new_n902), .B2(new_n904), .ZN(G54));
  NAND2_X1  g719(.A1(KEYINPUT58), .A2(G475), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n318), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .A4(new_n306), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n907), .A2(new_n894), .A3(new_n908), .ZN(G60));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n629), .B1(new_n835), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n629), .B(new_n912), .C1(new_n833), .C2(new_n900), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n894), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(G63));
  XNOR2_X1  g730(.A(new_n595), .B(KEYINPUT122), .ZN(new_n917));
  XNOR2_X1  g731(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n917), .B(new_n918), .Z(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n821), .B2(new_n804), .ZN(new_n920));
  AND4_X1   g734(.A1(new_n816), .A2(new_n796), .A3(new_n804), .A4(new_n829), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n893), .B1(new_n922), .B2(new_n602), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT61), .B1(new_n923), .B2(KEYINPUT123), .ZN(new_n924));
  INV_X1    g738(.A(new_n919), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n819), .B2(new_n830), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n894), .B1(new_n926), .B2(new_n603), .ZN(new_n927));
  INV_X1    g741(.A(new_n651), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n928), .B(new_n925), .C1(new_n819), .C2(new_n830), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT124), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n651), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n923), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n924), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  OAI211_X1 g749(.A(KEYINPUT123), .B(new_n894), .C1(new_n926), .C2(new_n603), .ZN(new_n936));
  AOI22_X1  g750(.A1(new_n930), .A2(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n934), .A2(new_n937), .ZN(G66));
  INV_X1    g752(.A(new_n315), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n260), .B1(new_n939), .B2(G224), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n783), .A2(new_n732), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n820), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n943), .B2(new_n260), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n430), .B(new_n369), .C1(G898), .C2(new_n260), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n944), .B(new_n945), .Z(G69));
  AND3_X1   g760(.A1(new_n664), .A2(new_n694), .A3(new_n735), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n685), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(KEYINPUT62), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n632), .B1(new_n640), .B2(new_n321), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n683), .A3(new_n737), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n566), .A3(new_n605), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n779), .A2(new_n774), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n948), .A2(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n260), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n513), .B1(new_n518), .B2(KEYINPUT30), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n301), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n755), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n752), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT126), .Z(new_n965));
  NAND4_X1  g779(.A1(new_n773), .A2(new_n860), .A3(new_n433), .A4(new_n723), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n779), .A2(new_n774), .A3(new_n947), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n260), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n954), .B2(new_n955), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT125), .B1(new_n972), .B2(new_n960), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n962), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n962), .A2(new_n973), .A3(new_n977), .A4(new_n971), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n956), .B2(new_n943), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n671), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n819), .A2(new_n825), .ZN(new_n984));
  INV_X1    g798(.A(new_n981), .ZN(new_n985));
  INV_X1    g799(.A(new_n563), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n525), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n894), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n985), .B1(new_n968), .B2(new_n942), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n519), .A2(new_n520), .A3(new_n529), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(G57));
endmodule


