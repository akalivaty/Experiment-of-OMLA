//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT67), .B(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(KEYINPUT3), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT68), .B(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(new_n464), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n463), .B(G2104), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  INV_X1    g050(.A(G113), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n464), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n479), .B2(new_n461), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n483), .B1(new_n486), .B2(G2104), .ZN(new_n487));
  AOI211_X1 g062(.A(KEYINPUT69), .B(new_n464), .C1(new_n484), .C2(new_n485), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT70), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT67), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G112), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n489), .A2(new_n461), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G124), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G162));
  NAND2_X1  g079(.A1(G126), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT4), .A4(G138), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n467), .A2(new_n472), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n470), .A2(G2104), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n482), .A2(new_n509), .A3(G138), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n510), .B2(new_n498), .ZN(new_n511));
  OAI21_X1  g086(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n512));
  INV_X1    g087(.A(G114), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(G2105), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G164));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n518), .B2(new_n519), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G88), .B1(G50), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n525), .B(KEYINPUT71), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(G50), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(new_n521), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n527), .A2(new_n526), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n528), .A2(new_n535), .ZN(G166));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT73), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT7), .Z(new_n539));
  AOI22_X1  g114(.A1(new_n520), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n540));
  INV_X1    g115(.A(new_n521), .ZN(new_n541));
  INV_X1    g116(.A(new_n524), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT72), .B(G51), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n539), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n522), .A2(G90), .B1(G52), .B2(new_n524), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT74), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n526), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT75), .B(G43), .Z(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n532), .B1(new_n542), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n526), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n524), .A2(G53), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT9), .Z(new_n564));
  AOI22_X1  g139(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n526), .B1(new_n532), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  OAI21_X1  g146(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n522), .A2(new_n575), .A3(G87), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT76), .B1(new_n532), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n524), .A2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n524), .A2(G48), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n532), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n526), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT78), .Z(G305));
  AOI22_X1  g163(.A1(new_n522), .A2(G85), .B1(G47), .B2(new_n524), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n541), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n526), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n594), .B2(new_n593), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n590), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n520), .A2(new_n521), .A3(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT81), .Z(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n526), .B1(new_n603), .B2(new_n604), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n542), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n524), .A2(KEYINPUT82), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n605), .A2(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n599), .B(KEYINPUT81), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n602), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n598), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n598), .B1(new_n614), .B2(G868), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n568), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(G868), .B2(new_n568), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n614), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI22_X1  g198(.A1(new_n623), .A2(KEYINPUT84), .B1(G868), .B2(new_n557), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(KEYINPUT84), .B2(new_n623), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT85), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n478), .A2(new_n474), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2100), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n490), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n501), .A2(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n461), .C2(G111), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(G156));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n650), .ZN(G401));
  NOR2_X1   g229(.A1(G2072), .A2(G2078), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n442), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n663), .B(new_n660), .C1(new_n656), .C2(new_n659), .ZN(new_n664));
  INV_X1    g239(.A(new_n656), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n665), .A2(new_n660), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n677), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  AOI211_X1 g256(.A(new_n679), .B(new_n681), .C1(new_n674), .C2(new_n678), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XOR2_X1   g258(.A(new_n682), .B(new_n683), .Z(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G20), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT23), .Z(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G299), .B2(G16), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G1956), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n697), .A2(G35), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n503), .B2(G29), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G2090), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n696), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n702), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n705), .B(KEYINPUT95), .C1(KEYINPUT94), .C2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(G28), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n697), .B1(new_n708), .B2(G28), .ZN(new_n710));
  AND2_X1   g285(.A1(KEYINPUT31), .A2(G11), .ZN(new_n711));
  NOR2_X1   g286(.A1(KEYINPUT31), .A2(G11), .ZN(new_n712));
  OAI22_X1  g287(.A1(new_n709), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n557), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G19), .ZN(new_n715));
  INV_X1    g290(.A(G1341), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G171), .A2(new_n691), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G5), .B2(new_n691), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n717), .B1(new_n716), .B2(new_n715), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT25), .Z(new_n724));
  AOI22_X1  g299(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n461), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G139), .B2(new_n490), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n697), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n697), .A2(G33), .ZN(new_n729));
  OAI21_X1  g304(.A(G2072), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n728), .A2(G2072), .A3(new_n729), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n722), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G168), .A2(new_n691), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n691), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G27), .A2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G164), .B2(G29), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G2078), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n697), .B1(new_n740), .B2(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n740), .B2(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G160), .B2(G29), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G2084), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G2084), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n736), .A2(new_n739), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n721), .A2(new_n732), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n490), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n501), .A2(G129), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(G105), .B2(new_n474), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n748), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(new_n697), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n697), .B2(G32), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n738), .A2(G2078), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n762), .B1(new_n635), .B2(new_n697), .C1(new_n734), .C2(new_n735), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G4), .A2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n602), .A2(new_n611), .A3(new_n613), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n691), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G1348), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n697), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT28), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n490), .A2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n501), .A2(G128), .ZN(new_n773));
  OAI221_X1 g348(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n461), .C2(G116), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n771), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G2067), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n769), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n747), .A2(new_n760), .A3(new_n764), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n701), .A2(G2090), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n706), .A2(KEYINPUT94), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n704), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n707), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(G6), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G305), .B2(new_n691), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT91), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n789), .B(new_n790), .Z(new_n791));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n792));
  NAND2_X1  g367(.A1(G166), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G16), .B2(G22), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(G1971), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(G1971), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n797), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n799), .A2(new_n795), .A3(KEYINPUT92), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n691), .A2(G23), .ZN(new_n802));
  INV_X1    g377(.A(G288), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n691), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT33), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1976), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT34), .B1(new_n791), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n789), .B(new_n790), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n809), .A2(new_n810), .A3(new_n801), .A4(new_n806), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n697), .A2(G25), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n501), .A2(G119), .ZN(new_n813));
  OAI221_X1 g388(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n461), .C2(G107), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n490), .A2(G131), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(new_n697), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XOR2_X1   g395(.A(new_n819), .B(new_n820), .Z(new_n821));
  NOR2_X1   g396(.A1(G16), .A2(G24), .ZN(new_n822));
  INV_X1    g397(.A(G290), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT90), .B(G1986), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n808), .A2(new_n811), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n808), .A2(new_n811), .A3(new_n830), .A4(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n786), .A2(new_n832), .ZN(G311));
  AND3_X1   g408(.A1(new_n786), .A2(new_n832), .A3(KEYINPUT96), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT96), .B1(new_n786), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n541), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n526), .B1(new_n839), .B2(KEYINPUT97), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(KEYINPUT97), .B2(new_n839), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n522), .A2(G93), .B1(G55), .B2(new_n524), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT99), .B(G860), .Z(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n614), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  INV_X1    g424(.A(new_n557), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n843), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT98), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n845), .B1(new_n852), .B2(new_n853), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n847), .B1(new_n855), .B2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n503), .B(new_n635), .ZN(new_n858));
  XNOR2_X1  g433(.A(G160), .B(KEYINPUT100), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n817), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n629), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n817), .B(KEYINPUT101), .ZN(new_n864));
  INV_X1    g439(.A(new_n629), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n490), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n501), .A2(G130), .ZN(new_n868));
  OAI221_X1 g443(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n461), .C2(G118), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n863), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n863), .B2(new_n866), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n775), .B(G164), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(new_n755), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n755), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n727), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n727), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n875), .A2(new_n876), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT102), .B1(new_n886), .B2(new_n874), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n875), .B2(new_n884), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n874), .A3(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n860), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT104), .B(G37), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n885), .A2(new_n887), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n860), .B1(new_n886), .B2(new_n874), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n893), .A2(new_n898), .A3(KEYINPUT40), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT40), .B1(new_n893), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(G395));
  XNOR2_X1  g476(.A(G305), .B(G288), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(G303), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n622), .B(new_n851), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n614), .A2(new_n568), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n767), .A2(G299), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT105), .B1(new_n912), .B2(KEYINPUT41), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n917), .B2(KEYINPUT105), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n911), .B1(new_n918), .B2(new_n907), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n906), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n906), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(G868), .B2(new_n844), .ZN(G295));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n844), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  XNOR2_X1  g503(.A(G301), .B(G286), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(new_n851), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n851), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n917), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(KEYINPUT108), .A3(new_n851), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n930), .A2(new_n912), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n934), .A2(KEYINPUT109), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n917), .A2(new_n941), .A3(new_n933), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n904), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n939), .A2(new_n932), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n930), .B1(new_n936), .B2(new_n937), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n904), .B(new_n947), .C1(new_n918), .C2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n945), .A2(new_n946), .A3(new_n894), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n894), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n904), .B1(new_n940), .B2(new_n942), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT110), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n928), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G37), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n947), .B1(new_n918), .B2(new_n948), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n944), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT43), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT44), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n928), .B1(new_n956), .B2(new_n958), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(G397));
  OR2_X1    g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT112), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(G1986), .B2(G290), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n817), .B(new_n820), .Z(new_n969));
  XNOR2_X1  g544(.A(new_n775), .B(new_n777), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n755), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n506), .A2(new_n505), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n487), .B2(new_n488), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n461), .A2(new_n478), .A3(G138), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n514), .B1(new_n978), .B2(new_n508), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n473), .A2(new_n480), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(KEYINPUT111), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(KEYINPUT111), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n975), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT115), .B(G8), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(G286), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT119), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n507), .B2(new_n516), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT114), .B(new_n994), .C1(new_n507), .C2(new_n516), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G2084), .ZN(new_n1000));
  INV_X1    g575(.A(new_n462), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n487), .B2(new_n488), .ZN(new_n1002));
  INV_X1    g577(.A(new_n475), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n482), .A2(new_n509), .A3(G125), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n476), .B2(new_n464), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n1005), .B2(new_n498), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1006), .A3(G40), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n507), .B2(new_n516), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(KEYINPUT50), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n999), .A2(new_n1000), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n1008), .C1(new_n507), .C2(new_n516), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n983), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n735), .B1(new_n1013), .B2(new_n981), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n993), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT51), .B1(new_n992), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(KEYINPUT120), .A3(new_n990), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n991), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT120), .B1(new_n1017), .B2(new_n990), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n991), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT118), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n999), .A2(new_n1010), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1013), .A2(new_n981), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2078), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n720), .A2(new_n1027), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G2078), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1007), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n980), .A2(new_n1034), .A3(KEYINPUT45), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT113), .B1(new_n1009), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1032), .B(new_n1033), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1029), .ZN(new_n1039));
  AOI21_X1  g614(.A(G301), .B1(new_n1031), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n528), .A2(new_n535), .A3(G8), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1034), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1009), .A2(KEYINPUT113), .A3(new_n1036), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1971), .B1(new_n1046), .B2(new_n1033), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n999), .A2(new_n1048), .A3(new_n1010), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1043), .B(G8), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n983), .A2(new_n980), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n574), .A2(new_n579), .A3(G1976), .A4(new_n580), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1052), .A2(new_n990), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  OAI21_X1  g631(.A(G1981), .B1(new_n584), .B2(new_n586), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n584), .A2(new_n586), .A3(G1981), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1981), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n587), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(KEYINPUT49), .A3(new_n1057), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(new_n990), .A3(new_n1063), .A4(new_n1053), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1053), .A2(new_n990), .A3(new_n1054), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1055), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1033), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1068));
  INV_X1    g643(.A(G1971), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1071), .A2(new_n983), .A3(new_n995), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1048), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n989), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1050), .B(new_n1067), .C1(new_n1074), .C2(new_n1043), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1026), .A2(new_n1040), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1053), .A2(new_n990), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1064), .A2(new_n1051), .A3(new_n803), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(new_n1062), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1067), .B(KEYINPUT116), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1050), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(G286), .B(new_n989), .C1(new_n1011), .C2(new_n1014), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(KEYINPUT63), .ZN(new_n1086));
  OAI21_X1  g661(.A(G8), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1043), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND4_X1   g664(.A1(new_n1050), .A2(new_n1082), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT63), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1084), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1013), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1010), .A2(new_n995), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT117), .B(G1956), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n568), .B(KEYINPUT57), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1095), .A2(new_n1100), .A3(new_n1098), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1348), .B1(new_n999), .B2(new_n1010), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1053), .A2(G2067), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n614), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1102), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n614), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1093), .A2(new_n971), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1053), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n850), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1111), .B1(new_n1115), .B2(KEYINPUT59), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1115), .A2(KEYINPUT59), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1109), .A2(new_n767), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1110), .B1(new_n1118), .B2(new_n1107), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1102), .A2(KEYINPUT61), .A3(new_n1103), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT61), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1108), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1009), .A2(new_n1036), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT122), .B(G2078), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1033), .A2(KEYINPUT53), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1961), .B1(new_n999), .B2(new_n1010), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(KEYINPUT121), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n1093), .B2(new_n1032), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1131), .B(G1961), .C1(new_n999), .C2(new_n1010), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1040), .B1(new_n1133), .B2(G301), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT123), .B1(new_n1134), .B2(KEYINPUT54), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1027), .A2(new_n720), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1131), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1128), .A2(KEYINPUT121), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n1039), .A3(new_n1140), .A4(new_n1127), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1136), .B(new_n1137), .C1(new_n1142), .C2(new_n1040), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1031), .A2(G301), .A3(new_n1039), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1144), .A2(KEYINPUT54), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(G171), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1075), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1135), .A2(new_n1143), .A3(new_n1147), .A4(new_n1025), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1124), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1147), .A2(new_n1025), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(KEYINPUT124), .A3(new_n1143), .A4(new_n1135), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1092), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1078), .B1(new_n1153), .B2(KEYINPUT125), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1155), .B(new_n1092), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n988), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n987), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n970), .B2(new_n756), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT126), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n987), .A2(new_n971), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT46), .Z(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT47), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n967), .A2(KEYINPUT48), .A3(new_n987), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n974), .B2(new_n1158), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT48), .B1(new_n967), .B2(new_n987), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n818), .A2(new_n820), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n973), .A2(new_n1169), .B1(G2067), .B2(new_n775), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1170), .A2(new_n987), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1164), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1157), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g748(.A(G319), .ZN(new_n1175));
  NOR3_X1   g749(.A1(G401), .A2(G227), .A3(new_n1175), .ZN(new_n1176));
  XOR2_X1   g750(.A(new_n1176), .B(KEYINPUT127), .Z(new_n1177));
  NAND2_X1  g751(.A1(new_n1177), .A2(new_n689), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n893), .B2(new_n898), .ZN(new_n1179));
  OR2_X1    g753(.A1(new_n962), .A2(new_n963), .ZN(new_n1180));
  AND2_X1   g754(.A1(new_n1179), .A2(new_n1180), .ZN(G308));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(G225));
endmodule


