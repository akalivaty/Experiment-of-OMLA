//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1318, new_n1319, new_n1320, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1388, new_n1389,
    new_n1390;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AND2_X1   g0014(.A1(KEYINPUT65), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(KEYINPUT65), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n204), .A2(new_n205), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n214), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n223), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n236), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(new_n217), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n251), .A2(new_n252), .B1(new_n209), .B2(G68), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT72), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n255), .B1(new_n209), .B2(G68), .C1(new_n251), .C2(new_n252), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n254), .B(new_n256), .C1(new_n221), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT73), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n218), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n259), .B2(new_n262), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT11), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n259), .A2(new_n262), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT11), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n269), .A3(new_n263), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n271), .A2(new_n209), .A3(G1), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n203), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT12), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n272), .A2(new_n262), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n203), .B1(new_n208), .B2(G20), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n266), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  AND2_X1   g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  AOI21_X1  g0085(.A(G1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(G274), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n286), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(G238), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G226), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n292), .A2(new_n296), .A3(G226), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NOR2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n238), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n280), .B(new_n291), .C1(new_n304), .C2(new_n283), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n283), .B1(new_n298), .B2(new_n303), .ZN(new_n306));
  INV_X1    g0106(.A(new_n291), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT13), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT14), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n310), .A3(G169), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(G179), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n309), .B2(G169), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n279), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n309), .A2(G200), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n305), .A2(G190), .A3(new_n308), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n279), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n283), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G226), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n287), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n292), .A2(G222), .A3(new_n293), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n292), .A2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n326), .B1(new_n252), .B2(new_n292), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n329), .B2(new_n289), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(G179), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  INV_X1    g0133(.A(G150), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n251), .A2(new_n333), .B1(new_n334), .B2(new_n258), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n209), .B1(new_n220), .B2(new_n221), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n262), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n221), .B1(new_n208), .B2(G20), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n276), .A2(new_n338), .B1(new_n221), .B2(new_n272), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n330), .A2(G169), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n332), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT9), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n337), .A2(new_n339), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n344), .A2(new_n345), .B1(new_n330), .B2(G190), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(KEYINPUT9), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n331), .A2(G200), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(KEYINPUT10), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT10), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n340), .A2(KEYINPUT9), .B1(new_n331), .B2(G200), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n346), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n343), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n292), .A2(G232), .A3(new_n293), .ZN(new_n355));
  INV_X1    g0155(.A(G107), .ZN(new_n356));
  INV_X1    g0156(.A(G238), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n355), .B1(new_n356), .B2(new_n292), .C1(new_n327), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n289), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n288), .B1(G244), .B2(new_n290), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n262), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT69), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(G33), .A3(new_n217), .ZN(new_n368));
  INV_X1    g0168(.A(new_n333), .ZN(new_n369));
  OR2_X1    g0169(.A1(KEYINPUT65), .A2(G20), .ZN(new_n370));
  NAND2_X1  g0170(.A1(KEYINPUT65), .A2(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n369), .A2(new_n257), .B1(new_n372), .B2(G77), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n364), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n276), .B(G77), .C1(G1), .C2(new_n209), .ZN(new_n375));
  INV_X1    g0175(.A(new_n272), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n376), .A2(KEYINPUT70), .A3(G77), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT70), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n272), .B2(new_n252), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n363), .B1(G179), .B2(new_n361), .C1(new_n374), .C2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n374), .A2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n361), .A2(G200), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n361), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n354), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n333), .B1(new_n208), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n276), .B1(new_n272), .B2(new_n333), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT7), .B1(new_n292), .B2(G20), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n217), .A2(new_n301), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n393), .A3(G68), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT74), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n202), .A2(new_n203), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(G20), .C1(new_n220), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n257), .A2(G159), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n397), .B1(new_n402), .B2(G20), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n364), .B1(new_n396), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n220), .B2(new_n398), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT74), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n400), .A3(new_n399), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT7), .B1(new_n372), .B2(new_n292), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n301), .A2(new_n392), .A3(new_n209), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G68), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n406), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n390), .B1(new_n405), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n328), .A2(new_n293), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n324), .A2(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n299), .C2(new_n300), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n289), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n290), .A2(G232), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(G179), .A3(new_n287), .A4(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n287), .B1(new_n323), .B2(new_n238), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n283), .B1(new_n418), .B2(new_n419), .ZN(new_n425));
  OAI21_X1  g0225(.A(G169), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n423), .A2(KEYINPUT75), .A3(new_n426), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT18), .B1(new_n415), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n424), .A2(new_n425), .ZN(new_n433));
  XOR2_X1   g0233(.A(KEYINPUT76), .B(G190), .Z(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G200), .B2(new_n433), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n430), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT75), .B1(new_n423), .B2(new_n426), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT16), .B1(new_n404), .B2(new_n412), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n262), .B1(new_n409), .B2(new_n395), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n389), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n436), .B(new_n389), .C1(new_n441), .C2(new_n442), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n432), .A2(new_n437), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT77), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n449), .A2(KEYINPUT77), .ZN(new_n451));
  AND4_X1   g0251(.A1(new_n321), .A2(new_n387), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n376), .A2(G116), .ZN(new_n454));
  AOI211_X1 g0254(.A(new_n262), .B(new_n272), .C1(new_n208), .C2(G33), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G116), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n262), .B1(new_n209), .B2(G116), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT86), .ZN(new_n458));
  INV_X1    g0258(.A(G33), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G97), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n372), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n217), .A2(KEYINPUT86), .A3(new_n460), .A4(new_n461), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n457), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT20), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  AOI211_X1 g0267(.A(new_n467), .B(new_n457), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n456), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g0269(.A1(KEYINPUT3), .A2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT3), .A2(G33), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT85), .A2(G303), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT85), .A2(G303), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G257), .B(new_n293), .C1(new_n299), .C2(new_n300), .ZN(new_n475));
  OAI211_X1 g0275(.A(G264), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n289), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n208), .B(G45), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G41), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n283), .B(G270), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n285), .A2(G1), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT79), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(G41), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G274), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n281), .B2(new_n282), .ZN(new_n489));
  INV_X1    g0289(.A(new_n481), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n483), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n478), .A2(new_n482), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n469), .A2(G169), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n492), .A2(new_n434), .ZN(new_n496));
  INV_X1    g0296(.A(G200), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n491), .A2(new_n482), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n478), .ZN(new_n499));
  OR3_X1    g0299(.A1(new_n469), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n477), .A2(new_n289), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n482), .ZN(new_n502));
  OAI211_X1 g0302(.A(KEYINPUT21), .B(G169), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n478), .A2(G179), .A3(new_n482), .A4(new_n491), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT87), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(new_n506), .A3(new_n469), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(new_n469), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n495), .B(new_n500), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT84), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(new_n293), .C1(new_n299), .C2(new_n300), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n461), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n289), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n283), .B(G257), .C1(new_n479), .C2(new_n481), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n491), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n520), .A3(G190), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT80), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n517), .A2(new_n520), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT6), .ZN(new_n526));
  AND2_X1   g0326(.A1(G97), .A2(G107), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT6), .A2(G97), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT78), .B1(new_n530), .B2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT78), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(new_n356), .A3(KEYINPUT6), .A4(G97), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n372), .B1(G77), .B2(new_n257), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n410), .A2(G107), .A3(new_n411), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n364), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n272), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n276), .B1(G1), .B2(new_n459), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(new_n538), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n517), .A2(new_n520), .A3(KEYINPUT80), .A4(G190), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n523), .A2(new_n525), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n519), .B1(new_n289), .B2(new_n516), .ZN(new_n545));
  INV_X1    g0345(.A(G179), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT81), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND4_X1   g0347(.A1(KEYINPUT81), .A2(new_n517), .A3(new_n546), .A4(new_n520), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n545), .A2(G169), .B1(new_n537), .B2(new_n541), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G87), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n528), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n554), .A2(new_n459), .A3(new_n538), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(new_n372), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n370), .A2(G33), .A3(G97), .A4(new_n371), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n554), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n217), .A2(new_n292), .A3(G68), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n262), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n455), .A2(new_n367), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n365), .B(KEYINPUT69), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n272), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT83), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n208), .A2(G45), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G250), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n289), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n283), .A2(KEYINPUT82), .A3(G250), .A4(new_n568), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n570), .A2(new_n571), .B1(new_n489), .B2(new_n484), .ZN(new_n572));
  OAI211_X1 g0372(.A(G244), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n573));
  OAI211_X1 g0373(.A(G238), .B(new_n293), .C1(new_n299), .C2(new_n300), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G116), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n289), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G169), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n572), .A2(G179), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n560), .A2(new_n262), .B1(new_n563), .B2(new_n272), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n562), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n566), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n578), .A2(G200), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n455), .A2(G87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n572), .A2(G190), .A3(new_n577), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n586), .A2(new_n582), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n510), .B1(new_n551), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G257), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n592));
  OAI211_X1 g0392(.A(G250), .B(new_n293), .C1(new_n299), .C2(new_n300), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G294), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n289), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n283), .B(G264), .C1(new_n479), .C2(new_n481), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n491), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT88), .ZN(new_n599));
  INV_X1    g0399(.A(new_n597), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n289), .B2(new_n595), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT88), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n491), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n603), .A3(new_n384), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n596), .A2(KEYINPUT89), .A3(new_n597), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT89), .B1(new_n596), .B2(new_n597), .ZN(new_n606));
  INV_X1    g0406(.A(new_n491), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n604), .B1(new_n608), .B2(G200), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT25), .B1(new_n272), .B2(new_n356), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n272), .A2(KEYINPUT25), .A3(new_n356), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n455), .A2(G107), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT23), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n356), .C1(new_n215), .C2(new_n216), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n575), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n209), .ZN(new_n618));
  NAND2_X1  g0418(.A1(KEYINPUT23), .A2(G107), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n217), .A2(new_n292), .A3(G87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT22), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT22), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n217), .A2(new_n292), .A3(new_n623), .A4(G87), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT24), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n614), .B1(new_n627), .B2(new_n262), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n609), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n625), .A2(new_n626), .ZN(new_n630));
  AOI211_X1 g0430(.A(KEYINPUT24), .B(new_n620), .C1(new_n622), .C2(new_n624), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n262), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n613), .ZN(new_n633));
  NOR4_X1   g0433(.A1(new_n605), .A2(new_n606), .A3(new_n546), .A4(new_n607), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n362), .B1(new_n599), .B2(new_n603), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(KEYINPUT83), .A2(new_n565), .B1(new_n579), .B2(new_n580), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n586), .A2(new_n588), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n582), .A2(new_n587), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n638), .A2(new_n584), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n550), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n517), .A2(new_n520), .A3(new_n546), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT81), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n545), .A2(KEYINPUT81), .A3(new_n546), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n641), .A2(KEYINPUT84), .A3(new_n648), .A4(new_n544), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n591), .A2(new_n637), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n453), .A2(new_n509), .A3(new_n650), .ZN(G372));
  INV_X1    g0451(.A(new_n427), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT18), .B1(new_n415), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n443), .A2(new_n444), .A3(new_n427), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n437), .A2(new_n448), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n320), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n315), .A2(new_n381), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n349), .A2(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n352), .A2(new_n351), .A3(new_n346), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n343), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT91), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT91), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n666), .B(new_n343), .C1(new_n659), .C2(new_n663), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n580), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n362), .B1(new_n572), .B2(new_n577), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n565), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n550), .B1(new_n645), .B2(new_n646), .ZN(new_n673));
  XNOR2_X1  g0473(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n641), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n589), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n648), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n672), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n493), .A2(new_n494), .B1(new_n469), .B2(new_n505), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n636), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n523), .A2(new_n542), .A3(new_n525), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n683), .A2(new_n543), .B1(new_n647), .B2(new_n642), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n678), .B1(new_n609), .B2(new_n628), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n452), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n668), .A2(new_n688), .ZN(G369));
  NAND2_X1  g0489(.A1(new_n505), .A2(new_n469), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n495), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n271), .A2(G1), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n217), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n217), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n694), .A2(G213), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT92), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(new_n469), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n691), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n509), .B2(new_n700), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n629), .A2(new_n636), .ZN(new_n704));
  INV_X1    g0504(.A(new_n699), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n628), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n704), .A2(new_n706), .B1(new_n636), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n636), .A2(new_n699), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n690), .A2(KEYINPUT87), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n505), .A2(new_n506), .A3(new_n469), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n699), .B1(new_n712), .B2(new_n495), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n709), .B1(new_n713), .B2(new_n637), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n212), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n222), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n208), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n553), .A2(G116), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n722), .B2(new_n721), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  INV_X1    g0525(.A(KEYINPUT94), .ZN(new_n726));
  INV_X1    g0526(.A(new_n504), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n596), .A2(new_n597), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT89), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n572), .A2(new_n577), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n727), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n545), .A2(KEYINPUT30), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n726), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n734), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n605), .A2(new_n606), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n504), .A2(new_n578), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT94), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(G179), .B1(new_n498), .B2(new_n478), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n524), .A3(new_n578), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT96), .B1(new_n608), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n730), .A2(new_n731), .A3(new_n491), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n492), .A2(new_n578), .A3(new_n546), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT96), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n524), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n737), .A2(new_n545), .A3(new_n738), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n749), .A2(KEYINPUT95), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT95), .B1(new_n749), .B2(new_n750), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n740), .B(new_n748), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT97), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n750), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n749), .A2(KEYINPUT95), .A3(new_n750), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n735), .A2(new_n739), .B1(new_n743), .B2(new_n747), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT97), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT31), .B1(new_n763), .B2(new_n699), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n740), .B(new_n755), .C1(new_n608), .C2(new_n742), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n705), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n509), .A2(new_n699), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n650), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(G330), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n674), .B1(new_n590), .B2(new_n648), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n671), .A2(new_n589), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n673), .A3(KEYINPUT26), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n672), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n495), .B1(new_n507), .B2(new_n508), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n634), .A2(new_n635), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n628), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n684), .B(new_n685), .C1(new_n776), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n699), .B1(new_n680), .B2(new_n686), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(KEYINPUT29), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n771), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n725), .B1(new_n785), .B2(G1), .ZN(G364));
  NOR2_X1   g0586(.A1(new_n372), .A2(new_n271), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G45), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n719), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n703), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(G330), .B2(new_n702), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n716), .A2(new_n301), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G355), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G116), .B2(new_n212), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n716), .A2(new_n292), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n222), .B2(new_n285), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n249), .A2(G45), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n218), .B1(G20), .B2(new_n362), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n790), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n217), .A2(new_n546), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(KEYINPUT98), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n434), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n808), .A2(KEYINPUT98), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G322), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n810), .A2(new_n384), .A3(new_n812), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G311), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n497), .A2(G179), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n819), .A2(G20), .A3(G190), .ZN(new_n820));
  INV_X1    g0620(.A(G303), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n301), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G179), .A2(G200), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n217), .B1(G190), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G294), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n372), .A2(new_n384), .A3(new_n819), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n824), .A2(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n372), .A2(new_n384), .A3(new_n823), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n822), .B(new_n828), .C1(G329), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n808), .A2(G200), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n434), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(G190), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT33), .B(G317), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n833), .A2(G326), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n815), .A2(new_n818), .A3(new_n831), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G159), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n829), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n834), .A2(G68), .B1(new_n840), .B2(KEYINPUT32), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n824), .A2(new_n538), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n826), .A2(new_n356), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n292), .B1(new_n820), .B2(new_n552), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT32), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n833), .A2(G50), .B1(new_n846), .B2(new_n839), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n841), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n202), .A2(new_n813), .B1(new_n816), .B2(new_n252), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n837), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n807), .B1(new_n850), .B2(new_n804), .ZN(new_n851));
  INV_X1    g0651(.A(new_n803), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n702), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n792), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NOR2_X1   g0655(.A1(new_n381), .A2(new_n699), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n385), .B1(new_n705), .B2(new_n382), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n381), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n782), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n590), .A2(new_n648), .A3(new_n674), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT26), .B1(new_n773), .B2(new_n673), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n671), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n705), .B(new_n858), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n782), .A2(KEYINPUT101), .A3(new_n858), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n859), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(G330), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n753), .A2(KEYINPUT97), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n699), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n766), .ZN(new_n873));
  INV_X1    g0673(.A(new_n770), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT102), .ZN(new_n876));
  OR3_X1    g0676(.A1(new_n868), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n868), .B2(new_n875), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n790), .B1(new_n868), .B2(new_n875), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n804), .A2(new_n801), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n789), .B1(new_n252), .B2(new_n881), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n292), .B1(new_n221), .B2(new_n820), .C1(new_n826), .C2(new_n203), .ZN(new_n883));
  INV_X1    g0683(.A(G132), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n824), .A2(new_n202), .B1(new_n829), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(G137), .A2(new_n833), .B1(new_n834), .B2(G150), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n838), .B2(new_n816), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(G143), .B2(new_n814), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT100), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT34), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n883), .B(new_n885), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n817), .A2(G116), .B1(G283), .B2(new_n834), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT99), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n826), .A2(new_n552), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n301), .B1(new_n356), .B2(new_n820), .C1(new_n824), .C2(new_n538), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n896), .B(new_n897), .C1(G311), .C2(new_n830), .ZN(new_n898));
  INV_X1    g0698(.A(new_n833), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n898), .B1(new_n825), .B2(new_n813), .C1(new_n821), .C2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT99), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n893), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n891), .A2(new_n892), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n804), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n882), .B1(new_n802), .B2(new_n858), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n880), .A2(new_n905), .ZN(G384));
  OR2_X1    g0706(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n907), .A2(G116), .A3(new_n219), .A4(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT36), .Z(new_n910));
  OAI211_X1 g0710(.A(new_n222), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n221), .A2(G68), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n208), .B(G13), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n856), .B1(new_n866), .B2(new_n867), .ZN(new_n915));
  INV_X1    g0715(.A(new_n278), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n268), .A2(new_n263), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(KEYINPUT11), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n918), .A2(new_n270), .A3(new_n318), .A4(new_n317), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n279), .A2(new_n699), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n315), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n279), .B(new_n699), .C1(new_n313), .C2(new_n314), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n391), .A2(new_n393), .A3(G68), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n406), .B1(new_n409), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n390), .B1(new_n405), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n446), .B1(new_n928), .B2(new_n652), .ZN(new_n929));
  INV_X1    g0729(.A(new_n697), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT37), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT37), .B1(new_n440), .B2(new_n443), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n443), .A2(new_n697), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n446), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n449), .A2(new_n931), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT38), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n925), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n655), .A2(new_n930), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n316), .A2(new_n705), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n934), .B(new_n446), .C1(new_n415), .C2(new_n652), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT37), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n653), .A2(new_n437), .A3(new_n654), .A4(new_n448), .ZN(new_n949));
  INV_X1    g0749(.A(new_n934), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n948), .A2(new_n935), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n940), .B(new_n946), .C1(new_n951), .C2(KEYINPUT38), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT103), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT38), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n949), .A2(new_n950), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n446), .B1(new_n415), .B2(new_n930), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(KEYINPUT37), .A2(new_n947), .B1(new_n958), .B2(new_n933), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n955), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT103), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(new_n946), .A4(new_n940), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT38), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT39), .B1(new_n963), .B2(new_n938), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT104), .B1(new_n954), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT104), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n953), .A2(new_n967), .A3(new_n964), .A4(new_n962), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n945), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n944), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n783), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n452), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n668), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n970), .B(new_n973), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n960), .A2(new_n940), .ZN(new_n975));
  INV_X1    g0775(.A(new_n858), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n921), .B2(new_n922), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n767), .B1(new_n870), .B2(new_n871), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n591), .A2(new_n637), .A3(new_n649), .ZN(new_n979));
  INV_X1    g0779(.A(new_n769), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n975), .B(new_n977), .C1(new_n982), .C2(new_n764), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n923), .A2(new_n858), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n763), .A2(new_n767), .B1(new_n979), .B2(new_n980), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(new_n873), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT40), .B1(new_n939), .B2(new_n940), .ZN(new_n987));
  AOI22_X1  g0787(.A1(KEYINPUT40), .A2(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n982), .A2(new_n764), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n453), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n983), .A2(KEYINPUT40), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n873), .A2(new_n985), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n977), .A3(new_n987), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(new_n452), .A3(new_n992), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n990), .A2(new_n995), .A3(G330), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n974), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n208), .B2(new_n787), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n974), .A2(new_n996), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n914), .B1(new_n998), .B2(new_n999), .ZN(G367));
  NAND2_X1  g0800(.A1(new_n236), .A2(new_n796), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n806), .B1(new_n367), .B2(new_n716), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n789), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n705), .A2(new_n640), .ZN(new_n1004));
  MUX2_X1   g0804(.A(new_n773), .B(new_n672), .S(new_n1004), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n826), .A2(new_n252), .ZN(new_n1006));
  INV_X1    g0806(.A(G137), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n292), .B1(new_n202), .B2(new_n820), .C1(new_n829), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n824), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1006), .B(new_n1008), .C1(G68), .C2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G143), .A2(new_n833), .B1(new_n834), .B2(G159), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n221), .B2(new_n816), .C1(new_n334), .C2(new_n813), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n826), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(G97), .ZN(new_n1015));
  INV_X1    g0815(.A(G317), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT46), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n820), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT112), .B1(new_n1018), .B2(G116), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1015), .B1(new_n1016), .B2(new_n829), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n292), .B1(new_n1019), .B2(new_n1017), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n834), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1021), .B1(new_n1022), .B2(new_n825), .ZN(new_n1023));
  XOR2_X1   g0823(.A(KEYINPUT111), .B(G311), .Z(new_n1024));
  AOI211_X1 g0824(.A(new_n1020), .B(new_n1023), .C1(new_n833), .C2(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n816), .A2(new_n827), .B1(new_n356), .B2(new_n824), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT110), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n472), .A2(new_n473), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1025), .B(new_n1028), .C1(new_n1029), .C2(new_n813), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1013), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT47), .Z(new_n1033));
  OAI221_X1 g0833(.A(new_n1003), .B1(new_n852), .B2(new_n1005), .C1(new_n1033), .C2(new_n904), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n788), .A2(G1), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n776), .A2(new_n636), .A3(new_n629), .A4(new_n705), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n707), .B2(new_n713), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n703), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n702), .A2(G330), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n1037), .C1(new_n707), .C2(new_n713), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n770), .B1(new_n872), .B2(new_n766), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n783), .B(new_n1042), .C1(new_n1043), .C2(new_n869), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT107), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT44), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT105), .B1(new_n648), .B2(new_n705), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT105), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n673), .A2(new_n1049), .A3(new_n699), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n699), .B1(new_n537), .B2(new_n541), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n684), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1047), .B1(new_n714), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n709), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1037), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1048), .A2(new_n1050), .B1(new_n684), .B2(new_n1052), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(KEYINPUT44), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT45), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1054), .A2(new_n1037), .A3(KEYINPUT45), .A4(new_n1056), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1060), .A2(new_n708), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n708), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n771), .A2(KEYINPUT107), .A3(new_n783), .A4(new_n1042), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1046), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT108), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT108), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1046), .A2(new_n1067), .A3(new_n1071), .A4(new_n1068), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n784), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n717), .B(KEYINPUT41), .Z(new_n1074));
  OAI21_X1  g0874(.A(new_n1036), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n703), .A2(new_n707), .A3(new_n1054), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT106), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1077), .B(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1058), .A2(new_n1037), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT42), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n648), .B1(new_n1058), .B2(new_n636), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n705), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1082), .A2(new_n1084), .B1(KEYINPUT43), .B2(new_n1005), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1080), .B(new_n1085), .Z(new_n1086));
  AND3_X1   g0886(.A1(new_n1075), .A2(KEYINPUT109), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT109), .B1(new_n1075), .B2(new_n1086), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1034), .B1(new_n1087), .B2(new_n1088), .ZN(G387));
  OAI22_X1  g0889(.A1(new_n1016), .A2(new_n813), .B1(new_n816), .B2(new_n1029), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n833), .A2(G322), .B1(new_n834), .B2(new_n1024), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT48), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1009), .A2(G283), .B1(new_n1018), .B2(G294), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT49), .Z(new_n1100));
  AOI21_X1  g0900(.A(new_n292), .B1(new_n830), .B2(G326), .ZN(new_n1101));
  INV_X1    g0901(.A(G116), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n826), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1009), .A2(new_n367), .B1(G150), .B2(new_n830), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n301), .B1(new_n1018), .B2(G77), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1105), .A2(new_n1015), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G159), .A2(new_n833), .B1(new_n834), .B2(new_n369), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n221), .C2(new_n813), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G68), .B2(new_n817), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n804), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n720), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n793), .A2(new_n1112), .B1(new_n356), .B2(new_n716), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n241), .A2(new_n285), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n369), .A2(new_n221), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT50), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n720), .B(new_n285), .C1(new_n203), .C2(new_n252), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n796), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1113), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n789), .B1(new_n1119), .B2(new_n805), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1111), .B(new_n1120), .C1(new_n707), .C2(new_n852), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1042), .A2(new_n1035), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1046), .A2(new_n1068), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1124), .B(new_n717), .C1(new_n785), .C2(new_n1042), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(G393));
  INV_X1    g0926(.A(new_n717), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1067), .B1(new_n1046), .B2(new_n1068), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1067), .A2(new_n1035), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1058), .A2(new_n803), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n814), .A2(G311), .B1(G317), .B2(new_n833), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT52), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n292), .B(new_n843), .C1(G283), .C2(new_n1018), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1009), .A2(G116), .B1(new_n830), .B2(G322), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n825), .B2(new_n816), .C1(new_n1029), .C2(new_n1022), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n813), .A2(new_n838), .B1(new_n334), .B2(new_n899), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT51), .Z(new_n1140));
  NOR2_X1   g0940(.A1(new_n824), .A2(new_n252), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n292), .B1(new_n203), .B2(new_n820), .C1(new_n826), .C2(new_n552), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G143), .C2(new_n830), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n221), .B2(new_n1022), .C1(new_n333), .C2(new_n816), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1134), .A2(new_n1138), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n804), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n246), .A2(new_n797), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n805), .B1(new_n538), .B2(new_n212), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n790), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1130), .B1(new_n1132), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1129), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G390));
  OAI21_X1  g0952(.A(new_n945), .B1(new_n915), .B2(new_n924), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n966), .A2(new_n1153), .A3(new_n968), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n875), .A2(new_n858), .A3(new_n923), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n857), .A2(new_n381), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n780), .A2(new_n705), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n381), .B2(new_n699), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n923), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n945), .A3(new_n975), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1154), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n992), .A2(G330), .A3(new_n977), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n992), .A2(new_n452), .A3(G330), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n668), .A2(new_n972), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n915), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n923), .B1(new_n875), .B2(new_n858), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n989), .A2(new_n869), .A3(new_n984), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(G330), .B(new_n858), .C1(new_n982), .C2(new_n764), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1158), .B1(new_n1171), .B2(new_n924), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1155), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1166), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1127), .B1(new_n1164), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT114), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1169), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1154), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1166), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1172), .A2(new_n1155), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n924), .B1(new_n771), .B2(new_n976), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n915), .B1(new_n1183), .B2(new_n1162), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1181), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1176), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1176), .B(new_n1185), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1175), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n966), .A2(new_n801), .A3(new_n968), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n881), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n790), .B1(new_n369), .B2(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n356), .A2(new_n1022), .B1(new_n899), .B2(new_n827), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n301), .B1(new_n552), .B2(new_n820), .C1(new_n826), .C2(new_n203), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n829), .A2(new_n825), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1193), .A2(new_n1141), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n538), .B2(new_n816), .C1(new_n1102), .C2(new_n813), .ZN(new_n1197));
  INV_X1    g0997(.A(G128), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n813), .A2(new_n884), .B1(new_n1198), .B2(new_n899), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT116), .Z(new_n1200));
  NOR3_X1   g1000(.A1(new_n820), .A2(KEYINPUT53), .A3(new_n334), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT53), .B1(new_n820), .B2(new_n334), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n292), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n834), .C2(G137), .ZN(new_n1204));
  INV_X1    g1004(.A(G125), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n824), .A2(new_n838), .B1(new_n829), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G50), .B2(new_n1014), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT54), .B(G143), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1204), .B(new_n1207), .C1(new_n816), .C2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1197), .B1(new_n1200), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1192), .B1(new_n1210), .B2(new_n804), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1190), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT115), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1180), .B2(new_n1036), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1164), .A2(KEYINPUT115), .A3(new_n1035), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1213), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1189), .A2(new_n1217), .ZN(G378));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n340), .A2(new_n930), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n662), .B2(new_n343), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1220), .B(new_n342), .C1(new_n660), .C2(new_n661), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT117), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n354), .A2(new_n1220), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT117), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n662), .A2(new_n343), .A3(new_n1221), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1229));
  AND3_X1   g1029(.A1(new_n1224), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1230), .A2(new_n1231), .A3(KEYINPUT118), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n994), .B2(G330), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n869), .B(new_n1232), .C1(new_n991), .C2(new_n993), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1234), .A2(new_n1235), .B1(new_n969), .B2(new_n944), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1232), .B1(new_n988), .B2(new_n869), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n994), .A2(G330), .A3(new_n1233), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n945), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n962), .A2(new_n964), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n967), .B1(new_n1240), .B2(new_n953), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n968), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1239), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n925), .A2(new_n941), .B1(new_n655), .B2(new_n930), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1237), .A2(new_n1238), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1236), .A2(new_n1245), .A3(KEYINPUT119), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT119), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n970), .A2(new_n1247), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1166), .B1(new_n1164), .B2(new_n1174), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1219), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1183), .A2(new_n1162), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1252), .A2(new_n1167), .B1(new_n1172), .B2(new_n1155), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1181), .B1(new_n1180), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1219), .B1(new_n1236), .B2(new_n1245), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1127), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1251), .A2(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n538), .A2(new_n1022), .B1(new_n899), .B2(new_n1102), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n292), .A2(G41), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n252), .B2(new_n820), .C1(new_n824), .C2(new_n203), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n202), .A2(new_n826), .B1(new_n829), .B2(new_n827), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1258), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n356), .B2(new_n813), .C1(new_n563), .C2(new_n816), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT58), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1259), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G50), .B1(new_n459), .B2(new_n284), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1263), .A2(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n824), .A2(new_n334), .B1(new_n820), .B2(new_n1208), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n899), .A2(new_n1205), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(G132), .C2(new_n834), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1270), .B1(new_n1198), .B2(new_n813), .C1(new_n1007), .C2(new_n816), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT59), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n459), .B(new_n284), .C1(new_n826), .C2(new_n838), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G124), .B2(new_n830), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1271), .A2(KEYINPUT59), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n1267), .B1(new_n1264), .B2(new_n1263), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n804), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1278), .B(new_n790), .C1(G50), .C2(new_n1191), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1230), .A2(new_n1231), .A3(new_n802), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1249), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1035), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1257), .A2(new_n1283), .ZN(G375));
  NAND2_X1  g1084(.A1(new_n1253), .A2(new_n1166), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1074), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1185), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n924), .A2(new_n801), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n790), .B1(G68), .B2(new_n1191), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n884), .A2(new_n899), .B1(new_n1022), .B2(new_n1208), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n826), .A2(new_n202), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n292), .B1(new_n820), .B2(new_n838), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n824), .A2(new_n221), .B1(new_n829), .B2(new_n1198), .ZN(new_n1293));
  NOR4_X1   g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n1294), .B1(new_n1007), .B2(new_n813), .C1(new_n334), .C2(new_n816), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n814), .A2(G283), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n292), .B(new_n1006), .C1(G97), .C2(new_n1018), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1009), .A2(new_n367), .B1(G303), .B2(new_n830), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(G116), .A2(new_n834), .B1(new_n833), .B2(G294), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n816), .A2(new_n356), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1295), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1289), .B1(new_n1302), .B2(new_n804), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1288), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1253), .B2(new_n1036), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1287), .A2(new_n1306), .ZN(G381));
  NOR2_X1   g1107(.A1(G375), .A2(G378), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G387), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1123), .A2(new_n854), .A3(new_n1125), .ZN(new_n1311));
  NOR4_X1   g1111(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT120), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1309), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1315), .B2(new_n1314), .ZN(G407));
  INV_X1    g1117(.A(G213), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1318), .A2(G343), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(KEYINPUT121), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G407), .B(G213), .C1(new_n1309), .C2(new_n1320), .ZN(G409));
  NAND2_X1  g1121(.A1(G393), .A2(G396), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT125), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1322), .A2(new_n1323), .A3(new_n1311), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1322), .B2(new_n1311), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G387), .A2(new_n1151), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1034), .B(G390), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1327), .A2(new_n1326), .A3(new_n1328), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1257), .A2(G378), .A3(new_n1283), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1254), .A2(new_n1286), .A3(new_n1248), .A4(new_n1246), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1236), .A2(new_n1245), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1281), .B1(new_n1335), .B2(new_n1035), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n1189), .A3(new_n1217), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1319), .B1(new_n1333), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT60), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1285), .B1(new_n1174), .B2(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1170), .A2(KEYINPUT60), .A3(new_n1166), .A4(new_n1173), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1342), .A2(new_n717), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(G384), .B1(new_n1344), .B2(new_n1306), .ZN(new_n1345));
  INV_X1    g1145(.A(G384), .ZN(new_n1346));
  AOI211_X1 g1146(.A(new_n1346), .B(new_n1305), .C1(new_n1341), .C2(new_n1343), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1339), .A2(KEYINPUT122), .A3(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(KEYINPUT122), .B1(new_n1339), .B2(new_n1348), .ZN(new_n1351));
  NOR3_X1   g1151(.A1(new_n1350), .A2(KEYINPUT62), .A3(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1333), .A2(new_n1338), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1320), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1348), .ZN(new_n1355));
  OAI21_X1  g1155(.A(KEYINPUT62), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(G2897), .ZN(new_n1357));
  OAI22_X1  g1157(.A1(new_n1345), .A2(new_n1347), .B1(new_n1357), .B2(new_n1320), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1357), .B1(new_n1348), .B2(KEYINPUT124), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT124), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1319), .B1(new_n1360), .B2(G2897), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1358), .B1(new_n1359), .B2(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT61), .B1(new_n1354), .B2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1356), .A2(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1332), .B1(new_n1352), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT123), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1362), .B1(new_n1339), .B2(new_n1366), .ZN(new_n1367));
  AOI211_X1 g1167(.A(KEYINPUT123), .B(new_n1319), .C1(new_n1333), .C2(new_n1338), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1353), .A2(KEYINPUT63), .A3(new_n1320), .A4(new_n1348), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT61), .ZN(new_n1371));
  NAND4_X1  g1171(.A1(new_n1370), .A2(new_n1371), .A3(new_n1330), .A4(new_n1331), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1369), .A2(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT63), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1374), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1375));
  AOI21_X1  g1175(.A(KEYINPUT126), .B1(new_n1373), .B2(new_n1375), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1327), .A2(new_n1326), .A3(new_n1328), .ZN(new_n1377));
  NOR3_X1   g1177(.A1(new_n1377), .A2(new_n1329), .A3(KEYINPUT61), .ZN(new_n1378));
  OAI211_X1 g1178(.A(new_n1378), .B(new_n1370), .C1(new_n1368), .C2(new_n1367), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1319), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1353), .A2(new_n1380), .A3(new_n1348), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT122), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(KEYINPUT63), .B1(new_n1383), .B2(new_n1349), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT126), .ZN(new_n1385));
  NOR3_X1   g1185(.A1(new_n1379), .A2(new_n1384), .A3(new_n1385), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1365), .B1(new_n1376), .B2(new_n1386), .ZN(G405));
  AND2_X1   g1187(.A1(G375), .A2(G378), .ZN(new_n1388));
  NOR2_X1   g1188(.A1(new_n1388), .A2(new_n1308), .ZN(new_n1389));
  XNOR2_X1  g1189(.A(new_n1389), .B(new_n1348), .ZN(new_n1390));
  XNOR2_X1  g1190(.A(new_n1390), .B(new_n1332), .ZN(G402));
endmodule


