//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n466), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n466), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(G136), .B2(new_n465), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT66), .Z(G162));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(KEYINPUT68), .C1(new_n463), .C2(new_n462), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT67), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n483), .B(new_n486), .C1(new_n463), .C2(new_n462), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(KEYINPUT4), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n484), .A2(KEYINPUT67), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n488), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  OR2_X1    g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n505), .A2(new_n510), .ZN(G166));
  NAND2_X1  g086(.A1(new_n509), .A2(KEYINPUT69), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n512), .A2(new_n515), .A3(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT70), .B(G51), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n519));
  AND3_X1   g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  NAND2_X1  g097(.A1(G63), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n509), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n521), .A2(new_n522), .B1(new_n525), .B2(new_n502), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n502), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n509), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G651), .B1(new_n533), .B2(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n516), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  AOI22_X1  g112(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n504), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(new_n533), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n512), .A2(new_n515), .A3(G543), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n539), .A2(KEYINPUT72), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  AOI22_X1  g127(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(KEYINPUT74), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n504), .B1(new_n553), .B2(KEYINPUT74), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n554), .A2(new_n555), .B1(G91), .B2(new_n533), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n516), .A2(new_n557), .A3(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n544), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n559), .B1(new_n558), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(G299));
  XNOR2_X1  g139(.A(new_n527), .B(KEYINPUT75), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND2_X1  g141(.A1(new_n516), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n533), .A2(G87), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n500), .B2(new_n501), .ZN(new_n572));
  AND2_X1   g147(.A1(G73), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n500), .B2(new_n501), .ZN(new_n576));
  AND2_X1   g151(.A1(G48), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n513), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT76), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n504), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n542), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n583), .A2(new_n584), .B1(new_n544), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT78), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  INV_X1    g169(.A(G79), .ZN(new_n595));
  INV_X1    g170(.A(G543), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n530), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n599), .B1(new_n595), .B2(new_n596), .C1(new_n530), .C2(new_n594), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(G651), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n502), .A2(new_n513), .A3(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n516), .A2(G54), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n593), .B1(new_n608), .B2(G868), .ZN(G284));
  XNOR2_X1  g184(.A(G284), .B(KEYINPUT81), .ZN(G321));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g186(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n608), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n608), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(G111), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G2105), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n465), .A2(G135), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT83), .ZN(new_n623));
  AOI211_X1 g198(.A(new_n621), .B(new_n623), .C1(G123), .C2(new_n475), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT82), .B(G2100), .ZN(new_n626));
  INV_X1    g201(.A(new_n464), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n467), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n626), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n631), .B(new_n632), .C1(new_n625), .C2(new_n624), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT84), .ZN(G156));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT86), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n638), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n645), .A3(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n635), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n653), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n656), .A2(KEYINPUT87), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(KEYINPUT87), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(G401));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT88), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n625), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT89), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n683), .C1(new_n674), .C2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT90), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n689), .A2(new_n692), .A3(new_n690), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n580), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(G23), .ZN(new_n707));
  INV_X1    g282(.A(G288), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n701), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n700), .A2(new_n706), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT34), .Z(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G24), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n590), .B2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT93), .B(G1986), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(G107), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G2105), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G119), .B2(new_n475), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n465), .A2(G131), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT91), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(new_n720), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n714), .A2(new_n719), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT36), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n701), .A2(G5), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G171), .B2(new_n701), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1961), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT31), .B(G11), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT30), .B(G28), .Z(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G29), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n624), .B2(G29), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n720), .B1(KEYINPUT24), .B2(G34), .ZN(new_n745));
  OAI22_X1  g320(.A1(G160), .A2(new_n720), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n743), .B1(G2084), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n739), .B(new_n747), .C1(G2084), .C2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n701), .A2(G19), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n547), .B2(new_n701), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1341), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n720), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n465), .A2(G140), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n475), .A2(G128), .ZN(new_n755));
  OR2_X1    g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(new_n720), .ZN(new_n760));
  INV_X1    g335(.A(G2067), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n701), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G168), .B2(new_n701), .ZN(new_n764));
  INV_X1    g339(.A(G1966), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n748), .A2(new_n751), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G129), .B2(new_n475), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n465), .A2(G141), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n467), .A2(G105), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n467), .A2(KEYINPUT98), .A3(G105), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n770), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n778), .A2(KEYINPUT100), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(KEYINPUT100), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G29), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT101), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G29), .B2(G32), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n784), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  AOI21_X1  g363(.A(new_n767), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G4), .A2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  INV_X1    g366(.A(new_n608), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n701), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n789), .B(new_n794), .C1(new_n787), .C2(new_n788), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n627), .A2(G127), .ZN(new_n796));
  NAND2_X1  g371(.A1(G115), .A2(G2104), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n466), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(KEYINPUT97), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(KEYINPUT97), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT25), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n465), .A2(G139), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n800), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n720), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n720), .B2(G33), .ZN(new_n808));
  INV_X1    g383(.A(G2072), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n720), .A2(G27), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G164), .B2(new_n720), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n808), .A2(new_n809), .B1(G2078), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(G2078), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n812), .B(new_n813), .C1(new_n809), .C2(new_n808), .ZN(new_n814));
  NOR2_X1   g389(.A1(G29), .A2(G35), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G162), .B2(G29), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT29), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G2090), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n701), .A2(G20), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT23), .ZN(new_n822));
  INV_X1    g397(.A(G299), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n701), .ZN(new_n824));
  INV_X1    g399(.A(G1956), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n820), .B(new_n826), .C1(new_n819), .C2(new_n818), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n736), .A2(new_n795), .A3(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(G67), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n530), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n504), .B1(new_n832), .B2(KEYINPUT102), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(KEYINPUT102), .B2(new_n832), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT103), .B(G55), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n516), .A2(new_n835), .B1(G93), .B2(new_n533), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n608), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT104), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  INV_X1    g417(.A(new_n837), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n547), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n842), .B(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n839), .B1(new_n846), .B2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n729), .B(new_n629), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n494), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n489), .A2(KEYINPUT105), .A3(new_n493), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n488), .A2(new_n497), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n758), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n780), .A2(new_n781), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n780), .B2(new_n781), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n806), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT106), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n856), .B(KEYINPUT107), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n778), .A2(new_n779), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n806), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT106), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n857), .A2(new_n865), .A3(new_n806), .A4(new_n858), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n860), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n465), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n475), .A2(G130), .ZN(new_n869));
  OR2_X1    g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n867), .A2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n851), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n850), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G162), .B(new_n473), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n624), .Z(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n877), .A2(new_n879), .A3(new_n882), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g463(.A(new_n615), .B(new_n844), .ZN(new_n889));
  XNOR2_X1  g464(.A(G299), .B(new_n605), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(KEYINPUT41), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n590), .B(new_n580), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(G303), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT42), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n893), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G868), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(G868), .B2(new_n843), .ZN(G331));
  XOR2_X1   g475(.A(G331), .B(KEYINPUT108), .Z(G295));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n902));
  NOR2_X1   g477(.A1(G171), .A2(G168), .ZN(new_n903));
  INV_X1    g478(.A(G286), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(G171), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n844), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n892), .ZN(new_n908));
  INV_X1    g483(.A(new_n890), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n896), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n885), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n896), .B1(new_n908), .B2(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n902), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n908), .A2(KEYINPUT109), .A3(new_n910), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n908), .A2(KEYINPUT109), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(new_n896), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n913), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n917), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n918), .ZN(new_n923));
  INV_X1    g498(.A(new_n913), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n916), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n913), .B2(new_n914), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n927), .A2(KEYINPUT110), .A3(new_n902), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT110), .B1(new_n927), .B2(new_n902), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(G397));
  INV_X1    g505(.A(G1384), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT45), .B1(new_n855), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n468), .A2(G40), .A3(new_n472), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n758), .B(G2067), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT112), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n862), .A3(G1996), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n729), .B(new_n732), .Z(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n934), .ZN(new_n941));
  INV_X1    g516(.A(G1996), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT111), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n782), .ZN(new_n945));
  NOR2_X1   g520(.A1(G290), .A2(G1986), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n934), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT48), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n939), .A2(new_n941), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  AND4_X1   g524(.A1(new_n732), .A2(new_n939), .A3(new_n730), .A4(new_n945), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n758), .A2(G2067), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n934), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n944), .A2(KEYINPUT46), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT124), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n862), .A2(new_n935), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n944), .A2(KEYINPUT46), .B1(new_n934), .B2(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n954), .B2(new_n957), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n949), .B(new_n952), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT54), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n498), .A2(new_n931), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n933), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(G2078), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT114), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n466), .A2(G138), .ZN(new_n970));
  INV_X1    g545(.A(new_n463), .ZN(new_n971));
  NAND2_X1  g546(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n486), .B1(new_n973), .B2(KEYINPUT68), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n497), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n853), .A2(new_n854), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n969), .B(new_n931), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n969), .B1(new_n855), .B2(new_n931), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n966), .B(new_n968), .C1(new_n981), .C2(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(new_n933), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n979), .B2(new_n980), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n963), .A2(new_n984), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n983), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT119), .B(G1961), .Z(new_n989));
  OAI21_X1  g564(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT120), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n982), .B(new_n992), .C1(new_n988), .C2(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n963), .A2(new_n964), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n855), .A2(KEYINPUT45), .A3(new_n931), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n933), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n967), .B1(new_n997), .B2(G2078), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT121), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G301), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n468), .A2(G40), .A3(new_n968), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT122), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n471), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n466), .B1(new_n471), .B2(new_n1003), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n996), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n988), .A2(new_n989), .B1(new_n932), .B2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n999), .A2(G171), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n962), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n558), .A2(new_n561), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n556), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(G299), .A2(KEYINPUT57), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n855), .A2(new_n931), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n984), .B1(new_n1017), .B2(new_n978), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n933), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n825), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n997), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT56), .B(G2072), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1015), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1020), .A2(new_n1015), .A3(new_n1023), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(new_n605), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT50), .B1(new_n1017), .B2(new_n978), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n933), .B1(new_n1027), .B2(new_n986), .ZN(new_n1028));
  INV_X1    g603(.A(G1348), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n981), .A2(new_n761), .A3(new_n933), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1024), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT61), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1015), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT50), .B1(new_n979), .B2(new_n980), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1019), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1956), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1020), .A2(new_n1023), .A3(new_n1015), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(KEYINPUT61), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1017), .A2(new_n933), .A3(new_n978), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  AOI22_X1  g620(.A1(new_n1021), .A2(new_n942), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n547), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT59), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n997), .A2(G1996), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(new_n547), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1035), .A2(new_n1043), .A3(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT60), .B(new_n1031), .C1(new_n988), .C2(G1348), .ZN(new_n1055));
  INV_X1    g630(.A(new_n605), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n605), .A4(new_n1031), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1057), .A2(new_n1058), .B1(new_n1059), .B2(new_n1032), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1033), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n994), .A2(G301), .A3(new_n1000), .ZN(new_n1062));
  OAI21_X1  g637(.A(G171), .B1(new_n999), .B2(new_n1008), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(KEYINPUT54), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G303), .A2(G8), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT55), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1017), .A2(new_n978), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1019), .B1(new_n1067), .B2(KEYINPUT50), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1068), .A2(new_n819), .B1(new_n704), .B2(new_n997), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1066), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n933), .A2(new_n819), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n985), .B2(new_n987), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n997), .A2(new_n704), .ZN(new_n1075));
  OAI211_X1 g650(.A(G8), .B(new_n1072), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1981), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n574), .A2(new_n578), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n574), .B2(new_n578), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT115), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT115), .B(KEYINPUT49), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1044), .A2(G8), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1044), .A2(new_n1087), .A3(new_n1084), .A4(G8), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n708), .A2(G1976), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1044), .A2(G8), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1092));
  INV_X1    g667(.A(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1044), .A2(G8), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1071), .A2(new_n1076), .A3(new_n1089), .A4(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n983), .A2(G2084), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1027), .B2(new_n986), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT45), .B1(new_n1017), .B2(new_n978), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n765), .B1(new_n1100), .B2(new_n965), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n1102), .B2(new_n527), .ZN(new_n1103));
  AOI21_X1  g678(.A(G168), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(G8), .C1(new_n1102), .C2(new_n527), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1097), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1010), .A2(new_n1061), .A3(new_n1064), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT62), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1114), .A2(new_n1071), .A3(new_n1076), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1105), .A2(new_n1116), .A3(new_n1107), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1111), .A2(new_n1001), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1102), .A2(G8), .A3(new_n904), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1097), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1119), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n819), .B(new_n933), .C1(new_n1027), .C2(new_n986), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n997), .A2(new_n704), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1070), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1125), .A2(new_n1072), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1122), .A2(new_n1126), .A3(new_n1114), .A4(new_n1076), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1044), .A2(G8), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(G1976), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1089), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1078), .B(KEYINPUT117), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1112), .A2(new_n1076), .A3(new_n1113), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1128), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1096), .A2(new_n1072), .A3(new_n1125), .A4(new_n1089), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1132), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1089), .B2(new_n1130), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1136), .B(KEYINPUT118), .C1(new_n1129), .C2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1121), .A2(new_n1127), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1109), .A2(new_n1118), .A3(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(G290), .A2(G1986), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n934), .B1(new_n1142), .B2(new_n946), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n939), .A2(new_n1143), .A3(new_n941), .A4(new_n945), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT113), .Z(new_n1145));
  AND3_X1   g720(.A1(new_n1141), .A2(KEYINPUT123), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT123), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n961), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n961), .B(KEYINPUT125), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g727(.A(new_n658), .ZN(new_n1154));
  NOR2_X1   g728(.A1(new_n656), .A2(KEYINPUT87), .ZN(new_n1155));
  OAI21_X1  g729(.A(new_n654), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g730(.A(G229), .ZN(new_n1157));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1158));
  NOR2_X1   g732(.A1(new_n460), .A2(G227), .ZN(new_n1159));
  NAND4_X1  g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n694), .A2(new_n695), .A3(new_n1159), .ZN(new_n1161));
  OAI21_X1  g735(.A(KEYINPUT126), .B1(G401), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g736(.A1(new_n926), .A2(new_n925), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g737(.A1(new_n887), .A2(new_n1163), .A3(KEYINPUT127), .ZN(new_n1164));
  AOI21_X1  g738(.A(KEYINPUT127), .B1(new_n887), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n1165), .ZN(G308));
  NAND2_X1  g740(.A1(new_n887), .A2(new_n1163), .ZN(G225));
endmodule


