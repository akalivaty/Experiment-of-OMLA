//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR3_X1   g040(.A1(new_n464), .A2(new_n465), .A3(G2105), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT66), .B1(new_n462), .B2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G101), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n462), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n471), .A2(new_n472), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n481), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT68), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(KEYINPUT69), .B1(new_n462), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n462), .A3(G138), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n482), .A2(KEYINPUT70), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n500), .A2(new_n462), .A3(G138), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n461), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(G138), .B(new_n462), .C1(new_n471), .C2(new_n472), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n499), .B1(new_n506), .B2(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(KEYINPUT71), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n517), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  AND3_X1   g105(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n532), .B1(new_n519), .B2(new_n520), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n524), .B(new_n529), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g111(.A1(KEYINPUT6), .A2(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT72), .B1(new_n519), .B2(new_n520), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(new_n539), .A3(G543), .ZN(new_n540));
  INV_X1    g115(.A(G51), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n534), .A2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n540), .A2(new_n545), .B1(new_n546), .B2(new_n533), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n516), .B2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AND3_X1   g127(.A1(new_n538), .A2(new_n539), .A3(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n531), .A2(new_n532), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(new_n533), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G81), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n540), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n535), .A2(new_n537), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(KEYINPUT72), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n573), .A2(new_n574), .A3(G53), .A4(new_n538), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n556), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n560), .B2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G166), .ZN(G303));
  OAI21_X1  g157(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n533), .A2(KEYINPUT74), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT74), .B1(new_n533), .B2(new_n586), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n553), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AND3_X1   g166(.A1(new_n572), .A2(G48), .A3(G543), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n533), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n514), .A2(new_n572), .A3(KEYINPUT77), .A4(G86), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(G61), .B1(new_n531), .B2(new_n532), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n516), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI211_X1 g177(.A(KEYINPUT76), .B(new_n516), .C1(new_n598), .C2(new_n599), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n560), .A2(G85), .ZN(new_n605));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  OAI221_X1 g182(.A(new_n605), .B1(new_n540), .B2(new_n606), .C1(new_n516), .C2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n560), .A2(G92), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT10), .Z(new_n613));
  AOI22_X1  g188(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n516), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G54), .B2(new_n553), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n611), .B1(new_n618), .B2(G868), .ZN(G321));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(G299), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(G168), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(new_n621), .B2(G168), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NOR2_X1   g201(.A1(new_n617), .A2(G559), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT79), .Z(new_n628));
  OAI21_X1  g203(.A(KEYINPUT80), .B1(new_n628), .B2(new_n621), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(KEYINPUT79), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(new_n631), .A3(G868), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n632), .C1(G868), .C2(new_n563), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g209(.A1(new_n468), .A2(new_n482), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n480), .A2(G123), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n483), .A2(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n462), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT17), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT84), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  INV_X1    g248(.A(new_n666), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n670), .C1(new_n674), .C2(new_n668), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n668), .A3(new_n669), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n686), .A2(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n693), .C1(new_n683), .C2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  XNOR2_X1  g275(.A(KEYINPUT86), .B(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(G6), .A2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(G305), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(G23), .ZN(new_n712));
  INV_X1    g287(.A(G288), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n707), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n711), .B(new_n716), .C1(new_n708), .C2(new_n709), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n480), .A2(G119), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n483), .A2(G131), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n462), .A2(G107), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G25), .B(new_n724), .S(G29), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n718), .B2(KEYINPUT34), .ZN(new_n729));
  MUX2_X1   g304(.A(G24), .B(G290), .S(new_n701), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT87), .ZN(new_n731));
  INV_X1    g306(.A(G1986), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n719), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT36), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n480), .A2(G129), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n483), .A2(G141), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT26), .Z(new_n739));
  INV_X1    g314(.A(G105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n737), .B(new_n739), .C1(new_n740), .C2(new_n468), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n743), .B2(G32), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n707), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n707), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n745), .A2(new_n746), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n747), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n701), .A2(G19), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n563), .B2(new_n701), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1341), .Z(new_n755));
  OR2_X1    g330(.A1(G29), .A2(G33), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n461), .A2(G127), .ZN(new_n757));
  AND2_X1   g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  OAI21_X1  g333(.A(G2105), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n483), .A2(G139), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n756), .B1(new_n764), .B2(new_n743), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  NAND2_X1  g344(.A1(G160), .A2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n771), .B2(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT24), .B2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  INV_X1    g351(.A(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n780), .B1(new_n645), .B2(new_n743), .C1(new_n774), .C2(new_n769), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n745), .B2(new_n746), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n752), .A2(new_n755), .A3(new_n775), .A4(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2090), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n743), .A2(G35), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT91), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G162), .B2(new_n743), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT29), .Z(new_n788));
  AOI21_X1  g363(.A(new_n783), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n743), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n480), .A2(G128), .ZN(new_n792));
  NOR2_X1   g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT88), .Z(new_n794));
  INV_X1    g369(.A(G116), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n465), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n794), .A2(new_n796), .B1(new_n483), .B2(G140), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n798), .A2(KEYINPUT89), .A3(G29), .ZN(new_n799));
  AOI21_X1  g374(.A(KEYINPUT89), .B1(new_n798), .B2(G29), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n791), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G2067), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n618), .A2(new_n707), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G4), .B2(new_n707), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n743), .A2(G27), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G164), .B2(new_n743), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G2078), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n805), .B2(new_n806), .ZN(new_n811));
  NOR2_X1   g386(.A1(G5), .A2(G16), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G171), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT90), .B(G1961), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AND4_X1   g390(.A1(new_n803), .A2(new_n807), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n789), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n788), .A2(new_n784), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT92), .B(KEYINPUT23), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  INV_X1    g395(.A(G20), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n701), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G16), .B2(G299), .ZN(new_n824));
  INV_X1    g399(.A(G1956), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n818), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n817), .B1(KEYINPUT94), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(KEYINPUT94), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n735), .A2(new_n828), .A3(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NAND2_X1  g406(.A1(new_n560), .A2(G93), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n832), .B1(new_n540), .B2(new_n833), .C1(new_n516), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n618), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n835), .B(new_n562), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT95), .Z(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n841), .B2(new_n842), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n837), .B1(new_n844), .B2(new_n846), .ZN(G145));
  XOR2_X1   g422(.A(KEYINPUT98), .B(G37), .Z(new_n848));
  XOR2_X1   g423(.A(new_n645), .B(G160), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n488), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT70), .B1(new_n482), .B2(new_n501), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n461), .A2(new_n504), .A3(new_n503), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n508), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(G126), .A2(new_n479), .B1(new_n494), .B2(new_n496), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n798), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n742), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n764), .A2(KEYINPUT96), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n764), .A2(KEYINPUT96), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n483), .A2(G142), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n462), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G130), .B2(new_n480), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n724), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n637), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n860), .A2(new_n862), .ZN(new_n872));
  INV_X1    g447(.A(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n851), .B(new_n871), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT99), .B1(new_n872), .B2(new_n873), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n848), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n874), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n872), .A2(new_n879), .A3(new_n873), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n851), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(G395));
  XNOR2_X1  g461(.A(G290), .B(G303), .ZN(new_n887));
  XNOR2_X1  g462(.A(G288), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n840), .B(KEYINPUT100), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n630), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n617), .B(G299), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT41), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n630), .A2(new_n890), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n893), .ZN(new_n897));
  INV_X1    g472(.A(new_n890), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n628), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n899), .B2(new_n891), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n896), .A2(new_n900), .A3(KEYINPUT42), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n893), .B(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n905), .A3(new_n891), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n902), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n889), .B1(new_n901), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n896), .B2(new_n900), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n902), .A3(new_n906), .ZN(new_n910));
  INV_X1    g485(.A(new_n889), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n621), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n835), .A2(new_n621), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT101), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n901), .A2(new_n907), .A3(new_n889), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n909), .B2(new_n910), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n914), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n916), .A2(new_n921), .ZN(G295));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n914), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n840), .B(G301), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(G168), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(G168), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n894), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n897), .B1(new_n926), .B2(new_n927), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n889), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n889), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n924), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n936), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n931), .A2(new_n848), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n935), .B1(new_n940), .B2(new_n924), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT44), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n937), .A2(new_n939), .A3(new_n924), .A4(new_n938), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n933), .B2(new_n934), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(G397));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  XOR2_X1   g524(.A(KEYINPUT103), .B(G1384), .Z(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(G164), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G160), .A2(G40), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT104), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT46), .Z(new_n957));
  XNOR2_X1  g532(.A(new_n798), .B(new_n802), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT105), .ZN(new_n959));
  INV_X1    g534(.A(new_n742), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n953), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n965), .B(KEYINPUT106), .Z(new_n966));
  INV_X1    g541(.A(new_n953), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n967), .A2(new_n954), .A3(new_n742), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n956), .B2(new_n742), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n724), .A2(new_n727), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n724), .A2(new_n727), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n953), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n967), .A2(G290), .A3(G1986), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT48), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n964), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n972), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n792), .A2(new_n802), .A3(new_n797), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n967), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(KEYINPUT107), .A2(KEYINPUT55), .ZN(new_n982));
  AND2_X1   g557(.A1(KEYINPUT107), .A2(KEYINPUT55), .ZN(new_n983));
  OAI211_X1 g558(.A(G303), .B(G8), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(G166), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n986), .B2(new_n983), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n470), .A2(new_n989), .A3(new_n475), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n854), .B2(new_n855), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT50), .B(G1384), .C1(new_n854), .C2(new_n855), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n950), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n856), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n990), .C1(KEYINPUT45), .C2(new_n991), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n995), .A2(new_n784), .B1(new_n998), .B2(new_n704), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n988), .B1(new_n999), .B2(new_n985), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n998), .A2(new_n704), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n993), .A2(new_n994), .A3(G2090), .ZN(new_n1002));
  OAI211_X1 g577(.A(G8), .B(new_n987), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n597), .B(new_n1005), .C1(new_n602), .C2(new_n603), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n572), .A2(G48), .A3(G543), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n594), .B2(new_n533), .ZN(new_n1008));
  OAI21_X1  g583(.A(G1981), .B1(new_n1008), .B2(new_n600), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(KEYINPUT49), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1006), .B(new_n1009), .C1(new_n1011), .C2(KEYINPUT49), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n1015), .B(new_n985), .C1(new_n991), .C2(new_n990), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n991), .A2(new_n990), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT108), .B1(new_n1017), .B2(G8), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1013), .B(new_n1014), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n713), .A2(G1976), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1020), .B(new_n1022), .C1(new_n1018), .C2(new_n1016), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G288), .A2(new_n1021), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1017), .A2(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n1015), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1017), .A2(KEYINPUT108), .A3(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1019), .B(new_n1023), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1018), .A2(new_n1016), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n1033), .B2(new_n1024), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(KEYINPUT110), .A3(new_n1019), .A4(new_n1023), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1004), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n825), .B1(new_n993), .B2(new_n994), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n856), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n949), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT56), .B(G2072), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n990), .A3(new_n997), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n576), .A2(new_n1043), .A3(new_n580), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n576), .B2(new_n580), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1037), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT113), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT61), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT122), .B(G2078), .Z(new_n1052));
  NOR3_X1   g627(.A1(new_n952), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n997), .A3(new_n951), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT119), .B(G1961), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n993), .B2(new_n994), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n990), .B1(new_n991), .B2(KEYINPUT45), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n949), .B(new_n950), .C1(new_n854), .C2(new_n855), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(G2078), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1054), .B(new_n1056), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1050), .B1(new_n1062), .B2(G171), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1040), .A2(new_n1064), .A3(new_n990), .A4(new_n997), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n991), .A2(new_n992), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n990), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1065), .A2(new_n1060), .B1(new_n1068), .B2(new_n1055), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1057), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT111), .B(new_n990), .C1(new_n991), .C2(KEYINPUT45), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1051), .A2(G2078), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(G301), .A3(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1048), .A2(new_n1049), .B1(new_n1063), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G286), .A2(G8), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1078), .B(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1068), .B2(G2084), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n995), .A2(KEYINPUT112), .A3(new_n769), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1083), .A2(new_n1084), .B1(new_n1085), .B2(new_n747), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1081), .B1(new_n1086), .B2(new_n985), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT111), .B1(new_n1040), .B2(new_n990), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n747), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT112), .B1(new_n995), .B2(new_n769), .ZN(new_n1093));
  NOR4_X1   g668(.A1(new_n993), .A2(new_n994), .A3(new_n1082), .A4(G2084), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1089), .B1(new_n1095), .B2(new_n1080), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1081), .B(new_n1089), .C1(new_n1086), .C2(new_n985), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1036), .A2(new_n1077), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1065), .A2(new_n1060), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(G301), .A3(new_n1056), .A4(new_n1054), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT123), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1069), .A2(new_n1104), .A3(G301), .A4(new_n1054), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g681(.A(KEYINPUT121), .B(G301), .C1(new_n1069), .C2(new_n1075), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1101), .A2(new_n1075), .A3(new_n1056), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(G171), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1100), .B1(new_n1111), .B2(KEYINPUT54), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n995), .A2(G1348), .B1(G2067), .B2(new_n1017), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n617), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1114), .B2(new_n1113), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1017), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT58), .B(G1341), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n998), .A2(G1996), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n563), .A3(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1121), .A2(KEYINPUT116), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(KEYINPUT61), .A3(new_n1047), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1068), .A2(new_n806), .B1(new_n802), .B2(new_n1117), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n617), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1116), .A2(new_n1122), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1121), .A2(KEYINPUT116), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1119), .A2(new_n563), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(KEYINPUT59), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1126), .A2(new_n617), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1132), .A2(KEYINPUT114), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1124), .B1(new_n1132), .B2(KEYINPUT114), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1128), .A2(new_n1131), .B1(new_n1135), .B2(new_n1048), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1110), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1109), .A2(new_n1108), .A3(G171), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT124), .B(new_n1050), .C1(new_n1139), .C2(new_n1106), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1099), .A2(new_n1112), .A3(new_n1136), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1006), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G288), .A2(G1976), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1019), .B2(new_n1143), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1030), .A2(new_n1003), .B1(new_n1144), .B2(new_n1033), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1004), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1086), .A2(new_n985), .A3(G286), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1004), .A2(new_n1150), .A3(new_n1030), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1148), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1145), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1141), .A2(KEYINPUT125), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT125), .B1(new_n1141), .B2(new_n1154), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1036), .B(new_n1139), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1158), .B2(new_n1157), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1155), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G290), .B(new_n732), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n970), .B(new_n973), .C1(new_n967), .C2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n981), .B1(new_n1161), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g739(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1166));
  OAI21_X1  g740(.A(new_n1166), .B1(new_n878), .B2(new_n883), .ZN(new_n1167));
  AOI21_X1  g741(.A(new_n1167), .B1(new_n944), .B2(new_n943), .ZN(G308));
  OAI211_X1 g742(.A(new_n945), .B(new_n1166), .C1(new_n883), .C2(new_n878), .ZN(G225));
endmodule


