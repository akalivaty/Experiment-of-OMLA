//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n462), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n463), .B2(new_n464), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n484), .B(new_n487), .C1(new_n464), .C2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n462), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n477), .A2(G126), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G50), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT66), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n508), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(new_n499), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n503), .A2(new_n502), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n497), .A2(new_n498), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n521), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n509), .A2(new_n510), .B1(new_n497), .B2(new_n498), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT67), .B(G90), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n530), .B1(new_n519), .B2(new_n531), .C1(new_n508), .C2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  AOI22_X1  g109(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n499), .A2(G43), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n506), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT68), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  NOR3_X1   g121(.A1(new_n503), .A2(new_n502), .A3(KEYINPUT70), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n509), .B2(new_n510), .ZN(new_n549));
  OAI21_X1  g124(.A(G65), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT69), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n509), .A2(new_n548), .A3(new_n510), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT70), .B1(new_n503), .B2(new_n502), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT71), .B1(new_n559), .B2(new_n553), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n560), .A3(G651), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n519), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n499), .A2(new_n564), .A3(G53), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n563), .A2(new_n565), .B1(G91), .B2(new_n528), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(G168), .A2(KEYINPUT72), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(new_n521), .B2(new_n526), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G286));
  OR2_X1    g147(.A1(new_n507), .A2(new_n515), .ZN(G303));
  NAND2_X1  g148(.A1(new_n528), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n499), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n522), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n499), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n528), .A2(new_n582), .A3(G86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n511), .A2(new_n523), .A3(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT73), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n528), .A2(G85), .B1(new_n499), .B2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n508), .B2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n528), .B2(G92), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  NOR3_X1   g170(.A1(new_n506), .A2(KEYINPUT74), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n528), .A2(new_n593), .A3(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT74), .B1(new_n506), .B2(new_n595), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT10), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n557), .B2(new_n558), .ZN(new_n603));
  AND2_X1   g178(.A1(G79), .A2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n499), .A2(G54), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n601), .A2(KEYINPUT75), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n597), .A2(new_n606), .A3(new_n605), .A4(new_n600), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n591), .B1(new_n613), .B2(new_n590), .ZN(G284));
  AOI21_X1  g189(.A(new_n591), .B1(new_n613), .B2(new_n590), .ZN(G321));
  NOR2_X1   g190(.A1(G299), .A2(G868), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n571), .ZN(G297));
  AOI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n571), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND3_X1  g195(.A1(new_n608), .A2(new_n619), .A3(new_n611), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n475), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n477), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n462), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT3), .B(G2104), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n469), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  AND2_X1   g210(.A1(new_n635), .A2(G2100), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(KEYINPUT77), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(KEYINPUT77), .ZN(new_n639));
  OAI221_X1 g214(.A(new_n630), .B1(G2100), .B2(new_n635), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT78), .ZN(G156));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT80), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT81), .Z(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT82), .Z(G401));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT83), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n664), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(KEYINPUT85), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(new_n670), .A3(new_n662), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n670), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(new_n664), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n674), .A2(new_n662), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(new_n669), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n672), .B(new_n680), .C1(new_n677), .C2(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT88), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n688), .B1(new_n692), .B2(KEYINPUT89), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(KEYINPUT89), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n688), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n696), .B(new_n688), .S(new_n697), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n695), .A2(new_n698), .A3(new_n700), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n705), .B1(new_n702), .B2(new_n706), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n686), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n709), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n711), .A2(new_n685), .A3(new_n707), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(G229));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1971), .Z(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G23), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G288), .B2(new_n717), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n716), .A2(new_n720), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n475), .A2(G131), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n477), .A2(G119), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n462), .A2(G107), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G25), .B(new_n734), .S(G29), .Z(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G24), .B(G290), .S(G16), .Z(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G1986), .Z(new_n739));
  NAND3_X1  g314(.A1(new_n729), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G33), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n631), .A2(G127), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n747), .A2(KEYINPUT95), .A3(G2105), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT95), .B1(new_n747), .B2(G2105), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n475), .A2(G139), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n748), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n744), .B1(new_n754), .B2(new_n743), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G2072), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n717), .A2(G19), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n540), .B2(new_n717), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  INV_X1    g335(.A(G168), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  INV_X1    g338(.A(G21), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n762), .B(new_n763), .C1(G16), .C2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n760), .B1(KEYINPUT100), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT100), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G11), .Z(new_n768));
  NOR2_X1   g343(.A1(new_n629), .A2(new_n743), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT99), .B(G28), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n768), .B(new_n769), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n475), .A2(G140), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n477), .A2(G128), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n462), .A2(G116), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n743), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT94), .B(G2067), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n767), .B(new_n774), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G5), .A2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT101), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G171), .B2(G16), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n743), .A2(G27), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n494), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2078), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n743), .B1(KEYINPUT24), .B2(G34), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(KEYINPUT24), .B2(G34), .ZN(new_n796));
  INV_X1    g371(.A(G160), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G2084), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n792), .A2(new_n793), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n790), .A2(new_n794), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n762), .B1(G16), .B2(new_n764), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G1966), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n783), .A2(new_n785), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n798), .A2(new_n799), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n789), .A2(G1961), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n766), .A2(new_n786), .A3(new_n802), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n743), .A2(G35), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G162), .B2(new_n743), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT29), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G2090), .Z(new_n813));
  NOR2_X1   g388(.A1(G29), .A2(G32), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n469), .A2(G105), .ZN(new_n815));
  NAND3_X1  g390(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT26), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n815), .B(new_n817), .C1(G129), .C2(new_n477), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n475), .A2(G141), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n814), .B1(new_n824), .B2(G29), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT27), .B(G1996), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  AND4_X1   g403(.A1(new_n756), .A2(new_n809), .A3(new_n813), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n717), .A2(G20), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT102), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT23), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G299), .B2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1956), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n613), .A2(new_n717), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G4), .B2(new_n717), .ZN(new_n836));
  INV_X1    g411(.A(G1348), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n829), .A2(new_n834), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n742), .A2(new_n840), .ZN(G311));
  OR2_X1    g416(.A1(new_n742), .A2(new_n840), .ZN(G150));
  XOR2_X1   g417(.A(KEYINPUT105), .B(G860), .Z(new_n843));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n613), .A2(new_n844), .A3(G559), .ZN(new_n845));
  INV_X1    g420(.A(new_n540), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n508), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT103), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n528), .A2(G93), .B1(new_n499), .B2(G55), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n848), .B2(KEYINPUT103), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n846), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n848), .A2(KEYINPUT103), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n854), .A2(new_n540), .A3(new_n849), .A4(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT38), .B1(new_n612), .B2(new_n619), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n845), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n857), .B1(new_n845), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n843), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT104), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(KEYINPUT104), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n850), .A2(new_n852), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n843), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(G145));
  NAND2_X1  g447(.A1(new_n475), .A2(G142), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n477), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n462), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n734), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n486), .A2(new_n880), .A3(new_n488), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n486), .B2(new_n488), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n493), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n779), .ZN(new_n884));
  INV_X1    g459(.A(new_n634), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n477), .A2(G126), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n490), .A2(new_n492), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n488), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n487), .B1(new_n631), .B2(new_n484), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT106), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n486), .A2(new_n880), .A3(new_n488), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n779), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(new_n634), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n879), .B1(new_n886), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n884), .A2(new_n885), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n634), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n878), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n822), .B(KEYINPUT97), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n754), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n754), .B1(new_n904), .B2(new_n822), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n904), .B2(new_n822), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n629), .B(G160), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(G162), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n897), .A2(new_n907), .A3(new_n900), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n909), .A2(new_n916), .A3(new_n913), .A4(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n909), .A2(new_n913), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n919), .B2(new_n911), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g497(.A(G305), .B(G290), .ZN(new_n923));
  XNOR2_X1  g498(.A(G166), .B(G288), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT42), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n621), .A2(new_n857), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n856), .A2(new_n619), .A3(new_n608), .A4(new_n611), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n601), .A2(new_n561), .A3(new_n566), .A4(new_n607), .ZN(new_n930));
  NAND2_X1  g505(.A1(G299), .A2(new_n609), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT109), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n932), .B2(KEYINPUT41), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n929), .B(KEYINPUT110), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n932), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n927), .A2(new_n928), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n935), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n938), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT110), .B1(new_n947), .B2(new_n929), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT111), .B1(new_n942), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n929), .B1(new_n936), .B2(new_n938), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n941), .A4(new_n939), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n926), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(new_n926), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n869), .A2(new_n590), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(G295));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n958), .ZN(G331));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g536(.A(G301), .B1(new_n568), .B2(new_n570), .ZN(new_n962));
  NOR2_X1   g537(.A1(G171), .A2(G168), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n856), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n853), .B(new_n855), .C1(new_n962), .C2(new_n963), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n933), .B2(new_n935), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n940), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n925), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G37), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n967), .B1(new_n945), .B2(new_n946), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n974), .A2(new_n925), .A3(new_n970), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n925), .B1(new_n974), .B2(new_n970), .ZN(new_n977));
  INV_X1    g552(.A(new_n925), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n936), .A2(new_n938), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n978), .B(new_n969), .C1(new_n979), .C2(new_n967), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n977), .A2(new_n980), .A3(new_n981), .A4(new_n972), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n961), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n973), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n977), .A2(new_n980), .A3(new_n972), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(KEYINPUT43), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n983), .B1(new_n961), .B2(new_n987), .ZN(G397));
  INV_X1    g563(.A(G1961), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n894), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(G160), .B2(G40), .ZN(new_n992));
  INV_X1    g567(.A(G40), .ZN(new_n993));
  NOR4_X1   g568(.A1(new_n467), .A2(new_n471), .A3(KEYINPUT113), .A4(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n489), .B2(new_n493), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n992), .A2(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n989), .B1(new_n990), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT124), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(G160), .A2(new_n991), .A3(G40), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n468), .A2(new_n470), .ZN(new_n1002));
  INV_X1    g577(.A(G125), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n473), .B2(new_n474), .ZN(new_n1004));
  INV_X1    g579(.A(new_n466), .ZN(new_n1005));
  OAI21_X1  g580(.A(G2105), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1006), .A3(G40), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT113), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n890), .A2(new_n891), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n889), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1001), .A2(new_n1008), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n883), .A2(new_n995), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT124), .A3(new_n989), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1000), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1001), .A2(new_n1008), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT112), .B(G1384), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n793), .A3(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1002), .A2(KEYINPUT125), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1006), .A2(KEYINPUT53), .A3(G40), .A4(new_n793), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1002), .A2(KEYINPUT125), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n883), .A2(new_n1021), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1018), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1017), .A2(new_n1023), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G301), .B1(new_n1016), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1023), .A2(new_n1017), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1018), .B1(new_n894), .B2(G1384), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1008), .A2(new_n1001), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT53), .A4(new_n793), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1033), .A2(G301), .A3(new_n998), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT54), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n990), .A2(new_n997), .A3(G2084), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1966), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n761), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT51), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n992), .A2(new_n994), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n883), .B2(new_n1009), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n763), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1012), .A2(new_n799), .A3(new_n1013), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1046), .B1(new_n1055), .B2(G8), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1048), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n995), .B1(new_n883), .B2(new_n1009), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n494), .A2(new_n995), .A3(new_n1009), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n992), .B2(new_n994), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1058), .A2(new_n1060), .A3(G2090), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1971), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G303), .A2(G8), .ZN(new_n1064));
  XOR2_X1   g639(.A(new_n1064), .B(KEYINPUT55), .Z(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n883), .B(new_n1009), .C1(new_n992), .C2(new_n994), .ZN(new_n1068));
  INV_X1    g643(.A(G288), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G1976), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(G8), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n499), .A2(G48), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(new_n584), .C1(new_n1075), .C2(new_n508), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(G1981), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n581), .A2(new_n583), .A3(new_n1079), .A4(new_n585), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1076), .B2(G1981), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1082), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(KEYINPUT49), .A3(new_n1080), .A4(new_n1078), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n892), .A2(new_n893), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1384), .B1(new_n1087), .B2(new_n493), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1008), .A2(new_n1001), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1083), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1976), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(G288), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1070), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1072), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1014), .A2(G2090), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1065), .B(G8), .C1(new_n1096), .C2(new_n1062), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1067), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1039), .A2(new_n1057), .A3(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT119), .B(G1996), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1019), .A2(new_n1022), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(G1341), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1068), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT59), .B1(new_n1105), .B2(new_n540), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1107), .B(new_n846), .C1(new_n1101), .C2(new_n1104), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1956), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1019), .A2(new_n1022), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n561), .B2(new_n566), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n561), .A2(new_n1116), .A3(new_n566), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n561), .A2(new_n1116), .A3(new_n566), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1121), .A2(new_n1117), .A3(KEYINPUT118), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1114), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1117), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(KEYINPUT61), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n609), .B(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n837), .B1(new_n990), .B2(new_n997), .ZN(new_n1129));
  INV_X1    g704(.A(G2067), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1088), .A2(new_n1089), .A3(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1348), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1088), .A2(new_n1130), .A3(new_n1089), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n609), .A2(KEYINPUT121), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1132), .B(new_n1136), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1124), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1111), .A2(new_n1113), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1109), .A2(new_n1126), .A3(new_n1139), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n609), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1125), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1146), .A2(new_n1123), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1023), .A2(new_n1017), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n998), .A2(new_n1036), .ZN(new_n1150));
  OAI21_X1  g725(.A(G171), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT123), .B(G171), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1016), .A2(G301), .A3(new_n1031), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1099), .A2(new_n1148), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1055), .A2(G8), .A3(new_n571), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(G8), .B1(new_n1096), .B2(new_n1062), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1066), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT117), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1166), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1168), .A2(new_n1164), .A3(new_n1162), .A4(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1098), .B2(new_n1160), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1167), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1098), .B1(new_n1154), .B2(new_n1153), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1057), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1048), .B(KEYINPUT62), .C1(new_n1050), .C2(new_n1056), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1097), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1091), .A2(new_n1092), .A3(new_n1069), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1080), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1179), .A2(new_n1095), .B1(new_n1181), .B2(new_n1090), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1159), .A2(new_n1173), .A3(new_n1178), .A4(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1029), .A2(new_n1018), .A3(new_n1089), .ZN(new_n1184));
  INV_X1    g759(.A(G1996), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n824), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n779), .B(G2067), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(G1996), .B2(new_n822), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1184), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT114), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n734), .B(new_n736), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1191), .B1(new_n1184), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1184), .ZN(new_n1194));
  XNOR2_X1  g769(.A(G290), .B(G1986), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1183), .A2(new_n1196), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1184), .A2(G1986), .A3(G290), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT48), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1193), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n736), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n734), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1191), .A2(new_n1202), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n779), .A2(G2067), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1184), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1194), .A2(new_n1185), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1206), .B(KEYINPUT46), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1187), .A2(new_n822), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1207), .B1(new_n1184), .B2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1209), .B(new_n1210), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1200), .A2(new_n1205), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1197), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g788(.A1(new_n682), .A2(G319), .A3(new_n683), .ZN(new_n1215));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g791(.A1(new_n682), .A2(KEYINPUT127), .A3(G319), .A4(new_n683), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AND4_X1   g793(.A1(new_n659), .A2(new_n712), .A3(new_n710), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n1220), .A2(new_n921), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n1221), .A2(new_n987), .ZN(G308));
  AND2_X1   g796(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1223));
  NOR3_X1   g797(.A1(new_n973), .A2(new_n975), .A3(KEYINPUT43), .ZN(new_n1224));
  OAI211_X1 g798(.A(new_n1220), .B(new_n921), .C1(new_n1223), .C2(new_n1224), .ZN(G225));
endmodule


