//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT77), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT77), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT3), .ZN(new_n196));
  AOI21_X1  g010(.A(G101), .B1(new_n188), .B2(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(KEYINPUT79), .A3(new_n196), .A4(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(G104), .B1(new_n191), .B2(new_n193), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n195), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT77), .B(G107), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n206), .A2(KEYINPUT81), .A3(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(G101), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT82), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n202), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n215), .B2(G116), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n213), .A3(G119), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT2), .B(G113), .Z(new_n220));
  AND2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(KEYINPUT5), .ZN(new_n222));
  INV_X1    g036(.A(G113), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT5), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n214), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n210), .A2(new_n212), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n188), .A2(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n194), .A2(new_n196), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G101), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(KEYINPUT80), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT78), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n235), .A3(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n202), .A2(new_n234), .A3(KEYINPUT4), .A4(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n219), .A2(new_n220), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n221), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n227), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G110), .B(G122), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT85), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n227), .A2(new_n241), .A3(new_n243), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n247), .A2(KEYINPUT6), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n249), .A3(new_n244), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n252), .A3(new_n244), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n242), .A2(KEYINPUT86), .A3(new_n252), .A4(new_n244), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G143), .B(G146), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G125), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT1), .B1(new_n260), .B2(G146), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n260), .A2(G146), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n258), .A2(G143), .ZN(new_n271));
  OAI211_X1 g085(.A(G128), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n259), .B(new_n261), .C1(KEYINPUT1), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n268), .B1(G125), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G224), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n251), .A2(new_n257), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n278), .A2(KEYINPUT7), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT87), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(KEYINPUT87), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n276), .B(new_n284), .Z(new_n285));
  XOR2_X1   g099(.A(new_n209), .B(new_n226), .Z(new_n286));
  XNOR2_X1  g100(.A(new_n243), .B(KEYINPUT8), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n283), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n288), .B2(new_n247), .ZN(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n280), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n280), .B2(new_n289), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n187), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G469), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT70), .B(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT12), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n298));
  INV_X1    g112(.A(new_n275), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n202), .A2(new_n208), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n209), .A2(new_n275), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n209), .A2(new_n301), .A3(new_n275), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(G137), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT11), .A3(G134), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(G137), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  INV_X1    g128(.A(G131), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n309), .A2(new_n311), .A3(new_n315), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n297), .B1(new_n306), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n297), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n298), .B(new_n319), .C1(new_n304), .C2(new_n305), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT10), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n275), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n210), .A2(new_n212), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n232), .A2(new_n237), .A3(new_n267), .ZN(new_n324));
  INV_X1    g138(.A(new_n317), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n300), .A2(new_n321), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G110), .B(G140), .ZN(new_n328));
  INV_X1    g142(.A(G227), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G953), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n318), .A2(new_n320), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n317), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n332), .B1(new_n336), .B2(new_n327), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n294), .B(new_n296), .C1(new_n334), .C2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n299), .B1(new_n202), .B2(new_n208), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n301), .B2(new_n300), .ZN(new_n340));
  INV_X1    g154(.A(new_n305), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT83), .B(new_n317), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n343));
  INV_X1    g157(.A(new_n319), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n306), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n327), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n331), .ZN(new_n347));
  INV_X1    g161(.A(new_n333), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n336), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(G469), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G902), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n294), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n338), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT9), .B(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(G221), .B1(new_n355), .B2(G902), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n293), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n359));
  INV_X1    g173(.A(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G125), .ZN(new_n361));
  INV_X1    g175(.A(G125), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G140), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n363), .A3(KEYINPUT16), .ZN(new_n364));
  OR3_X1    g178(.A1(new_n362), .A2(KEYINPUT16), .A3(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n258), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n365), .A3(G146), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n215), .A2(G128), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n215), .A2(G128), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT72), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n273), .A2(G119), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT72), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT24), .B(G110), .Z(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n273), .A2(KEYINPUT23), .A3(G119), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(new_n370), .C1(new_n372), .C2(KEYINPUT23), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT73), .B1(new_n380), .B2(G110), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n380), .A2(KEYINPUT73), .A3(G110), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n369), .B(new_n378), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G125), .B(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n258), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n377), .B1(new_n373), .B2(new_n376), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n380), .A2(G110), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n368), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n359), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT22), .B(G137), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n383), .A2(new_n359), .A3(new_n388), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n383), .A2(new_n393), .A3(new_n388), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(KEYINPUT75), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(KEYINPUT75), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n398), .A3(new_n296), .A4(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G234), .ZN(new_n404));
  OAI21_X1  g218(.A(G217), .B1(new_n295), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT71), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT75), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n397), .B(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n408), .A2(new_n296), .A3(new_n396), .A4(new_n401), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n408), .A2(new_n396), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n406), .A2(G902), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n308), .A2(G137), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n310), .A2(G134), .ZN(new_n417));
  OAI21_X1  g231(.A(G131), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n316), .A2(new_n418), .A3(KEYINPUT65), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT65), .B1(new_n316), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n299), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n317), .B2(new_n267), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n266), .B1(new_n314), .B2(new_n316), .ZN(new_n425));
  AND4_X1   g239(.A1(new_n316), .A2(new_n272), .A3(new_n274), .A4(new_n418), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n424), .A2(new_n240), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n429));
  INV_X1    g243(.A(G237), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n430), .A2(new_n277), .A3(G210), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT26), .B(G101), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n432), .B(new_n433), .Z(new_n434));
  INV_X1    g248(.A(new_n425), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n421), .A2(new_n435), .A3(new_n239), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT31), .B1(new_n428), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT67), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n240), .B1(new_n425), .B2(new_n426), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT28), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n316), .A2(new_n418), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n316), .A2(new_n418), .A3(KEYINPUT65), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n425), .B1(new_n446), .B2(new_n299), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n441), .B1(new_n447), .B2(new_n239), .ZN(new_n448));
  AND4_X1   g262(.A1(new_n441), .A2(new_n421), .A3(new_n435), .A4(new_n239), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n440), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n432), .B(new_n433), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n447), .B2(new_n239), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n424), .A2(new_n427), .A3(new_n240), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT31), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n439), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT31), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n454), .A2(new_n459), .A3(new_n434), .A4(new_n436), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n453), .A2(KEYINPUT68), .A3(new_n459), .A4(new_n454), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT69), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n459), .B1(new_n453), .B2(new_n454), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n451), .A2(new_n450), .B1(new_n466), .B2(new_n456), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n439), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(G472), .A2(G902), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT32), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G472), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n448), .A2(new_n449), .ZN(new_n477));
  INV_X1    g291(.A(new_n447), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n240), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT29), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n451), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n295), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n454), .A2(new_n436), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n451), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n484), .B(new_n480), .C1(new_n450), .C2(new_n451), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n476), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n472), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n465), .B2(new_n470), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT32), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n475), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G217), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n355), .A2(new_n495), .A3(G953), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G116), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n213), .A2(G122), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n206), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n260), .A2(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n273), .A2(G143), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G134), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n308), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n499), .B1(new_n500), .B2(KEYINPUT14), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n498), .A2(G116), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n501), .B(new_n507), .C1(new_n514), .C2(new_n190), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n191), .A2(new_n193), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n499), .A2(new_n500), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n501), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n506), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT13), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(G134), .C1(KEYINPUT13), .C2(new_n502), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n506), .A2(new_n520), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n519), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n515), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n526), .B1(new_n515), .B2(new_n525), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n497), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n515), .A2(new_n525), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT93), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n496), .A3(new_n527), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n533), .A3(new_n296), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT94), .A4(new_n296), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n494), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n493), .B1(new_n534), .B2(new_n535), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n277), .A2(G952), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n404), .B2(new_n430), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n277), .B(new_n296), .C1(G234), .C2(G237), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT21), .B(G898), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT20), .ZN(new_n548));
  NOR2_X1   g362(.A1(G475), .A2(G902), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n367), .A2(new_n368), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n430), .A2(new_n277), .A3(G214), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n260), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT17), .A3(G131), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(G131), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n551), .A2(new_n260), .ZN(new_n555));
  NOR2_X1   g369(.A1(G237), .A2(G953), .ZN(new_n556));
  AOI21_X1  g370(.A(G143), .B1(new_n556), .B2(G214), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n315), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n550), .B(new_n553), .C1(new_n560), .C2(KEYINPUT17), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n558), .B1(new_n562), .B2(new_n315), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n552), .A2(KEYINPUT18), .A3(G131), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n384), .A2(new_n258), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n565), .A2(KEYINPUT88), .A3(new_n385), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT88), .B1(new_n565), .B2(new_n385), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n563), .B(new_n564), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G113), .B(G122), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n188), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n561), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n384), .B1(KEYINPUT89), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n384), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n560), .B(new_n368), .C1(G146), .C2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n570), .B1(new_n576), .B2(new_n568), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n548), .B(new_n549), .C1(new_n571), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT90), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n561), .A2(new_n568), .A3(new_n570), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n576), .A2(new_n568), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n570), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT90), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n548), .A4(new_n549), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n549), .B1(new_n571), .B2(new_n577), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT20), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n579), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n570), .B1(new_n561), .B2(new_n568), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n351), .B1(new_n571), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G475), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n541), .A2(new_n547), .A3(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n358), .A2(new_n415), .A3(new_n491), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT95), .B(G101), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G3));
  INV_X1    g409(.A(new_n356), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n342), .A2(KEYINPUT12), .B1(new_n306), .B2(new_n344), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n348), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n336), .A2(new_n327), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n331), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n295), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n352), .B1(new_n601), .B2(new_n294), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n602), .B2(new_n350), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n471), .A2(new_n296), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n489), .B1(new_n604), .B2(G472), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n603), .A2(new_n605), .A3(KEYINPUT96), .A4(new_n415), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n354), .A2(new_n415), .A3(new_n356), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n295), .B1(new_n465), .B2(new_n470), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n473), .B1(new_n476), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n280), .A2(new_n289), .A3(KEYINPUT97), .A4(new_n290), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n187), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n291), .A2(new_n292), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n534), .A2(new_n492), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT33), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT33), .B1(new_n530), .B2(new_n533), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n296), .A2(G478), .ZN(new_n623));
  OAI211_X1 g437(.A(KEYINPUT98), .B(new_n618), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n530), .A2(new_n533), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n623), .B1(new_n628), .B2(new_n619), .ZN(new_n629));
  INV_X1    g443(.A(new_n618), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n587), .A2(new_n590), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n547), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n617), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n612), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NAND2_X1  g454(.A1(new_n280), .A2(new_n289), .ZN(new_n641));
  INV_X1    g455(.A(new_n290), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n280), .A2(new_n289), .A3(new_n290), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n616), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n613), .A2(new_n187), .ZN(new_n646));
  INV_X1    g460(.A(new_n547), .ZN(new_n647));
  INV_X1    g461(.A(new_n586), .ZN(new_n648));
  INV_X1    g462(.A(new_n578), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n647), .B(new_n590), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n645), .A2(new_n646), .A3(new_n541), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n612), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  INV_X1    g470(.A(new_n395), .ZN(new_n657));
  OAI22_X1  g471(.A1(new_n657), .A2(new_n389), .B1(KEYINPUT36), .B2(new_n394), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n394), .A2(KEYINPUT36), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n390), .A2(new_n395), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n656), .B1(new_n661), .B2(new_n412), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n661), .A2(new_n656), .A3(new_n412), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n410), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n410), .A2(KEYINPUT100), .A3(new_n663), .A4(new_n664), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n592), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n358), .A2(new_n605), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND4_X1  g486(.A1(new_n354), .A2(new_n667), .A3(new_n356), .A4(new_n668), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT101), .B(G900), .Z(new_n675));
  AOI21_X1  g489(.A(new_n544), .B1(new_n545), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n590), .B(new_n677), .C1(new_n648), .C2(new_n649), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n540), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n617), .A2(new_n674), .A3(new_n491), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XOR2_X1   g495(.A(new_n676), .B(KEYINPUT39), .Z(new_n682));
  AND2_X1   g496(.A1(new_n603), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n478), .A2(new_n240), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n434), .B1(new_n685), .B2(new_n436), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n455), .B1(new_n686), .B2(KEYINPUT102), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n351), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G472), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n475), .A2(new_n490), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n615), .A2(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n291), .B2(new_n292), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n541), .A2(new_n187), .A3(new_n591), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n695), .A2(new_n665), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n684), .A2(new_n691), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND4_X1  g513(.A1(new_n591), .A2(new_n624), .A3(new_n631), .A4(new_n677), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n617), .A2(new_n674), .A3(new_n491), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NAND2_X1  g517(.A1(KEYINPUT103), .A2(G469), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n337), .B1(new_n597), .B2(new_n348), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n705), .B1(new_n706), .B2(new_n295), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n598), .A2(new_n600), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n296), .A3(new_n704), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n709), .A3(new_n356), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n707), .A2(new_n709), .A3(KEYINPUT104), .A4(new_n356), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n491), .A2(new_n415), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n637), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NOR2_X1   g531(.A1(new_n714), .A2(new_n652), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n213), .ZN(G18));
  AND3_X1   g533(.A1(new_n707), .A2(new_n356), .A3(new_n709), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n617), .A2(new_n491), .A3(new_n669), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND3_X1  g536(.A1(new_n712), .A2(new_n647), .A3(new_n713), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n645), .A2(new_n646), .A3(new_n541), .A4(new_n591), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n438), .B1(new_n479), .B2(new_n434), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n472), .B1(new_n725), .B2(new_n464), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n415), .B(new_n726), .C1(new_n609), .C2(new_n476), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n723), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n498), .ZN(G24));
  NAND3_X1  g543(.A1(new_n645), .A2(new_n720), .A3(new_n646), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n604), .A2(G472), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n701), .A3(new_n665), .A4(new_n726), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT105), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n665), .B(new_n726), .C1(new_n609), .C2(new_n476), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n700), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n617), .A2(new_n735), .A3(new_n736), .A4(new_n720), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT106), .B(G125), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G27));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n347), .A2(new_n741), .A3(G469), .A4(new_n349), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n338), .A3(new_n353), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n346), .A2(new_n331), .B1(new_n348), .B2(new_n336), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n741), .B1(new_n744), .B2(G469), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n356), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n643), .A2(new_n187), .A3(new_n644), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT108), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n187), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n291), .A2(new_n292), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n350), .A2(KEYINPUT107), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n602), .A2(new_n752), .A3(new_n742), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n750), .A2(new_n751), .A3(new_n356), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n491), .A2(new_n415), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n757), .A3(new_n701), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n756), .B1(new_n748), .B2(new_n754), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT109), .B(G131), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G33));
  NAND3_X1  g579(.A1(new_n755), .A2(new_n757), .A3(new_n679), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  INV_X1    g581(.A(new_n338), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n347), .A2(new_n349), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n744), .A2(KEYINPUT45), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(G469), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n353), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n768), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n353), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n596), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n633), .A2(new_n624), .A3(new_n631), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT43), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n610), .A3(new_n665), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n779), .A2(new_n682), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n750), .B1(new_n787), .B2(new_n788), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n310), .ZN(G39));
  NOR4_X1   g609(.A1(new_n491), .A2(new_n747), .A3(new_n415), .A4(new_n700), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n776), .A2(new_n777), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n356), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n800), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n778), .B2(new_n596), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n798), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT114), .B(G140), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G42));
  NOR2_X1   g620(.A1(G952), .A2(G953), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n489), .A2(KEYINPUT32), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n474), .B(new_n488), .C1(new_n465), .C2(new_n470), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n810), .A3(new_n486), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n536), .A2(new_n537), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n493), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  INV_X1    g628(.A(new_n539), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT116), .B1(new_n538), .B2(new_n539), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n678), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n643), .A2(new_n818), .A3(new_n187), .A4(new_n644), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n811), .A2(new_n673), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n755), .B2(new_n735), .ZN(new_n821));
  AND4_X1   g635(.A1(KEYINPUT42), .A2(new_n755), .A3(new_n757), .A4(new_n701), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT42), .B1(new_n761), .B2(new_n701), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n766), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n612), .A2(new_n293), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n816), .A2(new_n817), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n547), .A3(new_n591), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n636), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n714), .B1(new_n637), .B2(new_n652), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n728), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n593), .A2(new_n721), .A3(new_n670), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n824), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n742), .A2(new_n338), .A3(new_n353), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n596), .B1(new_n835), .B2(new_n752), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n665), .A2(new_n676), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n691), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n680), .B(new_n702), .C1(new_n724), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n733), .A2(new_n737), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT52), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n645), .A2(new_n646), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n673), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n843), .B(new_n491), .C1(new_n679), .C2(new_n701), .ZN(new_n844));
  INV_X1    g658(.A(new_n724), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n691), .A3(new_n836), .A4(new_n837), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n738), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n834), .A2(KEYINPUT53), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n831), .A2(new_n829), .A3(new_n728), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n821), .A2(new_n766), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n763), .A2(new_n852), .A3(new_n853), .A4(new_n828), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n667), .A2(new_n668), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n603), .A3(new_n645), .A4(new_n646), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n491), .A2(new_n679), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n491), .A2(new_n701), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n838), .A2(new_n724), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n847), .B1(new_n861), .B2(new_n738), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n847), .A2(new_n844), .A3(new_n738), .A4(new_n846), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT117), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n841), .A2(new_n865), .A3(new_n848), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n854), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n808), .B(new_n851), .C1(new_n867), .C2(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT118), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n841), .A2(new_n865), .A3(new_n848), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n865), .B1(new_n841), .B2(new_n848), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n834), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n808), .A4(new_n851), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n834), .B(KEYINPUT53), .C1(new_n870), .C2(new_n871), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n854), .B2(new_n849), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT54), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n747), .A2(new_n710), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n786), .A2(new_n544), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n756), .ZN(new_n883));
  XNOR2_X1  g697(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n691), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n881), .A3(new_n415), .A4(new_n544), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(new_n635), .ZN(new_n888));
  INV_X1    g702(.A(new_n727), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n544), .A2(new_n889), .A3(new_n784), .A4(new_n785), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n617), .A3(new_n720), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n885), .A2(new_n542), .A3(new_n888), .A4(new_n891), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n187), .B(new_n710), .C1(new_n692), .C2(new_n694), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n893), .A2(KEYINPUT50), .A3(new_n890), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT50), .B1(new_n893), .B2(new_n890), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n632), .A2(new_n633), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n882), .A2(new_n734), .B1(new_n887), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT119), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n890), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n747), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n707), .A2(new_n709), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n356), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n803), .B2(new_n801), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g720(.A(KEYINPUT120), .B(new_n903), .C1(new_n803), .C2(new_n801), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT51), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n896), .A2(new_n898), .ZN(new_n910));
  NAND2_X1  g724(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n911));
  OR3_X1    g725(.A1(new_n900), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n910), .B(new_n911), .C1(new_n904), .C2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n892), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n869), .A2(new_n876), .A3(new_n880), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n807), .B1(new_n915), .B2(KEYINPUT122), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n808), .B1(new_n877), .B2(new_n878), .ZN(new_n917));
  INV_X1    g731(.A(new_n868), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n875), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n869), .A4(new_n914), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n414), .A2(new_n596), .A3(new_n749), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT115), .ZN(new_n924));
  INV_X1    g738(.A(new_n780), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(new_n925), .C1(KEYINPUT49), .C2(new_n902), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(KEYINPUT49), .B2(new_n902), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n886), .A3(new_n695), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n922), .A2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n277), .A2(G952), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n874), .A2(new_n851), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n295), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n935), .B2(new_n290), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n251), .A2(new_n257), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n279), .Z(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT55), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n933), .B(new_n939), .C1(new_n935), .C2(new_n290), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n932), .B1(new_n941), .B2(new_n942), .ZN(G51));
  NAND2_X1  g757(.A1(new_n864), .A2(new_n866), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n944), .B2(new_n834), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n854), .A2(new_n873), .A3(new_n849), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n808), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n918), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n352), .B(KEYINPUT57), .Z(new_n950));
  OAI21_X1  g764(.A(new_n708), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n935), .A2(new_n773), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n930), .B1(new_n951), .B2(new_n952), .ZN(G54));
  NAND2_X1  g767(.A1(KEYINPUT58), .A2(G475), .ZN(new_n954));
  OAI221_X1 g768(.A(new_n580), .B1(new_n570), .B2(new_n581), .C1(new_n935), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n935), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n956), .A2(KEYINPUT58), .A3(G475), .A4(new_n582), .ZN(new_n957));
  INV_X1    g771(.A(new_n930), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(G60));
  XOR2_X1   g773(.A(new_n622), .B(KEYINPUT124), .Z(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT59), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n931), .B1(new_n949), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n869), .A2(new_n876), .A3(new_n880), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n960), .B1(new_n965), .B2(new_n962), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n934), .A2(new_n661), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n947), .A2(new_n969), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n931), .B(new_n971), .C1(new_n972), .C2(new_n411), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G66));
  INV_X1    g789(.A(new_n546), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n277), .B1(new_n976), .B2(G224), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n833), .B2(new_n277), .ZN(new_n978));
  INV_X1    g792(.A(G898), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n937), .B1(new_n979), .B2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G69));
  NOR2_X1   g795(.A1(new_n277), .A2(G900), .ZN(new_n982));
  INV_X1    g796(.A(new_n794), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n779), .A2(new_n757), .A3(new_n682), .A4(new_n845), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n840), .A2(new_n859), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(new_n766), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n983), .A2(new_n763), .A3(new_n804), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n988), .B2(new_n277), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  INV_X1    g805(.A(new_n804), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n794), .A2(new_n986), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(G953), .B1(new_n993), .B2(new_n763), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n991), .B1(new_n994), .B2(new_n982), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n424), .A2(new_n427), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(new_n575), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n985), .A2(new_n698), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT62), .Z(new_n1001));
  OAI21_X1  g815(.A(new_n635), .B1(new_n826), .B2(new_n591), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n750), .B1(new_n1003), .B2(KEYINPUT125), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(KEYINPUT125), .B2(new_n1003), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n757), .A3(new_n683), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1001), .A2(new_n983), .A3(new_n804), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n998), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1007), .A2(new_n277), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n982), .B1(new_n329), .B2(G953), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n999), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1008), .B1(new_n990), .B2(new_n995), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1009), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1012), .A2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n1007), .B2(new_n833), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n483), .B(KEYINPUT127), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1019), .A2(new_n434), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1018), .B1(new_n988), .B2(new_n833), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1020), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1022), .A2(new_n451), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1021), .A2(new_n958), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1018), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n484), .B2(new_n455), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1025), .B1(new_n879), .B2(new_n1027), .ZN(G57));
endmodule


