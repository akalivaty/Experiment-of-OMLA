

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(n717), .A2(KEYINPUT33), .ZN(n719) );
  NOR2_X1 U553 ( .A1(n727), .A2(n636), .ZN(n637) );
  NOR2_X1 U554 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U555 ( .A1(n739), .A2(G1966), .ZN(n635) );
  NAND2_X1 U556 ( .A1(n634), .A2(n633), .ZN(n693) );
  INV_X1 U557 ( .A(KEYINPUT99), .ZN(n718) );
  AND2_X1 U558 ( .A1(n651), .A2(n650), .ZN(n652) );
  INV_X1 U559 ( .A(KEYINPUT40), .ZN(n754) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n535), .Z(n796) );
  XNOR2_X1 U561 ( .A(n754), .B(KEYINPUT106), .ZN(n755) );
  XNOR2_X1 U562 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n516) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  XNOR2_X2 U564 ( .A(n516), .B(n515), .ZN(n887) );
  NAND2_X1 U565 ( .A1(G138), .A2(n887), .ZN(n518) );
  INV_X1 U566 ( .A(G2105), .ZN(n519) );
  AND2_X1 U567 ( .A1(n519), .A2(G2104), .ZN(n886) );
  NAND2_X1 U568 ( .A1(G102), .A2(n886), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n518), .A2(n517), .ZN(n523) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U571 ( .A1(G114), .A2(n881), .ZN(n521) );
  NOR2_X1 U572 ( .A1(G2104), .A2(n519), .ZN(n882) );
  NAND2_X1 U573 ( .A1(G126), .A2(n882), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U575 ( .A1(n523), .A2(n522), .ZN(G164) );
  NAND2_X1 U576 ( .A1(n887), .A2(G137), .ZN(n526) );
  NAND2_X1 U577 ( .A1(G101), .A2(n886), .ZN(n524) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n524), .Z(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n530) );
  NAND2_X1 U580 ( .A1(G113), .A2(n881), .ZN(n528) );
  NAND2_X1 U581 ( .A1(G125), .A2(n882), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U583 ( .A1(n530), .A2(n529), .ZN(G160) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n791) );
  NAND2_X1 U585 ( .A1(n791), .A2(G85), .ZN(n532) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n573) );
  XOR2_X1 U587 ( .A(G651), .B(KEYINPUT66), .Z(n534) );
  NOR2_X1 U588 ( .A1(n573), .A2(n534), .ZN(n792) );
  NAND2_X1 U589 ( .A1(n792), .A2(G72), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U591 ( .A(KEYINPUT67), .B(n533), .Z(n538) );
  NOR2_X1 U592 ( .A1(G543), .A2(n534), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n796), .A2(G60), .ZN(n536) );
  XOR2_X1 U594 ( .A(KEYINPUT68), .B(n536), .Z(n537) );
  NOR2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n541) );
  NOR2_X1 U596 ( .A1(G651), .A2(n573), .ZN(n539) );
  XNOR2_X1 U597 ( .A(KEYINPUT64), .B(n539), .ZN(n799) );
  NAND2_X1 U598 ( .A1(G47), .A2(n799), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(G290) );
  NAND2_X1 U600 ( .A1(n791), .A2(G89), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G76), .A2(n792), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U604 ( .A(n545), .B(KEYINPUT5), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G63), .A2(n796), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G51), .A2(n799), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n548), .Z(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n551), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U611 ( .A1(G90), .A2(n791), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G77), .A2(n792), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U614 ( .A(KEYINPUT9), .B(n554), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n799), .A2(G52), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G64), .A2(n796), .ZN(n555) );
  AND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(G301) );
  INV_X1 U619 ( .A(G301), .ZN(G171) );
  NAND2_X1 U620 ( .A1(n799), .A2(G53), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT70), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G65), .A2(n796), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G91), .A2(n791), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G78), .A2(n792), .ZN(n562) );
  XNOR2_X1 U626 ( .A(KEYINPUT69), .B(n562), .ZN(n563) );
  NOR2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(G299) );
  NAND2_X1 U629 ( .A1(G88), .A2(n791), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G75), .A2(n792), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G62), .A2(n796), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G50), .A2(n799), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n572), .A2(n571), .ZN(G166) );
  INV_X1 U636 ( .A(G166), .ZN(G303) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(n573), .A2(G87), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G49), .A2(n799), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n796), .A2(n576), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G651), .A2(G74), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U644 ( .A1(G61), .A2(n796), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G86), .A2(n791), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G73), .A2(n792), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT2), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n582), .B(KEYINPUT77), .ZN(n583) );
  NOR2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G48), .A2(n799), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(G305) );
  XNOR2_X1 U653 ( .A(G2067), .B(KEYINPUT37), .ZN(n596) );
  NAND2_X1 U654 ( .A1(G104), .A2(n886), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G140), .A2(n887), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U657 ( .A(KEYINPUT34), .B(n589), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G116), .A2(n881), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G128), .A2(n882), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U661 ( .A(KEYINPUT35), .B(n592), .Z(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U663 ( .A(KEYINPUT36), .B(n595), .ZN(n895) );
  NAND2_X1 U664 ( .A1(n596), .A2(n895), .ZN(n964) );
  NOR2_X1 U665 ( .A1(n596), .A2(n895), .ZN(n947) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n634) );
  AND2_X1 U667 ( .A1(G160), .A2(G40), .ZN(n633) );
  INV_X1 U668 ( .A(n633), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n634), .A2(n597), .ZN(n746) );
  NAND2_X1 U670 ( .A1(n947), .A2(n746), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT82), .ZN(n743) );
  XNOR2_X1 U672 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n627) );
  NAND2_X1 U673 ( .A1(n887), .A2(G141), .ZN(n606) );
  XOR2_X1 U674 ( .A(KEYINPUT38), .B(KEYINPUT86), .Z(n600) );
  NAND2_X1 U675 ( .A1(G105), .A2(n886), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n600), .B(n599), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G117), .A2(n881), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G129), .A2(n882), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U682 ( .A(KEYINPUT87), .B(n607), .Z(n869) );
  NOR2_X1 U683 ( .A1(G1996), .A2(n869), .ZN(n952) );
  NAND2_X1 U684 ( .A1(G1996), .A2(n869), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G107), .A2(n881), .ZN(n609) );
  NAND2_X1 U686 ( .A1(G119), .A2(n882), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G95), .A2(n886), .ZN(n611) );
  NAND2_X1 U689 ( .A1(G131), .A2(n887), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U691 ( .A(KEYINPUT83), .B(n612), .Z(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U693 ( .A(KEYINPUT84), .B(n615), .Z(n899) );
  NAND2_X1 U694 ( .A1(G1991), .A2(n899), .ZN(n616) );
  XOR2_X1 U695 ( .A(KEYINPUT85), .B(n616), .Z(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT88), .B(n619), .Z(n949) );
  INV_X1 U698 ( .A(n949), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n620), .A2(n746), .ZN(n749) );
  INV_X1 U700 ( .A(n749), .ZN(n624) );
  NOR2_X1 U701 ( .A1(G1986), .A2(G290), .ZN(n622) );
  NOR2_X1 U702 ( .A1(n899), .A2(G1991), .ZN(n621) );
  XNOR2_X1 U703 ( .A(n621), .B(KEYINPUT102), .ZN(n944) );
  NOR2_X1 U704 ( .A1(n622), .A2(n944), .ZN(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n952), .A2(n625), .ZN(n626) );
  XOR2_X1 U707 ( .A(n627), .B(n626), .Z(n628) );
  NAND2_X1 U708 ( .A1(n743), .A2(n628), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n964), .A2(n629), .ZN(n630) );
  XNOR2_X1 U710 ( .A(KEYINPUT104), .B(n630), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n631), .A2(n746), .ZN(n632) );
  XNOR2_X1 U712 ( .A(KEYINPUT105), .B(n632), .ZN(n753) );
  NAND2_X1 U713 ( .A1(G8), .A2(n693), .ZN(n739) );
  NOR2_X1 U714 ( .A1(G2084), .A2(n693), .ZN(n727) );
  XNOR2_X1 U715 ( .A(n635), .B(KEYINPUT89), .ZN(n709) );
  NAND2_X1 U716 ( .A1(G8), .A2(n709), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT30), .B(n637), .Z(n638) );
  NOR2_X1 U718 ( .A1(G168), .A2(n638), .ZN(n643) );
  XOR2_X1 U719 ( .A(KEYINPUT25), .B(G2078), .Z(n1001) );
  NOR2_X1 U720 ( .A1(n1001), .A2(n693), .ZN(n639) );
  XNOR2_X1 U721 ( .A(n639), .B(KEYINPUT91), .ZN(n641) );
  XOR2_X1 U722 ( .A(G1961), .B(KEYINPUT90), .Z(n914) );
  NAND2_X1 U723 ( .A1(n914), .A2(n693), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n646) );
  NOR2_X1 U725 ( .A1(G171), .A2(n646), .ZN(n642) );
  XOR2_X1 U726 ( .A(n644), .B(KEYINPUT98), .Z(n645) );
  XNOR2_X1 U727 ( .A(n645), .B(KEYINPUT31), .ZN(n707) );
  NAND2_X1 U728 ( .A1(n646), .A2(G171), .ZN(n692) );
  XNOR2_X1 U729 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n690) );
  NAND2_X1 U730 ( .A1(n796), .A2(G66), .ZN(n647) );
  XNOR2_X1 U731 ( .A(KEYINPUT72), .B(n647), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n799), .A2(G54), .ZN(n651) );
  NAND2_X1 U733 ( .A1(G92), .A2(n791), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G79), .A2(n792), .ZN(n648) );
  AND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n654), .B(KEYINPUT15), .ZN(n977) );
  NAND2_X1 U738 ( .A1(n796), .A2(G56), .ZN(n655) );
  XOR2_X1 U739 ( .A(KEYINPUT14), .B(n655), .Z(n661) );
  NAND2_X1 U740 ( .A1(n791), .A2(G81), .ZN(n656) );
  XNOR2_X1 U741 ( .A(n656), .B(KEYINPUT12), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G68), .A2(n792), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U744 ( .A(KEYINPUT13), .B(n659), .Z(n660) );
  NOR2_X1 U745 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U746 ( .A1(G43), .A2(n799), .ZN(n662) );
  NAND2_X1 U747 ( .A1(n663), .A2(n662), .ZN(n978) );
  INV_X1 U748 ( .A(n693), .ZN(n679) );
  AND2_X1 U749 ( .A1(n679), .A2(G1996), .ZN(n665) );
  XOR2_X1 U750 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n664) );
  XNOR2_X1 U751 ( .A(n665), .B(n664), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n693), .A2(G1341), .ZN(n666) );
  NAND2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U754 ( .A1(n978), .A2(n668), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n977), .A2(n675), .ZN(n673) );
  AND2_X1 U756 ( .A1(n679), .A2(G2067), .ZN(n669) );
  XNOR2_X1 U757 ( .A(n669), .B(KEYINPUT95), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n693), .A2(G1348), .ZN(n670) );
  NAND2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U760 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U761 ( .A(n674), .B(KEYINPUT96), .ZN(n677) );
  OR2_X1 U762 ( .A1(n675), .A2(n977), .ZN(n676) );
  NAND2_X1 U763 ( .A1(n677), .A2(n676), .ZN(n683) );
  INV_X1 U764 ( .A(G299), .ZN(n970) );
  NAND2_X1 U765 ( .A1(n679), .A2(G2072), .ZN(n678) );
  XNOR2_X1 U766 ( .A(n678), .B(KEYINPUT27), .ZN(n681) );
  XOR2_X1 U767 ( .A(G1956), .B(KEYINPUT92), .Z(n926) );
  NOR2_X1 U768 ( .A1(n679), .A2(n926), .ZN(n680) );
  NOR2_X1 U769 ( .A1(n681), .A2(n680), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n970), .A2(n684), .ZN(n682) );
  NAND2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n688) );
  NOR2_X1 U772 ( .A1(n970), .A2(n684), .ZN(n686) );
  XNOR2_X1 U773 ( .A(KEYINPUT93), .B(KEYINPUT28), .ZN(n685) );
  XNOR2_X1 U774 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n706) );
  INV_X1 U778 ( .A(G8), .ZN(n698) );
  NOR2_X1 U779 ( .A1(G1971), .A2(n739), .ZN(n695) );
  NOR2_X1 U780 ( .A1(G2090), .A2(n693), .ZN(n694) );
  NOR2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U782 ( .A1(n696), .A2(G303), .ZN(n697) );
  OR2_X1 U783 ( .A1(n698), .A2(n697), .ZN(n700) );
  AND2_X1 U784 ( .A1(n706), .A2(n700), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n707), .A2(n699), .ZN(n704) );
  INV_X1 U786 ( .A(n700), .ZN(n702) );
  AND2_X1 U787 ( .A1(G286), .A2(G8), .ZN(n701) );
  OR2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U789 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U790 ( .A(n705), .B(KEYINPUT32), .ZN(n730) );
  NAND2_X1 U791 ( .A1(n707), .A2(n706), .ZN(n708) );
  AND2_X1 U792 ( .A1(n709), .A2(n708), .ZN(n728) );
  INV_X1 U793 ( .A(n728), .ZN(n710) );
  NAND2_X1 U794 ( .A1(G1976), .A2(G288), .ZN(n969) );
  AND2_X1 U795 ( .A1(n710), .A2(n969), .ZN(n711) );
  NAND2_X1 U796 ( .A1(n730), .A2(n711), .ZN(n715) );
  INV_X1 U797 ( .A(n969), .ZN(n713) );
  NOR2_X1 U798 ( .A1(G1976), .A2(G288), .ZN(n720) );
  NOR2_X1 U799 ( .A1(G1971), .A2(G303), .ZN(n712) );
  NOR2_X1 U800 ( .A1(n720), .A2(n712), .ZN(n976) );
  OR2_X1 U801 ( .A1(n713), .A2(n976), .ZN(n714) );
  AND2_X1 U802 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U803 ( .A1(n739), .A2(n716), .ZN(n717) );
  XNOR2_X1 U804 ( .A(n719), .B(n718), .ZN(n726) );
  XNOR2_X1 U805 ( .A(G1981), .B(G305), .ZN(n986) );
  NAND2_X1 U806 ( .A1(n720), .A2(KEYINPUT33), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n721), .A2(n739), .ZN(n722) );
  XNOR2_X1 U808 ( .A(KEYINPUT100), .B(n722), .ZN(n723) );
  NOR2_X1 U809 ( .A1(n986), .A2(n723), .ZN(n724) );
  AND2_X1 U810 ( .A1(n724), .A2(n743), .ZN(n725) );
  NAND2_X1 U811 ( .A1(n726), .A2(n725), .ZN(n745) );
  NAND2_X1 U812 ( .A1(G8), .A2(n727), .ZN(n729) );
  NAND2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U814 ( .A1(n731), .A2(n730), .ZN(n734) );
  NOR2_X1 U815 ( .A1(G2090), .A2(G303), .ZN(n732) );
  NAND2_X1 U816 ( .A1(G8), .A2(n732), .ZN(n733) );
  NAND2_X1 U817 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U818 ( .A1(n739), .A2(n735), .ZN(n736) );
  XOR2_X1 U819 ( .A(KEYINPUT101), .B(n736), .Z(n741) );
  NOR2_X1 U820 ( .A1(G1981), .A2(G305), .ZN(n737) );
  XOR2_X1 U821 ( .A(n737), .B(KEYINPUT24), .Z(n738) );
  OR2_X1 U822 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U823 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U824 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U825 ( .A1(n745), .A2(n744), .ZN(n751) );
  XNOR2_X1 U826 ( .A(G1986), .B(G290), .ZN(n980) );
  NAND2_X1 U827 ( .A1(n980), .A2(n746), .ZN(n747) );
  XOR2_X1 U828 ( .A(n747), .B(KEYINPUT81), .Z(n748) );
  NAND2_X1 U829 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U830 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U831 ( .A1(n753), .A2(n752), .ZN(n756) );
  XNOR2_X1 U832 ( .A(n756), .B(n755), .ZN(G329) );
  XOR2_X1 U833 ( .A(G2446), .B(G2451), .Z(n758) );
  XNOR2_X1 U834 ( .A(G2454), .B(KEYINPUT107), .ZN(n757) );
  XNOR2_X1 U835 ( .A(n758), .B(n757), .ZN(n765) );
  XOR2_X1 U836 ( .A(G2438), .B(G2430), .Z(n760) );
  XNOR2_X1 U837 ( .A(G2435), .B(G2443), .ZN(n759) );
  XNOR2_X1 U838 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U839 ( .A(n761), .B(G2427), .Z(n763) );
  XNOR2_X1 U840 ( .A(G1341), .B(G1348), .ZN(n762) );
  XNOR2_X1 U841 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U842 ( .A(n765), .B(n764), .ZN(n766) );
  AND2_X1 U843 ( .A1(n766), .A2(G14), .ZN(G401) );
  AND2_X1 U844 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U845 ( .A1(n881), .A2(G111), .ZN(n773) );
  NAND2_X1 U846 ( .A1(G99), .A2(n886), .ZN(n768) );
  NAND2_X1 U847 ( .A1(G135), .A2(n887), .ZN(n767) );
  NAND2_X1 U848 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U849 ( .A1(n882), .A2(G123), .ZN(n769) );
  XOR2_X1 U850 ( .A(KEYINPUT18), .B(n769), .Z(n770) );
  NOR2_X1 U851 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U852 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U853 ( .A(KEYINPUT73), .B(n774), .Z(n941) );
  XNOR2_X1 U854 ( .A(G2096), .B(n941), .ZN(n775) );
  OR2_X1 U855 ( .A1(G2100), .A2(n775), .ZN(G156) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  INV_X1 U858 ( .A(G120), .ZN(G236) );
  INV_X1 U859 ( .A(G69), .ZN(G235) );
  INV_X1 U860 ( .A(G57), .ZN(G237) );
  XOR2_X1 U861 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n777) );
  NAND2_X1 U862 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U863 ( .A(n777), .B(n776), .ZN(G223) );
  INV_X1 U864 ( .A(G223), .ZN(n831) );
  NAND2_X1 U865 ( .A1(n831), .A2(G567), .ZN(n778) );
  XOR2_X1 U866 ( .A(KEYINPUT11), .B(n778), .Z(G234) );
  INV_X1 U867 ( .A(G860), .ZN(n783) );
  OR2_X1 U868 ( .A1(n978), .A2(n783), .ZN(G153) );
  NAND2_X1 U869 ( .A1(G868), .A2(G301), .ZN(n780) );
  OR2_X1 U870 ( .A1(n977), .A2(G868), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(G284) );
  INV_X1 U872 ( .A(G868), .ZN(n811) );
  NOR2_X1 U873 ( .A1(G286), .A2(n811), .ZN(n782) );
  NOR2_X1 U874 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U875 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U876 ( .A1(n783), .A2(G559), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n784), .A2(n977), .ZN(n785) );
  XNOR2_X1 U878 ( .A(n785), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U879 ( .A1(G868), .A2(n978), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G868), .A2(n977), .ZN(n786) );
  NOR2_X1 U881 ( .A1(G559), .A2(n786), .ZN(n787) );
  NOR2_X1 U882 ( .A1(n788), .A2(n787), .ZN(G282) );
  XNOR2_X1 U883 ( .A(n978), .B(KEYINPUT74), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n977), .A2(G559), .ZN(n789) );
  XNOR2_X1 U885 ( .A(n790), .B(n789), .ZN(n809) );
  NOR2_X1 U886 ( .A1(G860), .A2(n809), .ZN(n803) );
  NAND2_X1 U887 ( .A1(G93), .A2(n791), .ZN(n794) );
  NAND2_X1 U888 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U890 ( .A(n795), .B(KEYINPUT75), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G67), .A2(n796), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n799), .A2(G55), .ZN(n800) );
  XOR2_X1 U894 ( .A(KEYINPUT76), .B(n800), .Z(n801) );
  OR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n812) );
  XOR2_X1 U896 ( .A(n803), .B(n812), .Z(G145) );
  XNOR2_X1 U897 ( .A(KEYINPUT19), .B(G290), .ZN(n804) );
  XNOR2_X1 U898 ( .A(n804), .B(G288), .ZN(n805) );
  XOR2_X1 U899 ( .A(n812), .B(n805), .Z(n807) );
  XNOR2_X1 U900 ( .A(G305), .B(G166), .ZN(n806) );
  XNOR2_X1 U901 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(G299), .ZN(n903) );
  XOR2_X1 U903 ( .A(n903), .B(n809), .Z(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n814) );
  NOR2_X1 U905 ( .A1(G868), .A2(n812), .ZN(n813) );
  NOR2_X1 U906 ( .A1(n814), .A2(n813), .ZN(G295) );
  XOR2_X1 U907 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n816) );
  NAND2_X1 U908 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U911 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U914 ( .A(G661), .ZN(n830) );
  NOR2_X1 U915 ( .A1(G235), .A2(G236), .ZN(n820) );
  XNOR2_X1 U916 ( .A(n820), .B(KEYINPUT79), .ZN(n821) );
  NOR2_X1 U917 ( .A1(G237), .A2(n821), .ZN(n822) );
  NAND2_X1 U918 ( .A1(G108), .A2(n822), .ZN(n838) );
  NAND2_X1 U919 ( .A1(G567), .A2(n838), .ZN(n827) );
  NOR2_X1 U920 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U922 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U923 ( .A1(G96), .A2(n825), .ZN(n839) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n839), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U926 ( .A(KEYINPUT80), .B(n828), .Z(n859) );
  NAND2_X1 U927 ( .A1(G483), .A2(n859), .ZN(n829) );
  NOR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(n831), .A2(G2106), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n832), .B(KEYINPUT108), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n833) );
  XNOR2_X1 U933 ( .A(KEYINPUT109), .B(n833), .ZN(n834) );
  NAND2_X1 U934 ( .A1(n834), .A2(G661), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n835) );
  XNOR2_X1 U936 ( .A(KEYINPUT110), .B(n835), .ZN(n837) );
  NAND2_X1 U937 ( .A1(n837), .A2(n836), .ZN(G188) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G325) );
  XNOR2_X1 U939 ( .A(KEYINPUT111), .B(G325), .ZN(G261) );
  XNOR2_X1 U940 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  XOR2_X1 U943 ( .A(KEYINPUT113), .B(G2090), .Z(n841) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2084), .ZN(n840) );
  XNOR2_X1 U945 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U946 ( .A(n842), .B(G2096), .Z(n844) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2072), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2678), .Z(n846) );
  XNOR2_X1 U950 ( .A(G2100), .B(KEYINPUT42), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U952 ( .A(n848), .B(n847), .Z(G227) );
  XNOR2_X1 U953 ( .A(G1996), .B(G2474), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1956), .B(G1961), .Z(n850) );
  XNOR2_X1 U955 ( .A(G1991), .B(G1981), .ZN(n849) );
  XNOR2_X1 U956 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U957 ( .A(G1966), .B(G1971), .Z(n852) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1976), .ZN(n851) );
  XNOR2_X1 U959 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U960 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U961 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U962 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U963 ( .A(n858), .B(n857), .ZN(G229) );
  XNOR2_X1 U964 ( .A(KEYINPUT112), .B(n859), .ZN(G319) );
  NAND2_X1 U965 ( .A1(G100), .A2(n886), .ZN(n861) );
  NAND2_X1 U966 ( .A1(G112), .A2(n881), .ZN(n860) );
  NAND2_X1 U967 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n862), .B(KEYINPUT115), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G136), .A2(n887), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n882), .A2(G124), .ZN(n865) );
  XOR2_X1 U972 ( .A(KEYINPUT44), .B(n865), .Z(n866) );
  NOR2_X1 U973 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U974 ( .A(G160), .B(G162), .Z(n868) );
  XNOR2_X1 U975 ( .A(n941), .B(n868), .ZN(n873) );
  XNOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U977 ( .A(n869), .B(G164), .ZN(n870) );
  XNOR2_X1 U978 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U979 ( .A(n873), .B(n872), .ZN(n897) );
  NAND2_X1 U980 ( .A1(G118), .A2(n881), .ZN(n875) );
  NAND2_X1 U981 ( .A1(G130), .A2(n882), .ZN(n874) );
  NAND2_X1 U982 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G106), .A2(n886), .ZN(n877) );
  NAND2_X1 U984 ( .A1(G142), .A2(n887), .ZN(n876) );
  NAND2_X1 U985 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U986 ( .A(n878), .B(KEYINPUT45), .Z(n879) );
  NOR2_X1 U987 ( .A1(n880), .A2(n879), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U989 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U990 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U991 ( .A(KEYINPUT47), .B(n885), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G103), .A2(n886), .ZN(n889) );
  NAND2_X1 U993 ( .A1(G139), .A2(n887), .ZN(n888) );
  NAND2_X1 U994 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U995 ( .A(KEYINPUT116), .B(n890), .Z(n891) );
  NAND2_X1 U996 ( .A1(n892), .A2(n891), .ZN(n956) );
  XNOR2_X1 U997 ( .A(n893), .B(n956), .ZN(n894) );
  XNOR2_X1 U998 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U999 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U1000 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(n978), .B(KEYINPUT117), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(G171), .B(n977), .ZN(n901) );
  XNOR2_X1 U1004 ( .A(n902), .B(n901), .ZN(n905) );
  XOR2_X1 U1005 ( .A(G286), .B(n903), .Z(n904) );
  XNOR2_X1 U1006 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n907), .B(KEYINPUT49), .ZN(n911) );
  INV_X1 U1010 ( .A(G319), .ZN(n908) );
  NOR2_X1 U1011 ( .A1(n908), .A2(G401), .ZN(n909) );
  XOR2_X1 U1012 ( .A(KEYINPUT118), .B(n909), .Z(n910) );
  NOR2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1017 ( .A(G1966), .B(G21), .Z(n916) );
  XNOR2_X1 U1018 ( .A(n914), .B(G5), .ZN(n915) );
  NAND2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(G1976), .B(G23), .ZN(n918) );
  XNOR2_X1 U1021 ( .A(G1971), .B(G22), .ZN(n917) );
  NOR2_X1 U1022 ( .A1(n918), .A2(n917), .ZN(n920) );
  XOR2_X1 U1023 ( .A(G1986), .B(G24), .Z(n919) );
  NAND2_X1 U1024 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1025 ( .A(KEYINPUT58), .B(n921), .ZN(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n935) );
  XOR2_X1 U1027 ( .A(G4), .B(KEYINPUT126), .Z(n925) );
  XNOR2_X1 U1028 ( .A(G1348), .B(KEYINPUT59), .ZN(n924) );
  XNOR2_X1 U1029 ( .A(n925), .B(n924), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(n926), .B(G20), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(G1981), .B(G6), .ZN(n928) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n927) );
  NOR2_X1 U1033 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1036 ( .A(n933), .B(KEYINPUT60), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n936) );
  XNOR2_X1 U1039 ( .A(n937), .B(n936), .ZN(n939) );
  INV_X1 U1040 ( .A(G16), .ZN(n938) );
  NAND2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n940), .A2(G11), .ZN(n995) );
  XNOR2_X1 U1043 ( .A(G160), .B(G2084), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1046 ( .A(KEYINPUT120), .B(n945), .Z(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(n950), .B(KEYINPUT121), .ZN(n955) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n953), .Z(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G2072), .B(KEYINPUT122), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(n957), .B(n956), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G2078), .B(G164), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(KEYINPUT123), .B(n958), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1059 ( .A(KEYINPUT50), .B(n961), .Z(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(n966), .B(KEYINPUT52), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n967), .A2(G29), .ZN(n993) );
  XNOR2_X1 U1064 ( .A(KEYINPUT56), .B(G16), .ZN(n991) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n970), .B(G1956), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(G171), .B(G1961), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n977), .B(G1348), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n989) );
  XOR2_X1 U1077 ( .A(G1966), .B(G168), .Z(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n987), .Z(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n1017) );
  XOR2_X1 U1084 ( .A(KEYINPUT124), .B(G34), .Z(n997) );
  XNOR2_X1 U1085 ( .A(G2084), .B(KEYINPUT54), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n997), .B(n996), .ZN(n1012) );
  XNOR2_X1 U1087 ( .A(G2090), .B(G35), .ZN(n1010) );
  XOR2_X1 U1088 ( .A(G1991), .B(G25), .Z(n998) );
  NAND2_X1 U1089 ( .A1(n998), .A2(G28), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G1996), .B(G32), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G33), .B(G2072), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G2067), .B(G26), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G27), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT53), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT125), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(G29), .A2(n1014), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(KEYINPUT55), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

