//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  NOR2_X1   g006(.A1(G237), .A2(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G143), .A3(G214), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n192), .B1(new_n191), .B2(new_n194), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT17), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n197), .B1(KEYINPUT17), .B2(new_n196), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT71), .A3(G140), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT16), .B(new_n200), .C1(new_n204), .C2(KEYINPUT71), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT16), .B1(new_n201), .B2(G125), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n205), .B2(new_n208), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n198), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G125), .B(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n199), .A2(KEYINPUT71), .A3(G140), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT71), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n215), .B1(new_n219), .B2(new_n206), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT18), .A2(G131), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n191), .A2(new_n194), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n191), .A2(new_n194), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT18), .A3(G131), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n213), .A2(new_n229), .A3(new_n225), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G475), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT19), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n218), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n214), .A2(KEYINPUT19), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n206), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n196), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(KEYINPUT85), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n205), .A2(new_n208), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT85), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n195), .B2(new_n196), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n241), .A2(new_n244), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n249), .A2(new_n225), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n237), .B1(new_n250), .B2(new_n229), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n225), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT86), .A3(new_n230), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n232), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n255));
  NOR2_X1   g069(.A1(G475), .A2(G902), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n254), .B2(new_n256), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n236), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT9), .B(G234), .ZN(new_n260));
  INV_X1    g074(.A(G217), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n260), .A2(new_n261), .A3(G953), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT66), .B(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G143), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n190), .A2(G128), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT88), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n267), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G134), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n268), .ZN(new_n275));
  INV_X1    g089(.A(G116), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(G122), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(G122), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n277), .A2(new_n278), .A3(G107), .ZN(new_n279));
  INV_X1    g093(.A(G107), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT89), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT14), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n276), .A2(G122), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n278), .B2(KEYINPUT14), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n280), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n285), .A2(KEYINPUT89), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n279), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(new_n275), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT13), .B1(new_n190), .B2(G128), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(KEYINPUT87), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n190), .A2(KEYINPUT13), .A3(G128), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n265), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G134), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n277), .A2(new_n278), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n280), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(new_n268), .C1(new_n296), .C2(new_n279), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT90), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n289), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n289), .B2(new_n297), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n263), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n289), .A2(new_n297), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT90), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n289), .A2(new_n297), .A3(new_n298), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n262), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n305), .A3(new_n234), .ZN(new_n306));
  INV_X1    g120(.A(G478), .ZN(new_n307));
  NOR2_X1   g121(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n306), .B(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT92), .B(G952), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(G234), .A2(G237), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT21), .B(G898), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(G902), .A3(G953), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n259), .A2(new_n312), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n206), .A2(G143), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n190), .A2(G146), .ZN(new_n324));
  AND2_X1   g138(.A1(KEYINPUT0), .A2(G128), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT64), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT64), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n324), .ZN(new_n330));
  NOR2_X1   g144(.A1(KEYINPUT0), .A2(G128), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n327), .A2(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G125), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n330), .B1(new_n336), .B2(new_n264), .ZN(new_n337));
  INV_X1    g151(.A(G128), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT1), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n323), .A3(new_n324), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n334), .B1(G125), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n188), .A2(G224), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n345));
  AND4_X1   g159(.A1(KEYINPUT7), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n347), .B(KEYINPUT8), .Z(new_n348));
  OR2_X1    g162(.A1(KEYINPUT67), .A2(G119), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT67), .A2(G119), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(G116), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G119), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(G116), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(KEYINPUT5), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n355), .B(G113), .C1(KEYINPUT5), .C2(new_n351), .ZN(new_n356));
  INV_X1    g170(.A(G113), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT2), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G113), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n351), .A2(new_n354), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n280), .A3(G104), .ZN(new_n366));
  INV_X1    g180(.A(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n228), .A2(G107), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n364), .A2(new_n366), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n228), .A2(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n280), .A2(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(G101), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n369), .A2(new_n372), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n356), .A2(new_n362), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n348), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n343), .A2(new_n345), .B1(KEYINPUT7), .B2(new_n344), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n346), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G101), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n351), .A2(new_n354), .A3(new_n361), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n361), .B1(new_n351), .B2(new_n354), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n380), .A2(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT82), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n361), .ZN(new_n390));
  INV_X1    g204(.A(new_n350), .ZN(new_n391));
  NOR2_X1   g205(.A1(KEYINPUT67), .A2(G119), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(new_n276), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n390), .B1(new_n393), .B2(new_n353), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n362), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n380), .A2(G101), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n395), .A2(new_n397), .A3(new_n398), .A4(new_n382), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n389), .A2(new_n347), .A3(new_n399), .A4(new_n376), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n399), .A2(new_n376), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n403), .A2(KEYINPUT83), .A3(new_n347), .A4(new_n389), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(G902), .B1(new_n379), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n347), .B1(new_n403), .B2(new_n389), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n407), .A2(KEYINPUT6), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n400), .A2(new_n401), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n400), .A2(new_n401), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT6), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n407), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n343), .B(new_n344), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n406), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G210), .B1(G237), .B2(G902), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n407), .B1(new_n405), .B2(KEYINPUT6), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n414), .B1(new_n420), .B2(new_n408), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n406), .A3(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT81), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n322), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT11), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n266), .B2(G137), .ZN(new_n429));
  INV_X1    g243(.A(G137), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT11), .A3(G134), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n266), .A2(G137), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n429), .A2(new_n431), .A3(new_n192), .A4(new_n432), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(KEYINPUT65), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n437), .A3(G131), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n333), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n440));
  INV_X1    g254(.A(new_n432), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n266), .A2(G137), .ZN(new_n442));
  OAI21_X1  g256(.A(G131), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n341), .A2(new_n435), .A3(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n440), .B1(new_n439), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n395), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n395), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(new_n448), .A3(new_n444), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n193), .A2(G210), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT27), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT26), .B(G101), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n447), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n447), .A2(KEYINPUT68), .A3(new_n449), .A4(new_n453), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(KEYINPUT31), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n453), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT28), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n439), .A2(new_n444), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n395), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n462), .B2(new_n449), .ZN(new_n463));
  INV_X1    g277(.A(new_n449), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT28), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT31), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n447), .A2(new_n467), .A3(new_n449), .A4(new_n453), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n458), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G472), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n234), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT32), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n458), .B2(new_n469), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT32), .A3(new_n471), .ZN(new_n476));
  OR3_X1    g290(.A1(new_n463), .A2(new_n465), .A3(new_n459), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n478));
  INV_X1    g292(.A(new_n447), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n459), .B1(new_n479), .B2(new_n464), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n234), .B1(new_n477), .B2(new_n478), .ZN(new_n482));
  OAI21_X1  g296(.A(G472), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n474), .A2(new_n476), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT74), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n349), .A2(G128), .A3(new_n350), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT66), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G128), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n489), .A3(G119), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT24), .B(G110), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n491), .B2(new_n493), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G110), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n264), .A2(KEYINPUT23), .A3(G119), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n486), .A2(KEYINPUT70), .A3(KEYINPUT23), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n338), .B1(new_n391), .B2(new_n392), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT70), .B1(new_n486), .B2(KEYINPUT23), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n497), .B(new_n498), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n207), .B1(new_n218), .B2(KEYINPUT16), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n215), .B1(new_n505), .B2(new_n206), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n491), .A2(new_n493), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n246), .B2(new_n209), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G110), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n504), .A2(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n485), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n504), .A2(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n509), .A2(new_n511), .ZN(new_n518));
  AND4_X1   g332(.A1(new_n485), .A2(new_n517), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n521));
  OAI22_X1  g335(.A1(new_n210), .A2(new_n211), .B1(new_n491), .B2(new_n493), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n486), .A2(KEYINPUT23), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n499), .A3(new_n500), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n497), .B1(new_n526), .B2(new_n498), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n506), .B1(new_n503), .B2(new_n496), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n515), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT73), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n520), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(G217), .A2(G902), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n261), .B2(G234), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n536), .B(KEYINPUT69), .Z(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n517), .A2(new_n518), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT74), .B1(new_n541), .B2(new_n531), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n512), .A2(new_n485), .A3(new_n515), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n533), .A2(new_n542), .A3(new_n234), .A4(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n520), .A2(KEYINPUT25), .A3(new_n234), .A4(new_n533), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n540), .B1(new_n548), .B2(new_n537), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n342), .A2(new_n373), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n335), .A2(G128), .B1(new_n323), .B2(new_n324), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n339), .A2(new_n323), .A3(new_n324), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT77), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n553), .A2(new_n373), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n330), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n338), .B1(new_n323), .B2(KEYINPUT1), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n340), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT77), .B1(new_n375), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n550), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n436), .A2(new_n438), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT78), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n436), .A2(new_n564), .A3(new_n438), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n560), .A2(new_n562), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n554), .B1(new_n553), .B2(new_n373), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n558), .A2(KEYINPUT77), .A3(new_n369), .A4(new_n372), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n567), .A2(new_n568), .B1(new_n342), .B2(new_n373), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n563), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n569), .A2(new_n570), .A3(new_n561), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT80), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G140), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n188), .A2(G227), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n397), .A2(new_n333), .A3(new_n382), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n337), .B2(new_n340), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n578), .A2(KEYINPUT76), .B1(new_n375), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n579), .B1(new_n555), .B2(new_n559), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n397), .A2(new_n333), .A3(new_n583), .A4(new_n382), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n581), .A2(new_n582), .A3(new_n561), .A4(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n572), .A2(new_n573), .A3(new_n577), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n562), .A2(KEYINPUT79), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n327), .A2(new_n329), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n330), .A2(new_n332), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n382), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT76), .B1(new_n591), .B2(new_n388), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n580), .A2(new_n375), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n584), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT10), .B1(new_n567), .B2(new_n568), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n581), .A2(new_n582), .A3(new_n587), .A4(new_n584), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n576), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n565), .A2(new_n563), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n560), .A2(new_n600), .A3(new_n562), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n570), .B1(new_n569), .B2(new_n561), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n585), .A2(new_n577), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n586), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G469), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n234), .ZN(new_n607));
  NAND2_X1  g421(.A1(G469), .A2(G902), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n585), .A2(new_n602), .A3(new_n601), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n576), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n596), .A2(new_n577), .A3(new_n597), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(G469), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G221), .B1(new_n260), .B2(G902), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT75), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n427), .A2(new_n484), .A3(new_n549), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  XNOR2_X1  g433(.A(new_n475), .B(new_n471), .ZN(new_n620));
  INV_X1    g434(.A(new_n549), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n617), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n307), .A2(G902), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n302), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n305), .A3(new_n301), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n301), .B2(new_n305), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n306), .A2(new_n307), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n259), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n321), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT93), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n419), .A2(new_n637), .A3(new_n422), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n421), .A2(KEYINPUT93), .A3(new_n406), .A4(new_n417), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n639), .A2(new_n426), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n635), .A2(new_n636), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n623), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  INV_X1    g459(.A(new_n311), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n306), .B(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n259), .A2(new_n647), .A3(new_n321), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n638), .A2(new_n648), .A3(new_n640), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT95), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n638), .A2(new_n648), .A3(new_n640), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n623), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NAND2_X1  g470(.A1(new_n530), .A2(new_n532), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n531), .A2(KEYINPUT36), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n548), .A2(new_n537), .B1(new_n538), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n620), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n427), .A2(new_n617), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT96), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n548), .A2(new_n537), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n661), .A2(new_n538), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n484), .A2(new_n617), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n316), .B1(G900), .B2(new_n319), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n259), .A2(new_n647), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n638), .A2(new_n674), .A3(new_n640), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT97), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n638), .A2(new_n674), .A3(new_n640), .A4(KEYINPUT97), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n671), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT98), .B(G128), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G30));
  XNOR2_X1  g495(.A(new_n423), .B(KEYINPUT38), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n456), .A2(new_n457), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n453), .B1(new_n462), .B2(new_n449), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n234), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n474), .A3(new_n476), .ZN(new_n687));
  INV_X1    g501(.A(new_n258), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n688), .A2(new_n689), .B1(G475), .B2(new_n235), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n647), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n426), .A3(new_n662), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n682), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n672), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n617), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n693), .B1(KEYINPUT40), .B2(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  AND2_X1   g513(.A1(new_n638), .A2(new_n640), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n633), .A2(new_n259), .A3(new_n672), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n671), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  AOI21_X1  g518(.A(new_n606), .B1(new_n605), .B2(new_n234), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT99), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n607), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n707), .B(new_n606), .C1(new_n605), .C2(new_n234), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n615), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n484), .A3(new_n549), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n641), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT100), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n713), .B(new_n715), .ZN(G15));
  AOI21_X1  g530(.A(new_n712), .B1(new_n650), .B2(new_n652), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n276), .ZN(G18));
  NAND3_X1  g532(.A1(new_n484), .A2(new_n322), .A3(new_n670), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n638), .A2(new_n640), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n607), .A2(new_n707), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n705), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n616), .B1(new_n722), .B2(new_n709), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n352), .ZN(G21));
  AOI21_X1  g539(.A(new_n471), .B1(new_n470), .B2(new_n234), .ZN(new_n726));
  AOI211_X1 g540(.A(G472), .B(G902), .C1(new_n458), .C2(new_n469), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n728), .A2(new_n549), .A3(new_n636), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n700), .A3(new_n691), .A4(new_n711), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR3_X1   g545(.A1(new_n723), .A2(new_n720), .A3(new_n701), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n662), .A2(new_n726), .A3(new_n727), .A4(KEYINPUT101), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT101), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n728), .B2(new_n670), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  NAND2_X1  g552(.A1(new_n484), .A2(new_n549), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n702), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n419), .A2(new_n426), .A3(new_n422), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n610), .A2(KEYINPUT102), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT102), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n609), .A2(new_n746), .A3(new_n576), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(G469), .A3(new_n611), .A4(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n607), .A2(new_n608), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n616), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n419), .A2(KEYINPUT103), .A3(new_n426), .A4(new_n422), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n744), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n744), .A2(new_n754), .A3(new_n750), .A4(new_n751), .ZN(new_n755));
  AOI211_X1 g569(.A(new_n739), .B(new_n741), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n755), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n474), .A2(new_n758), .A3(new_n476), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n472), .A2(KEYINPUT105), .A3(new_n473), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n483), .A3(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n757), .A2(new_n765), .A3(new_n549), .A4(new_n702), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n756), .B1(new_n766), .B2(KEYINPUT42), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND4_X1  g582(.A1(new_n757), .A2(new_n484), .A3(new_n549), .A4(new_n674), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n301), .A2(new_n305), .ZN(new_n772));
  INV_X1    g586(.A(new_n627), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n628), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n775), .A2(new_n624), .B1(new_n307), .B2(new_n306), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n771), .B1(new_n776), .B2(new_n259), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n690), .A2(new_n633), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n771), .A3(KEYINPUT43), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n728), .A2(new_n662), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(KEYINPUT44), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n744), .A2(new_n751), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n782), .A2(new_n783), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT44), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n612), .B1(new_n792), .B2(new_n606), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n745), .A2(KEYINPUT45), .A3(new_n611), .A4(new_n747), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT46), .B1(new_n797), .B2(new_n608), .ZN(new_n798));
  INV_X1    g612(.A(new_n607), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n608), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n615), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(new_n694), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n784), .A2(KEYINPUT109), .A3(new_n786), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n789), .A2(new_n791), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n800), .A2(new_n801), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n616), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n785), .A2(new_n484), .A3(new_n549), .A4(new_n701), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n807), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(new_n807), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  INV_X1    g634(.A(new_n622), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n779), .A2(new_n781), .A3(new_n317), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT113), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n779), .A2(new_n781), .A3(new_n824), .A4(new_n317), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n786), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n802), .B(new_n810), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n615), .B1(new_n722), .B2(new_n709), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n711), .A2(new_n744), .A3(new_n751), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n823), .B2(new_n825), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n831), .A2(new_n687), .A3(new_n621), .A4(new_n316), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n633), .A2(new_n259), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n832), .A2(new_n736), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n682), .A2(new_n426), .A3(new_n723), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n826), .A2(KEYINPUT50), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT50), .B1(new_n826), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n820), .B1(new_n830), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n811), .A2(new_n812), .A3(new_n829), .ZN(new_n842));
  INV_X1    g656(.A(new_n827), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n826), .A2(new_n836), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n837), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n844), .A2(new_n848), .A3(KEYINPUT51), .A4(new_n835), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n826), .A2(new_n700), .A3(new_n711), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n833), .A2(new_n635), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n850), .A2(new_n314), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n832), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n765), .A2(new_n549), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n853), .A2(KEYINPUT48), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT48), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n841), .A2(new_n849), .A3(new_n852), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n844), .A2(new_n848), .A3(new_n835), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n861), .A2(new_n820), .B1(new_n856), .B2(new_n855), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT114), .A3(new_n849), .A4(new_n852), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT101), .B1(new_n620), .B2(new_n662), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n728), .A2(new_n670), .A3(new_n734), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n635), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n753), .B2(new_n755), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n259), .A2(new_n312), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n786), .A2(new_n671), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n672), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n717), .A2(new_n724), .A3(new_n713), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n312), .B(new_n236), .C1(new_n258), .C2(new_n257), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n321), .B1(new_n634), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n425), .B1(new_n419), .B2(new_n422), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n622), .A2(new_n873), .A3(new_n617), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n730), .A2(new_n618), .A3(new_n664), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n870), .A2(new_n871), .A3(new_n769), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n766), .A2(KEYINPUT42), .ZN(new_n879));
  INV_X1    g693(.A(new_n756), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n616), .A2(new_n662), .A3(new_n672), .A4(new_n749), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n700), .A3(new_n687), .A4(new_n691), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n737), .A2(new_n679), .A3(new_n703), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT112), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT52), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT111), .B1(new_n885), .B2(KEYINPUT112), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n885), .B2(KEYINPUT111), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n882), .B2(new_n892), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n876), .A2(new_n717), .A3(new_n713), .A4(new_n724), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n767), .A2(new_n769), .A3(new_n894), .A4(new_n870), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n885), .B(KEYINPUT52), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n882), .A2(new_n892), .A3(KEYINPUT53), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n860), .A2(new_n863), .A3(new_n899), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(G952), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n188), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n722), .A2(new_n709), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT49), .ZN(new_n909));
  OR4_X1    g723(.A1(new_n621), .A2(new_n780), .A3(new_n615), .A4(new_n425), .ZN(new_n910));
  OR4_X1    g724(.A1(new_n687), .A2(new_n909), .A3(new_n682), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n907), .A2(KEYINPUT115), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(G75));
  NAND2_X1  g730(.A1(new_n905), .A2(G953), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT117), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n234), .B1(new_n900), .B2(new_n901), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n413), .B(new_n414), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(G51));
  INV_X1    g742(.A(new_n918), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n608), .B(KEYINPUT57), .Z(new_n930));
  AND3_X1   g744(.A1(new_n900), .A2(new_n902), .A3(new_n901), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n605), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n919), .A2(new_n795), .A3(new_n796), .A4(new_n794), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(G54));
  NAND3_X1  g750(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n254), .Z(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n929), .ZN(G60));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n775), .B(KEYINPUT118), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n931), .B2(new_n932), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT119), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT119), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n945), .C1(new_n931), .C2(new_n932), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n944), .B1(new_n899), .B2(new_n903), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n918), .B1(new_n951), .B2(new_n941), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n940), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n944), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n882), .A2(new_n892), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n896), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n902), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n954), .B1(new_n958), .B2(new_n931), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n929), .B1(new_n959), .B2(new_n942), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(KEYINPUT120), .A3(new_n947), .A4(new_n949), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n953), .A2(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(new_n900), .A2(new_n901), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n535), .B(KEYINPUT121), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n929), .B1(new_n966), .B2(new_n534), .ZN(new_n967));
  INV_X1    g781(.A(new_n661), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n966), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  INV_X1    g785(.A(new_n894), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n188), .ZN(new_n973));
  INV_X1    g787(.A(G224), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n318), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(KEYINPUT122), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(KEYINPUT122), .B2(new_n973), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n413), .B1(G898), .B2(new_n188), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT123), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n977), .B(new_n979), .ZN(G69));
  AND2_X1   g794(.A1(new_n679), .A2(new_n703), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n737), .ZN(new_n982));
  INV_X1    g796(.A(new_n854), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n803), .A2(new_n700), .A3(new_n691), .A4(new_n983), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n769), .A2(new_n805), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n818), .A2(new_n985), .A3(new_n188), .A4(new_n767), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n445), .A2(new_n446), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n239), .A2(new_n240), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n986), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n634), .A2(new_n872), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n785), .A2(new_n739), .A3(new_n695), .A4(new_n997), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT124), .Z(new_n999));
  NAND2_X1  g813(.A1(new_n805), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n817), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n815), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n698), .A2(new_n737), .A3(new_n981), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT62), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n996), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1000), .B1(new_n816), .B2(new_n817), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1004), .B(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1007), .A2(KEYINPUT125), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(G953), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n993), .B(new_n995), .C1(new_n1011), .C2(new_n989), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT126), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1003), .A2(new_n996), .A3(new_n1005), .ZN(new_n1016));
  AOI21_X1  g830(.A(KEYINPUT125), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n188), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n990), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1013), .B1(new_n986), .B2(new_n991), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1015), .B(new_n1020), .C1(new_n1011), .C2(new_n989), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1014), .B1(new_n1021), .B2(new_n1023), .ZN(G72));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT63), .Z(new_n1026));
  NAND3_X1  g840(.A1(new_n818), .A2(new_n985), .A3(new_n767), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1026), .B1(new_n1027), .B2(new_n972), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1028), .A2(new_n449), .A3(new_n447), .A4(new_n459), .ZN(new_n1029));
  INV_X1    g843(.A(new_n480), .ZN(new_n1030));
  OAI221_X1 g844(.A(new_n1026), .B1(new_n683), .B2(new_n1030), .C1(new_n893), .C2(new_n898), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1029), .A2(new_n918), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1006), .A2(new_n894), .A3(new_n1010), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1026), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n459), .B1(new_n447), .B2(new_n449), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(G57));
endmodule


