//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n207), .C1(new_n203), .C2(new_n204), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(G190gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n210), .B1(new_n212), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(new_n215), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n216), .A2(new_n211), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n224), .B2(new_n208), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n214), .B2(KEYINPUT27), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT27), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT27), .B1(new_n217), .B2(new_n218), .ZN(new_n233));
  NOR2_X1   g032(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT28), .B1(new_n238), .B2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT69), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n245), .A2(KEYINPUT26), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n245), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n246), .A2(new_n247), .B1(G183gat), .B2(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n227), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n235), .A2(new_n242), .A3(new_n239), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n242), .B1(new_n235), .B2(new_n239), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n227), .B(new_n248), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n226), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(G113gat), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(KEYINPUT71), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(KEYINPUT71), .B2(new_n257), .ZN(new_n259));
  XOR2_X1   g058(.A(G127gat), .B(G134gat), .Z(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G120gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n265), .B2(new_n256), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n202), .B1(new_n254), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(new_n252), .B1(new_n225), .B2(new_n221), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n259), .A2(new_n261), .B1(new_n266), .B2(new_n260), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(KEYINPUT72), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n268), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n269), .A2(new_n270), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT34), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT32), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n269), .A2(new_n276), .A3(new_n275), .ZN(new_n280));
  INV_X1    g079(.A(new_n270), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT33), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  XNOR2_X1  g082(.A(G15gat), .B(G43gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n282), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  AOI221_X4 g087(.A(new_n279), .B1(KEYINPUT33), .B2(new_n286), .C1(new_n280), .C2(new_n281), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n278), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT73), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n283), .A2(new_n287), .ZN(new_n292));
  INV_X1    g091(.A(new_n282), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n278), .ZN(new_n295));
  INV_X1    g094(.A(new_n289), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n291), .B1(new_n299), .B2(KEYINPUT73), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT74), .B(G197gat), .Z(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G204gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT74), .B(G197gat), .ZN(new_n307));
  INV_X1    g106(.A(G204gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310));
  INV_X1    g109(.A(G211gat), .ZN(new_n311));
  INV_X1    g110(.A(G218gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n306), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n271), .A2(new_n317), .A3(new_n226), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(KEYINPUT29), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n316), .B(new_n318), .C1(new_n273), .C2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n317), .B(new_n226), .C1(new_n249), .C2(new_n253), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n271), .A2(new_n226), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n319), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n328));
  INV_X1    g127(.A(new_n323), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n254), .A2(new_n319), .B1(new_n317), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(KEYINPUT75), .A3(new_n316), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n327), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n327), .B2(new_n331), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n304), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n304), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n327), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n342), .B(KEYINPUT79), .Z(new_n343));
  XOR2_X1   g142(.A(G141gat), .B(G148gat), .Z(new_n344));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT2), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n345), .B(KEYINPUT78), .Z(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  INV_X1    g149(.A(new_n345), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n344), .B(new_n346), .C1(new_n351), .C2(new_n342), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n353), .A2(new_n268), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n352), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT4), .B1(new_n268), .B2(new_n355), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n274), .A2(new_n349), .A3(new_n358), .A4(new_n352), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n354), .A2(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT5), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n360), .A2(KEYINPUT82), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n357), .A2(new_n359), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n268), .A3(new_n353), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n361), .A4(new_n362), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n360), .A2(new_n362), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n268), .B(new_n355), .ZN(new_n371));
  INV_X1    g170(.A(new_n362), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n361), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT81), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT80), .ZN(new_n378));
  XOR2_X1   g177(.A(G57gat), .B(G85gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n378), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n363), .A2(new_n368), .B1(new_n370), .B2(new_n373), .ZN(new_n384));
  INV_X1    g183(.A(new_n381), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT89), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n382), .A2(new_n386), .A3(new_n389), .A4(new_n383), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n384), .A2(new_n385), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT6), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT86), .B1(new_n316), .B2(KEYINPUT29), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n350), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n316), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n355), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n353), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n316), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n316), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n399), .A3(new_n355), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n316), .A2(new_n400), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n356), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n406), .A2(KEYINPUT85), .A3(new_n398), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT85), .B1(new_n406), .B2(new_n398), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT31), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT31), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n402), .B(new_n411), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(G22gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G50gat), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n410), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n410), .B2(new_n412), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(KEYINPUT35), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n301), .A2(new_n341), .A3(new_n393), .A4(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n334), .A2(new_n422), .A3(new_n338), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n387), .A2(new_n392), .B1(new_n337), .B2(new_n336), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n334), .B2(new_n338), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT83), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n333), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n327), .A2(new_n328), .A3(new_n331), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n335), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n336), .A2(new_n337), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT77), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n423), .A4(new_n424), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n298), .A2(new_n419), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n427), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT93), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT35), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n436), .B2(KEYINPUT35), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n421), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT37), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n327), .A2(new_n441), .A3(new_n331), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n330), .A2(new_n403), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n322), .A2(new_n324), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n316), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(KEYINPUT37), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n450));
  NOR2_X1   g249(.A1(new_n335), .A2(new_n450), .ZN(new_n451));
  AND4_X1   g250(.A1(new_n442), .A2(new_n448), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n393), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n327), .ZN(new_n454));
  INV_X1    g253(.A(new_n331), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n456), .B2(new_n335), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n304), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n428), .A2(new_n429), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(KEYINPUT37), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n453), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n360), .A2(new_n362), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n463));
  OR3_X1    g262(.A1(new_n371), .A2(new_n463), .A3(new_n372), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n371), .B2(new_n372), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(KEYINPUT39), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n466), .B2(KEYINPUT88), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(KEYINPUT88), .B2(new_n466), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n381), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n468), .A2(KEYINPUT40), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT40), .B1(new_n468), .B2(new_n470), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n471), .A2(new_n472), .A3(new_n391), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n419), .B1(new_n473), .B2(new_n340), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n461), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT92), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  INV_X1    g276(.A(new_n291), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT73), .B1(new_n290), .B2(new_n297), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n298), .B2(new_n477), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n427), .A2(new_n434), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n419), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n461), .A2(new_n484), .A3(new_n474), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n476), .A2(new_n481), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n440), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT106), .ZN(new_n488));
  INV_X1    g287(.A(G71gat), .ZN(new_n489));
  INV_X1    g288(.A(G78gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(G71gat), .A2(G78gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(KEYINPUT98), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(KEYINPUT98), .B2(new_n492), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n491), .A2(KEYINPUT9), .ZN(new_n495));
  XOR2_X1   g294(.A(G57gat), .B(G64gat), .Z(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n495), .B(new_n496), .C1(new_n491), .C2(new_n492), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(KEYINPUT99), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n498), .A2(KEYINPUT99), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G85gat), .ZN(new_n502));
  INV_X1    g301(.A(G92gat), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT101), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT101), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(G85gat), .A3(G92gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(KEYINPUT7), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508));
  OAI211_X1 g307(.A(KEYINPUT101), .B(new_n508), .C1(new_n502), .C2(new_n503), .ZN(new_n509));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510));
  AOI22_X1  g309(.A1(KEYINPUT8), .A2(new_n510), .B1(new_n502), .B2(new_n503), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G99gat), .B(G106gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n501), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n516), .B(KEYINPUT104), .Z(new_n517));
  AND2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT100), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n501), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT100), .B1(new_n499), .B2(new_n500), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT10), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n514), .B(KEYINPUT102), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n522), .A2(new_n524), .B1(new_n515), .B2(KEYINPUT10), .ZN(new_n525));
  INV_X1    g324(.A(new_n517), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n518), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT105), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n488), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AOI211_X1 g334(.A(KEYINPUT105), .B(KEYINPUT106), .C1(new_n527), .C2(new_n531), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n527), .A2(new_n531), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI22_X1  g338(.A1(new_n534), .A2(new_n536), .B1(new_n527), .B2(new_n531), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n501), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G15gat), .B(G22gat), .Z(new_n545));
  INV_X1    g344(.A(G1gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n548));
  AOI21_X1  g347(.A(G8gat), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n546), .A2(KEYINPUT16), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n547), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n549), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n520), .A2(new_n521), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n555), .B2(new_n543), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n556), .B2(new_n544), .ZN(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n214), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(new_n311), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n557), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G127gat), .B(G155gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n564), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OR3_X1    g367(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n569), .A2(new_n570), .B1(G29gat), .B2(G36gat), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n572));
  XNOR2_X1  g371(.A(G43gat), .B(G50gat), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT17), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n552), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n553), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G169gat), .B(G197gat), .Z(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT94), .B(KEYINPUT11), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT12), .Z(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n584), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT96), .B1(new_n581), .B2(new_n553), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n582), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n580), .B(KEYINPUT13), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n585), .A2(new_n591), .A3(new_n592), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT97), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n592), .A2(new_n597), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n591), .A4(new_n585), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n585), .ZN(new_n604));
  INV_X1    g403(.A(new_n591), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n578), .A2(new_n524), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(KEYINPUT103), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n609), .B(new_n613), .C1(new_n577), .C2(new_n524), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(KEYINPUT103), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n616), .B(new_n619), .ZN(new_n620));
  NOR4_X1   g419(.A1(new_n542), .A2(new_n568), .A3(new_n608), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n487), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n387), .A2(new_n392), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT107), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT108), .B(G1gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(G1324gat));
  NOR2_X1   g426(.A1(new_n622), .A2(new_n341), .ZN(new_n628));
  INV_X1    g427(.A(G8gat), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT42), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT16), .B(G8gat), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  MUX2_X1   g431(.A(KEYINPUT42), .B(new_n630), .S(new_n632), .Z(G1325gat));
  INV_X1    g432(.A(new_n622), .ZN(new_n634));
  AOI21_X1  g433(.A(G15gat), .B1(new_n634), .B2(new_n301), .ZN(new_n635));
  INV_X1    g434(.A(new_n481), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(G15gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT109), .Z(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n634), .B2(new_n638), .ZN(G1326gat));
  INV_X1    g438(.A(new_n419), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n622), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT43), .B(G22gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n620), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n440), .B2(new_n486), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n542), .A2(new_n608), .A3(new_n567), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n647), .A2(G29gat), .A3(new_n624), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n487), .B2(new_n620), .ZN(new_n652));
  AOI211_X1 g451(.A(KEYINPUT44), .B(new_n644), .C1(new_n440), .C2(new_n486), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n646), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G29gat), .B1(new_n654), .B2(new_n624), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(G1328gat));
  OR2_X1    g455(.A1(new_n341), .A2(G36gat), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT46), .B1(new_n647), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT111), .ZN(new_n659));
  OAI21_X1  g458(.A(G36gat), .B1(new_n654), .B2(new_n341), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n647), .A2(new_n657), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n659), .B(new_n660), .C1(KEYINPUT46), .C2(new_n661), .ZN(G1329gat));
  OAI21_X1  g461(.A(G43gat), .B1(new_n654), .B2(new_n481), .ZN(new_n663));
  OR3_X1    g462(.A1(new_n647), .A2(G43gat), .A3(new_n300), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1330gat));
  NOR3_X1   g466(.A1(new_n647), .A2(G50gat), .A3(new_n640), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n419), .B(new_n646), .C1(new_n652), .C2(new_n653), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(G50gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g470(.A1(new_n608), .A2(new_n567), .A3(new_n644), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n541), .B(new_n672), .C1(new_n440), .C2(new_n486), .ZN(new_n673));
  INV_X1    g472(.A(new_n624), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n340), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT49), .B(G64gat), .Z(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n677), .B2(new_n679), .ZN(G1333gat));
  AOI21_X1  g479(.A(new_n489), .B1(new_n673), .B2(new_n636), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n300), .A2(G71gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n673), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g483(.A1(new_n673), .A2(new_n419), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g485(.A1(new_n567), .A2(new_n607), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n541), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n652), .B2(new_n653), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(KEYINPUT112), .A3(new_n674), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G85gat), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT112), .B1(new_n691), .B2(new_n674), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n645), .A2(new_n687), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n541), .B1(new_n695), .B2(KEYINPUT51), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT51), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n645), .A2(new_n697), .A3(new_n687), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n674), .A2(new_n502), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n693), .A2(new_n694), .B1(new_n699), .B2(new_n700), .ZN(G1336gat));
  NAND2_X1  g500(.A1(new_n695), .A2(KEYINPUT51), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n341), .A2(G92gat), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n702), .A2(new_n542), .A3(new_n698), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT114), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT52), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n696), .A2(new_n707), .A3(new_n698), .A4(new_n703), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n340), .B(new_n689), .C1(new_n652), .C2(new_n653), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G92gat), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n705), .A2(new_n706), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT113), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n704), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(KEYINPUT52), .ZN(new_n714));
  AOI211_X1 g513(.A(KEYINPUT113), .B(new_n706), .C1(new_n710), .C2(new_n704), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(G1337gat));
  NOR2_X1   g515(.A1(new_n690), .A2(new_n481), .ZN(new_n717));
  INV_X1    g516(.A(G99gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n301), .A2(new_n718), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n699), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT115), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT115), .ZN(new_n723));
  OAI221_X1 g522(.A(new_n723), .B1(new_n699), .B2(new_n720), .C1(new_n717), .C2(new_n718), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1338gat));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n640), .A2(G106gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n696), .A2(new_n698), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT116), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G106gat), .B1(new_n690), .B2(new_n640), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n728), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n730), .B(new_n732), .ZN(G1339gat));
  NOR2_X1   g532(.A1(new_n624), .A2(new_n340), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n525), .A2(new_n526), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n531), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n525), .B2(new_n526), .ZN(new_n739));
  OAI221_X1 g538(.A(new_n517), .B1(new_n515), .B2(KEYINPUT10), .C1(new_n524), .C2(new_n522), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n739), .A2(KEYINPUT117), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT117), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI211_X1 g541(.A(KEYINPUT55), .B(new_n738), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n532), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT118), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(KEYINPUT118), .A3(new_n532), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n746), .A2(new_n607), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n579), .A2(new_n582), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n752), .A2(new_n580), .B1(new_n596), .B2(new_n594), .ZN(new_n753));
  INV_X1    g552(.A(new_n590), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n539), .A2(new_n540), .A3(new_n603), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n620), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n620), .A2(new_n603), .A3(new_n755), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n758), .A2(new_n746), .A3(new_n747), .A4(new_n750), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n568), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n672), .A2(new_n542), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n735), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n300), .A2(new_n419), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G113gat), .B1(new_n766), .B2(new_n608), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n435), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n607), .A2(new_n264), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT119), .Z(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(G1340gat));
  OAI21_X1  g570(.A(G120gat), .B1(new_n766), .B2(new_n541), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n542), .A2(new_n255), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n768), .B2(new_n773), .ZN(G1341gat));
  INV_X1    g573(.A(new_n768), .ZN(new_n775));
  AOI21_X1  g574(.A(G127gat), .B1(new_n775), .B2(new_n567), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n764), .A2(G127gat), .A3(new_n567), .A4(new_n765), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(KEYINPUT120), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(KEYINPUT120), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(G1342gat));
  OAI21_X1  g579(.A(G134gat), .B1(new_n766), .B2(new_n644), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n768), .A2(G134gat), .A3(new_n644), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n782), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT121), .B1(new_n782), .B2(KEYINPUT56), .ZN(new_n784));
  OAI221_X1 g583(.A(new_n781), .B1(KEYINPUT56), .B2(new_n782), .C1(new_n783), .C2(new_n784), .ZN(G1343gat));
  AOI21_X1  g584(.A(new_n640), .B1(new_n761), .B2(new_n763), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n481), .A2(new_n734), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(G141gat), .A3(new_n608), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n607), .A2(new_n750), .A3(new_n532), .A4(new_n743), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n756), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n644), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n567), .B1(new_n795), .B2(new_n759), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n419), .B1(new_n796), .B2(new_n762), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n787), .B1(new_n797), .B2(KEYINPUT57), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n786), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n798), .A2(new_n800), .A3(new_n607), .ZN(new_n801));
  INV_X1    g600(.A(G141gat), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n791), .B(new_n792), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n798), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n798), .B2(new_n800), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n607), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n790), .B1(new_n808), .B2(G141gat), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(G1344gat));
  OR3_X1    g610(.A1(new_n789), .A2(G148gat), .A3(new_n541), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G148gat), .ZN(new_n814));
  INV_X1    g613(.A(new_n807), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n805), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n542), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n786), .A2(KEYINPUT57), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n797), .A2(new_n799), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n542), .A3(new_n788), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n813), .B1(new_n821), .B2(G148gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n812), .B1(new_n817), .B2(new_n822), .ZN(G1345gat));
  INV_X1    g622(.A(new_n789), .ZN(new_n824));
  AOI21_X1  g623(.A(G155gat), .B1(new_n824), .B2(new_n567), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n567), .A2(G155gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n816), .B2(new_n826), .ZN(G1346gat));
  NOR3_X1   g626(.A1(new_n789), .A2(G162gat), .A3(new_n644), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT124), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n644), .B1(new_n815), .B2(new_n805), .ZN(new_n830));
  INV_X1    g629(.A(G162gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G1347gat));
  NOR2_X1   g631(.A1(new_n674), .A2(new_n341), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n761), .B2(new_n763), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n765), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G169gat), .B1(new_n837), .B2(new_n608), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n835), .A2(new_n435), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n203), .A3(new_n607), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1348gat));
  AOI21_X1  g640(.A(G176gat), .B1(new_n839), .B2(new_n542), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n541), .A2(new_n204), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n836), .B2(new_n843), .ZN(G1349gat));
  NAND2_X1  g643(.A1(new_n836), .A2(new_n567), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n568), .A2(new_n238), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n845), .A2(new_n219), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT125), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT126), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(KEYINPUT126), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n847), .B2(new_n849), .ZN(G1350gat));
  NAND3_X1  g652(.A1(new_n839), .A2(new_n215), .A3(new_n620), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n215), .B1(new_n836), .B2(new_n620), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(G1351gat));
  NOR2_X1   g658(.A1(new_n636), .A2(new_n834), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n786), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(G197gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n607), .ZN(new_n863));
  INV_X1    g662(.A(new_n860), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n818), .B2(new_n819), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n607), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n863), .B1(new_n866), .B2(new_n862), .ZN(G1352gat));
  NAND3_X1  g666(.A1(new_n861), .A2(new_n308), .A3(new_n542), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT62), .Z(new_n869));
  AOI211_X1 g668(.A(new_n541), .B(new_n864), .C1(new_n818), .C2(new_n819), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n308), .B2(new_n870), .ZN(G1353gat));
  NAND3_X1  g670(.A1(new_n861), .A2(new_n311), .A3(new_n567), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n865), .A2(new_n567), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT63), .B1(new_n873), .B2(G211gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(G1354gat));
  AND2_X1   g675(.A1(new_n865), .A2(KEYINPUT127), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n620), .B1(new_n865), .B2(KEYINPUT127), .ZN(new_n878));
  OAI21_X1  g677(.A(G218gat), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n312), .A3(new_n620), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1355gat));
endmodule


