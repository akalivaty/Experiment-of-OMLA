//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n210), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n213), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n212), .B1(new_n221), .B2(KEYINPUT0), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT0), .B2(new_n221), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT64), .Z(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n226), .B2(new_n213), .C1(new_n227), .C2(new_n219), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  INV_X1    g0029(.A(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G77), .ZN(new_n231));
  INV_X1    g0031(.A(G244), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n229), .B1(new_n202), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n216), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  AND2_X1   g0037(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n238));
  NOR3_X1   g0038(.A1(new_n224), .A2(new_n237), .A3(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT8), .B(G58), .Z(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n210), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n209), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n202), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n261), .B(new_n209), .C1(G1), .C2(new_n210), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n267), .B2(new_n202), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G274), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n271), .ZN(new_n276));
  OR2_X1    g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G223), .A3(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G222), .A3(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G77), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n280), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n273), .B1(new_n230), .B2(new_n276), .C1(new_n287), .C2(new_n275), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n270), .B(new_n289), .C1(new_n290), .C2(new_n288), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(G169), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n288), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n269), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G20), .A2(G77), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT15), .B(G87), .ZN(new_n298));
  INV_X1    g0098(.A(new_n255), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n297), .B1(new_n259), .B2(new_n298), .C1(new_n258), .C2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(new_n262), .ZN(new_n301));
  INV_X1    g0101(.A(new_n264), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n231), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n231), .B2(new_n266), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n273), .B1(new_n276), .B2(new_n232), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n279), .A2(G238), .A3(G1698), .ZN(new_n307));
  INV_X1    g0107(.A(G107), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n279), .A2(new_n281), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n307), .B1(new_n308), .B2(new_n279), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n275), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(G190), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(G200), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n305), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n305), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n314), .A2(new_n294), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AND4_X1   g0122(.A1(new_n292), .A2(new_n296), .A3(new_n317), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G13), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(G1), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(G20), .A3(new_n326), .ZN(new_n327));
  XOR2_X1   g0127(.A(new_n327), .B(KEYINPUT12), .Z(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(G68), .B2(new_n267), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n299), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n259), .A2(new_n231), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n262), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT11), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n333), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n329), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n279), .A2(G1698), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n338), .B1(new_n309), .B2(new_n230), .C1(new_n310), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n312), .ZN(new_n341));
  INV_X1    g0141(.A(new_n276), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(G238), .B1(G274), .B2(new_n272), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n345), .A2(KEYINPUT66), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n344), .B(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G179), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n345), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n341), .A2(KEYINPUT13), .A3(new_n343), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(G169), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT67), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT14), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n351), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n337), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n337), .B1(new_n347), .B2(G190), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n349), .A2(G200), .A3(new_n350), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n323), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n277), .A2(new_n210), .A3(new_n278), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n278), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n326), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G58), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(new_n326), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n201), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n255), .A2(G159), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT16), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n285), .B2(new_n210), .ZN(new_n376));
  NOR4_X1   g0176(.A1(new_n283), .A2(new_n284), .A3(new_n366), .A4(G20), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(new_n374), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n262), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n257), .A2(new_n266), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n302), .B2(new_n257), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT68), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n273), .B1(new_n276), .B2(new_n310), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n279), .A2(G223), .A3(new_n281), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G87), .ZN(new_n391));
  OAI211_X1 g0191(.A(G226), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n393), .B2(new_n312), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(G169), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n395), .B1(new_n294), .B2(new_n394), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT18), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n388), .A2(new_n399), .A3(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(new_n312), .ZN(new_n402));
  INV_X1    g0202(.A(new_n389), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n290), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G200), .B2(new_n394), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n383), .A2(new_n405), .A3(new_n387), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT17), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT69), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(KEYINPUT69), .A3(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n406), .A2(KEYINPUT17), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n401), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OR3_X1    g0214(.A1(new_n364), .A2(KEYINPUT70), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT70), .B1(new_n364), .B2(new_n414), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G41), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n214), .A2(G45), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT71), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G41), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n214), .A4(G45), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n422), .A2(G41), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(G270), .A3(new_n275), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n214), .B(G45), .C1(new_n418), .C2(KEYINPUT5), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n430), .B2(KEYINPUT71), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n275), .A2(G274), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n425), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(KEYINPUT75), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n279), .A2(G257), .A3(new_n281), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n285), .A2(G303), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(new_n436), .C1(new_n339), .C2(new_n220), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n312), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT75), .B1(new_n429), .B2(new_n433), .ZN(new_n440));
  INV_X1    g0240(.A(G116), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n214), .A2(new_n441), .A3(G13), .A4(G20), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n214), .A2(G33), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n264), .A2(new_n446), .A3(new_n209), .A4(new_n261), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n444), .A2(new_n445), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(new_n210), .C1(G33), .C2(new_n227), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n441), .A2(G20), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n262), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT20), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n448), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR4_X1   g0256(.A1(new_n439), .A2(new_n440), .A3(new_n456), .A4(new_n294), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n455), .ZN(new_n458));
  INV_X1    g0258(.A(new_n448), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n320), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT21), .B(new_n460), .C1(new_n439), .C2(new_n440), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT77), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT75), .ZN(new_n464));
  INV_X1    g0264(.A(G270), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n465), .B(new_n312), .C1(new_n431), .C2(new_n425), .ZN(new_n466));
  INV_X1    g0266(.A(new_n433), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n434), .A3(new_n438), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT77), .A3(KEYINPUT21), .A4(new_n460), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n457), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT21), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(new_n460), .C1(new_n439), .C2(new_n440), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n469), .B2(new_n460), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n439), .A2(new_n440), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G200), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n469), .A2(G190), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n456), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n471), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n262), .ZN(new_n483));
  NAND3_X1  g0283(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n210), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G87), .A2(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n308), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT19), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n485), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n210), .B(G68), .C1(new_n283), .C2(new_n284), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n483), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n447), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT73), .A3(G87), .ZN(new_n495));
  INV_X1    g0295(.A(new_n298), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n264), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT73), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n447), .B2(new_n226), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n493), .A2(new_n495), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  OAI21_X1  g0302(.A(G250), .B1(new_n502), .B2(G1), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n214), .A2(G45), .A3(G274), .ZN(new_n504));
  INV_X1    g0304(.A(new_n209), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n274), .ZN(new_n506));
  OAI211_X1 g0306(.A(G238), .B(new_n281), .C1(new_n283), .C2(new_n284), .ZN(new_n507));
  OAI211_X1 g0307(.A(G244), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G116), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n510), .B2(new_n312), .ZN(new_n511));
  INV_X1    g0311(.A(G200), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(new_n290), .B(new_n506), .C1(new_n510), .C2(new_n312), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n501), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n511), .A2(G169), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n447), .A2(new_n298), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n492), .A2(new_n497), .A3(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(G179), .B(new_n506), .C1(new_n510), .C2(new_n312), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT74), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n428), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n312), .B1(new_n431), .B2(new_n425), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n432), .B1(new_n523), .B2(G257), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G1698), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(G244), .C1(new_n284), .C2(new_n283), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n232), .B1(new_n277), .B2(new_n278), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n449), .C1(new_n528), .C2(KEYINPUT4), .ZN(new_n529));
  OAI21_X1  g0329(.A(G250), .B1(new_n283), .B2(new_n284), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n281), .B1(new_n530), .B2(KEYINPUT4), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n312), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n524), .A2(new_n294), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n523), .A2(G257), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n433), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n320), .ZN(new_n536));
  OAI21_X1  g0336(.A(G107), .B1(new_n376), .B2(new_n377), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  AND2_X1   g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n308), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n483), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n264), .A2(G97), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n494), .B2(G97), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n545), .A2(KEYINPUT72), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT72), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n308), .A2(KEYINPUT6), .A3(G97), .ZN(new_n551));
  XNOR2_X1  g0351(.A(G97), .B(G107), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n538), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n553), .A2(new_n210), .B1(new_n231), .B2(new_n299), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n308), .B1(new_n367), .B2(new_n368), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n262), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n550), .B1(new_n556), .B2(new_n547), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n533), .B(new_n536), .C1(new_n549), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n510), .A2(new_n312), .ZN(new_n559));
  INV_X1    g0359(.A(new_n506), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n320), .ZN(new_n562));
  INV_X1    g0362(.A(new_n517), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n493), .A2(new_n498), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n511), .A2(new_n294), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT74), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n511), .A2(G190), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n512), .B2(new_n511), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n566), .B(new_n567), .C1(new_n501), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n556), .A2(new_n547), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n535), .A2(G190), .ZN(new_n573));
  AOI21_X1  g0373(.A(G200), .B1(new_n524), .B2(new_n532), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n521), .A2(new_n558), .A3(new_n570), .A4(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G250), .B(new_n281), .C1(new_n283), .C2(new_n284), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n578));
  XOR2_X1   g0378(.A(KEYINPUT81), .B(G294), .Z(new_n579));
  INV_X1    g0379(.A(G33), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n312), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n428), .A2(G264), .A3(new_n275), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n433), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G169), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT82), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n523), .A2(KEYINPUT82), .A3(G264), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n433), .A4(new_n582), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n585), .B1(new_n589), .B2(new_n294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n325), .A2(G20), .A3(new_n308), .ZN(new_n591));
  NOR2_X1   g0391(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n592));
  XOR2_X1   g0392(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND2_X1  g0393(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n593), .A2(new_n594), .B1(G107), .B2(new_n494), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n279), .A2(new_n210), .A3(G87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT22), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n279), .A2(new_n598), .A3(new_n210), .A4(G87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT79), .B1(new_n210), .B2(G107), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n600), .A2(KEYINPUT24), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n262), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT24), .B1(new_n600), .B2(new_n606), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n595), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n590), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n584), .A2(G190), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n512), .B2(new_n589), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n576), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n417), .A2(new_n482), .A3(new_n615), .ZN(G372));
  AND2_X1   g0416(.A1(new_n558), .A2(new_n575), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n613), .A2(new_n610), .ZN(new_n618));
  INV_X1    g0418(.A(new_n515), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT84), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n617), .A2(KEYINPUT84), .A3(new_n618), .A4(new_n619), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n471), .A2(new_n477), .A3(new_n611), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n516), .A2(KEYINPUT83), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n518), .A2(new_n519), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n516), .A2(KEYINPUT83), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n521), .A2(new_n570), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(new_n558), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n536), .A2(new_n533), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT85), .B1(new_n635), .B2(new_n571), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n536), .A2(new_n533), .A3(KEYINPUT85), .A4(new_n571), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n629), .A2(new_n637), .A3(new_n619), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n630), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n625), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n417), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n400), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n399), .B1(new_n388), .B2(new_n396), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n359), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n353), .A3(new_n348), .ZN(new_n647));
  INV_X1    g0447(.A(new_n322), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n337), .B1(new_n363), .B2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n406), .A2(KEYINPUT69), .A3(KEYINPUT17), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT69), .B1(new_n406), .B2(KEYINPUT17), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n412), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n645), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n292), .B1(new_n269), .B2(new_n295), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n642), .A2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(new_n325), .ZN(new_n657));
  OR3_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .A3(G20), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT27), .B1(new_n657), .B2(G20), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n456), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n482), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n471), .A2(new_n477), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n610), .A2(new_n662), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n614), .A2(new_n669), .B1(new_n611), .B2(new_n663), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n666), .A2(new_n662), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n590), .A2(new_n610), .A3(new_n663), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(G399));
  NOR2_X1   g0480(.A1(new_n218), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G1), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n486), .A2(new_n308), .A3(new_n441), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT87), .Z(new_n685));
  OAI22_X1  g0485(.A1(new_n683), .A2(new_n685), .B1(new_n207), .B2(new_n682), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n662), .B1(new_n625), .B2(new_n640), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n632), .A2(new_n634), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT26), .B1(new_n636), .B2(new_n638), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n629), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n620), .B1(new_n666), .B2(new_n611), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT29), .B(new_n663), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n532), .A2(new_n433), .A3(new_n534), .A4(new_n511), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n587), .A2(new_n582), .A3(new_n588), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n478), .A3(KEYINPUT30), .A4(G179), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n511), .A2(G179), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n469), .A2(new_n589), .A3(new_n535), .A4(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n469), .A2(new_n294), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n698), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT88), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n699), .A2(new_n701), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT30), .B1(new_n703), .B2(new_n698), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT88), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n662), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n666), .A2(new_n615), .A3(new_n481), .A4(new_n663), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT89), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT31), .B(new_n662), .C1(new_n708), .C2(new_n709), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n482), .A2(KEYINPUT89), .A3(new_n615), .A4(new_n663), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n714), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n695), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n687), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n324), .A2(G20), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G45), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT90), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT90), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n681), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n218), .A2(new_n285), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n732), .A2(G355), .B1(new_n441), .B2(new_n218), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n208), .A2(G45), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n250), .B2(G45), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n218), .A2(new_n279), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n320), .A2(KEYINPUT91), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n320), .A2(KEYINPUT91), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n210), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n209), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n731), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n210), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n512), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n285), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n756), .A2(G329), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n210), .A2(new_n290), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n294), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n753), .B(new_n757), .C1(G322), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n579), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n210), .B1(new_n754), .B2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n294), .A2(new_n512), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n749), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT93), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n767), .A2(new_n758), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n749), .A2(new_n759), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n758), .A2(new_n750), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(G303), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n762), .A2(new_n766), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G58), .A2(new_n761), .B1(new_n779), .B2(G87), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n765), .A2(G97), .ZN(new_n783));
  INV_X1    g0583(.A(new_n768), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n285), .B1(new_n784), .B2(G68), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n755), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  INV_X1    g0589(.A(new_n775), .ZN(new_n790));
  INV_X1    g0590(.A(new_n751), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G77), .A2(new_n790), .B1(new_n791), .B2(G107), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n789), .B(new_n792), .C1(new_n202), .C2(new_n773), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n781), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n748), .B1(new_n742), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n745), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n667), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT94), .Z(new_n798));
  NOR2_X1   g0598(.A1(new_n667), .A2(G330), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n668), .A2(new_n731), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n641), .A2(new_n663), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n317), .B(new_n322), .C1(new_n305), .C2(new_n663), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n648), .B2(new_n662), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT97), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n803), .B(KEYINPUT96), .Z(new_n808));
  NAND2_X1  g0608(.A1(new_n648), .A2(new_n662), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n688), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n806), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n807), .B2(new_n806), .ZN(new_n813));
  INV_X1    g0613(.A(new_n721), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n731), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(KEYINPUT98), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(KEYINPUT98), .B2(new_n816), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n778), .A2(new_n308), .B1(new_n755), .B2(new_n776), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n751), .A2(new_n226), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n819), .A2(new_n279), .A3(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G294), .A2(new_n761), .B1(new_n790), .B2(G116), .ZN(new_n822));
  XOR2_X1   g0622(.A(KEYINPUT95), .B(G283), .Z(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n773), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n784), .A2(new_n824), .B1(new_n825), .B2(G303), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n821), .A2(new_n783), .A3(new_n822), .A4(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n825), .A2(G137), .B1(new_n790), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G143), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n760), .C1(new_n830), .C2(new_n768), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n279), .B1(new_n778), .B2(new_n202), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n751), .A2(new_n326), .B1(new_n755), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(G58), .C2(new_n765), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n831), .A2(new_n832), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n827), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n742), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n742), .A2(new_n743), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n731), .B1(new_n231), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(new_n810), .C2(new_n744), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n818), .A2(new_n844), .ZN(G384));
  OAI211_X1 g0645(.A(G116), .B(new_n211), .C1(new_n543), .C2(KEYINPUT35), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(KEYINPUT35), .B2(new_n543), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT36), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n207), .A2(new_n231), .A3(new_n371), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT99), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n849), .A2(KEYINPUT99), .B1(new_n202), .B2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n214), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  INV_X1    g0655(.A(new_n660), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n388), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(KEYINPUT101), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n397), .A2(new_n857), .A3(new_n406), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n858), .B(new_n859), .Z(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(new_n652), .B2(new_n645), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n383), .A2(new_n385), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n396), .B2(new_n856), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n386), .B1(new_n262), .B2(new_n382), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n855), .B1(new_n865), .B2(new_n405), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n859), .A2(new_n855), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n856), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n867), .C1(new_n413), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n652), .B2(new_n645), .ZN(new_n872));
  INV_X1    g0672(.A(new_n867), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n854), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n869), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n647), .A2(new_n337), .A3(new_n663), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n688), .A2(new_n810), .B1(new_n648), .B2(new_n663), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT100), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n360), .B2(new_n663), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n647), .A2(KEYINPUT100), .A3(new_n337), .A4(new_n662), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n337), .A2(new_n662), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n360), .A2(new_n363), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n875), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n401), .A2(new_n660), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n879), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n417), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n655), .B1(new_n892), .B2(new_n695), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n891), .B(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(G330), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT31), .B(new_n662), .C1(new_n707), .C2(new_n711), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n714), .A2(new_n717), .A3(new_n719), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n417), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(new_n810), .A3(new_n886), .A4(new_n875), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n862), .B2(new_n869), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n902), .A2(new_n810), .A3(new_n897), .A4(new_n886), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n898), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n894), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n214), .B2(new_n725), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n894), .A2(new_n895), .A3(new_n905), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n853), .B1(new_n907), .B2(new_n908), .ZN(G367));
  OAI21_X1  g0709(.A(new_n678), .B1(new_n677), .B2(KEYINPUT42), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n617), .B1(new_n572), .B2(new_n663), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n635), .A2(new_n571), .A3(new_n662), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT103), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n676), .A2(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n917), .B(new_n919), .C1(new_n558), .C2(new_n662), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n629), .A2(new_n501), .A3(new_n662), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n629), .A2(new_n619), .B1(new_n501), .B2(new_n662), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT102), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n925), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n672), .A2(new_n916), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n928), .B(new_n929), .Z(new_n930));
  XOR2_X1   g0730(.A(new_n681), .B(KEYINPUT41), .Z(new_n931));
  NOR2_X1   g0731(.A1(new_n679), .A2(new_n916), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n679), .A2(new_n916), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n935));
  XNOR2_X1  g0735(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n673), .A2(KEYINPUT105), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n668), .A2(new_n671), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n675), .B1(new_n940), .B2(new_n672), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n677), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n722), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n938), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n931), .B1(new_n945), .B2(new_n723), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n930), .B1(new_n946), .B2(new_n729), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n737), .A2(new_n246), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n745), .B(new_n742), .C1(new_n218), .C2(new_n496), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n731), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n779), .A2(KEYINPUT46), .A3(G116), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT46), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n778), .B2(new_n441), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(new_n579), .C2(new_n768), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT106), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n285), .B1(new_n764), .B2(new_n308), .C1(new_n823), .C2(new_n775), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n773), .A2(new_n776), .B1(new_n755), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(G303), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n760), .A2(new_n960), .B1(new_n751), .B2(new_n227), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n957), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT107), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n764), .A2(new_n326), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n285), .B(new_n965), .C1(G150), .C2(new_n761), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n768), .A2(new_n787), .B1(new_n751), .B2(new_n231), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n773), .A2(new_n829), .B1(new_n775), .B2(new_n202), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(G137), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n778), .A2(new_n370), .B1(new_n755), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n966), .A2(new_n969), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n964), .A2(KEYINPUT47), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n742), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT47), .B1(new_n964), .B2(new_n974), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n950), .B1(new_n796), .B2(new_n923), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n947), .A2(new_n978), .ZN(G387));
  INV_X1    g0779(.A(new_n942), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n671), .A2(new_n745), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n257), .A2(new_n202), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT50), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n502), .B1(new_n326), .B2(new_n231), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n983), .A2(new_n685), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n736), .B1(new_n243), .B2(new_n502), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n732), .A2(new_n685), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n217), .A2(G107), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n746), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n730), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G50), .A2(new_n761), .B1(new_n756), .B2(G150), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n992), .B(new_n279), .C1(new_n227), .C2(new_n751), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n258), .A2(new_n768), .B1(new_n326), .B2(new_n775), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n773), .A2(new_n787), .B1(new_n778), .B2(new_n231), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n764), .A2(new_n298), .ZN(new_n996));
  NOR4_X1   g0796(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n763), .A2(new_n779), .B1(new_n824), .B2(new_n765), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n825), .A2(G322), .B1(new_n790), .B2(G303), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n776), .B2(new_n768), .C1(new_n958), .C2(new_n760), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT48), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT109), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n285), .B1(new_n755), .B2(new_n774), .C1(new_n441), .C2(new_n751), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n1006), .B2(KEYINPUT49), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n997), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n742), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1010), .B2(KEYINPUT110), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n991), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n980), .A2(new_n729), .B1(new_n981), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n943), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n681), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n980), .A2(new_n723), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(G393));
  NAND2_X1  g0819(.A1(new_n937), .A2(new_n673), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n933), .A2(new_n672), .A3(new_n936), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n1016), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n945), .A2(new_n1022), .A3(new_n681), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n729), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n916), .A2(new_n796), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n737), .A2(new_n253), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n746), .B1(new_n227), .B2(new_n217), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n730), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G50), .A2(new_n784), .B1(new_n756), .B2(G143), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n326), .B2(new_n778), .C1(new_n258), .C2(new_n775), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n764), .A2(new_n231), .ZN(new_n1032));
  NOR4_X1   g0832(.A1(new_n1031), .A2(new_n285), .A3(new_n820), .A4(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n773), .A2(new_n830), .B1(new_n760), .B2(new_n787), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT51), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n773), .A2(new_n958), .B1(new_n760), .B2(new_n776), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT52), .Z(new_n1037));
  AOI22_X1  g0837(.A1(new_n784), .A2(G303), .B1(new_n765), .B2(G116), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(KEYINPUT111), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n285), .B1(new_n751), .B2(new_n308), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n790), .B1(new_n756), .B2(G322), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n778), .B2(new_n823), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1033), .A2(new_n1035), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT112), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1012), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1029), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1025), .B1(new_n1026), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1023), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(G390));
  NOR2_X1   g0853(.A1(new_n898), .A2(new_n895), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n893), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n897), .A2(G330), .A3(new_n810), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n887), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT114), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n814), .A2(new_n810), .A3(new_n886), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(KEYINPUT114), .A3(new_n887), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n663), .B(new_n804), .C1(new_n692), .C2(new_n693), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n648), .A2(new_n663), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT113), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1062), .A2(KEYINPUT113), .A3(new_n1063), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1056), .A2(new_n887), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n887), .B1(new_n721), .B2(new_n805), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1069), .B1(new_n1072), .B2(new_n880), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1055), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n878), .B1(new_n880), .B2(new_n887), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n877), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1066), .A2(new_n886), .A3(new_n1067), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n870), .A2(new_n878), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1076), .B(new_n1060), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1079), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n877), .A2(new_n1075), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1070), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n682), .B1(new_n1074), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1074), .B2(new_n1083), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n731), .B1(new_n258), .B2(new_n842), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n835), .A2(new_n760), .B1(new_n768), .B2(new_n970), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT54), .B(G143), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n825), .A2(G128), .B1(new_n790), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(G125), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n755), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1087), .B(new_n1092), .C1(G159), .C2(new_n765), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n779), .A2(G150), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n279), .B1(new_n751), .B2(new_n202), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(KEYINPUT116), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1096), .A2(KEYINPUT116), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n285), .B1(new_n778), .B2(new_n226), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT117), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n773), .A2(new_n752), .B1(new_n775), .B2(new_n227), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n308), .A2(new_n768), .B1(new_n760), .B2(new_n441), .ZN(new_n1103));
  INV_X1    g0903(.A(G294), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n751), .A2(new_n326), .B1(new_n755), .B2(new_n1104), .ZN(new_n1105));
  NOR4_X1   g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .A4(new_n1032), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1093), .A2(new_n1099), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1086), .B1(new_n1107), .B2(new_n1012), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n877), .B2(new_n743), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1080), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1082), .A2(new_n1070), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(KEYINPUT115), .A3(new_n729), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1083), .B2(new_n1024), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1109), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1085), .A2(new_n1116), .ZN(G378));
  OAI22_X1  g0917(.A1(new_n773), .A2(new_n1091), .B1(new_n768), .B2(new_n835), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1089), .A2(new_n779), .B1(new_n761), .B2(G128), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n970), .B2(new_n775), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(G150), .C2(new_n765), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n580), .B(new_n418), .C1(new_n751), .C2(new_n787), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G124), .B2(new_n756), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G77), .A2(new_n779), .B1(new_n784), .B2(G97), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n825), .A2(G116), .B1(new_n791), .B2(G58), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n279), .A2(G41), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n308), .B2(new_n760), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n775), .A2(new_n298), .B1(new_n755), .B2(new_n752), .ZN(new_n1133));
  NOR4_X1   g0933(.A1(new_n1130), .A2(new_n965), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(KEYINPUT58), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1134), .A2(KEYINPUT58), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G50), .B(new_n1131), .C1(new_n580), .C2(new_n418), .ZN(new_n1137));
  NOR4_X1   g0937(.A1(new_n1127), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1138), .A2(KEYINPUT118), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1012), .B1(new_n1138), .B2(KEYINPUT118), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n731), .B(new_n1141), .C1(new_n202), .C2(new_n842), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n292), .A2(new_n296), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n269), .A2(new_n856), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1143), .B(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n743), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n891), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n901), .A2(G330), .A3(new_n903), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(new_n1147), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1147), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT119), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(new_n1156), .A3(new_n1147), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1153), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT120), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1151), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1152), .A2(new_n1147), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1152), .A2(new_n1156), .A3(new_n1147), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1156), .B1(new_n1152), .B2(new_n1147), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(KEYINPUT120), .A3(new_n891), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1150), .B1(new_n1166), .B2(new_n729), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1073), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1055), .B1(new_n1168), .B2(new_n1083), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT57), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1164), .A2(new_n1151), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n891), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1171), .A3(KEYINPUT57), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n681), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1167), .B1(new_n1170), .B2(new_n1174), .ZN(G375));
  NAND2_X1  g0975(.A1(new_n887), .A2(new_n743), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n778), .A2(new_n227), .B1(new_n755), .B2(new_n960), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT121), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G116), .A2(new_n784), .B1(new_n790), .B2(G107), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n279), .B(new_n996), .C1(G77), .C2(new_n791), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G294), .A2(new_n825), .B1(new_n761), .B2(G283), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n279), .B1(new_n751), .B2(new_n370), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G150), .A2(new_n790), .B1(new_n756), .B2(G128), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n787), .B2(new_n778), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(G50), .C2(new_n765), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT122), .Z(new_n1187));
  AOI22_X1  g0987(.A1(G132), .A2(new_n825), .B1(new_n784), .B2(new_n1089), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n970), .B2(new_n760), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(new_n742), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n731), .B(new_n1191), .C1(new_n326), .C2(new_n842), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1073), .A2(new_n729), .B1(new_n1176), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n931), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1074), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1055), .A2(new_n1073), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1193), .B1(new_n1195), .B2(new_n1196), .ZN(G381));
  NAND3_X1  g0997(.A1(new_n947), .A2(new_n1052), .A3(new_n978), .ZN(new_n1198));
  OR2_X1    g0998(.A1(G393), .A2(G396), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1198), .A2(G384), .A3(G381), .A4(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(G375), .A2(G378), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(G407));
  INV_X1    g1003(.A(G213), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(G343), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(G407), .A2(G213), .A3(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1008(.A(KEYINPUT62), .ZN(new_n1209));
  INV_X1    g1009(.A(G384), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1074), .A2(new_n681), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT60), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1196), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT60), .B1(new_n1055), .B2(new_n1073), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1193), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1210), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n682), .B1(new_n1055), .B2(new_n1073), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1214), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1055), .A2(new_n1073), .A3(KEYINPUT60), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(G384), .A3(new_n1193), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1217), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1171), .A2(new_n729), .A3(new_n1172), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1149), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(KEYINPUT124), .A3(new_n1149), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1166), .A2(new_n1194), .A3(new_n1169), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G378), .B(new_n1167), .C1(new_n1170), .C2(new_n1174), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1205), .B(new_n1223), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT127), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1209), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1205), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1223), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1112), .A2(new_n1073), .A3(new_n1055), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1160), .A2(new_n1165), .B1(new_n1239), .B2(new_n1055), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1240), .A2(new_n1194), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G378), .B1(new_n1241), .B2(new_n1228), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1233), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1237), .B(new_n1238), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1205), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1205), .A2(G2897), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1223), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1217), .A2(new_n1222), .A3(new_n1248), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(KEYINPUT126), .B(new_n1246), .C1(new_n1247), .C2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1236), .A2(new_n1245), .A3(new_n1253), .ZN(new_n1254));
  XOR2_X1   g1054(.A(G393), .B(G396), .Z(new_n1255));
  AND3_X1   g1055(.A1(new_n947), .A2(new_n1052), .A3(new_n978), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1052), .B1(new_n947), .B2(new_n978), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(G390), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1255), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1198), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1237), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1262), .B1(new_n1265), .B2(KEYINPUT126), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1254), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(KEYINPUT125), .A3(new_n1264), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1234), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1244), .A2(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1262), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1267), .A2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(new_n1262), .A2(new_n1223), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1258), .A2(new_n1261), .A3(new_n1238), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(G375), .B(new_n1231), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1278), .A2(new_n1281), .A3(new_n1279), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(G402));
endmodule


