//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(new_n466), .B1(G101), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n461), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT67), .B(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n473), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n461), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G124), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n459), .B2(new_n460), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G138), .B1(new_n459), .B2(new_n460), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT4), .B1(new_n491), .B2(new_n473), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n466), .A2(new_n477), .A3(new_n493), .A4(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G50), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n498), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n502), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n500), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n502), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(new_n503), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT68), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n508), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(new_n499), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n504), .A2(new_n502), .ZN(new_n522));
  OAI21_X1  g097(.A(G89), .B1(new_n505), .B2(new_n506), .ZN(new_n523));
  NAND2_X1  g098(.A1(G63), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n526));
  OR3_X1    g101(.A1(new_n521), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n521), .B2(new_n525), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(new_n499), .A2(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n507), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT70), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT70), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n522), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n533), .A2(new_n534), .B1(G651), .B2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n522), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n509), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n543), .B1(new_n542), .B2(new_n541), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n510), .A2(new_n503), .B1(new_n497), .B2(new_n498), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G81), .B1(new_n499), .B2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n499), .A2(G53), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(KEYINPUT72), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n554), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n522), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n545), .B2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(new_n533), .A2(new_n534), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n537), .A2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  OR3_X1    g142(.A1(new_n504), .A2(new_n502), .A3(G74), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(new_n499), .B2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n545), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G288));
  OAI211_X1 g146(.A(G48), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n507), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n504), .B2(new_n502), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n509), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n509), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n499), .A2(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n507), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(new_n545), .A2(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n522), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n499), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n595), .B2(G171), .ZN(G284));
  OAI21_X1  g172(.A(new_n596), .B1(new_n595), .B2(G171), .ZN(G321));
  NOR2_X1   g173(.A1(G299), .A2(G868), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g175(.A(new_n599), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g176(.A(new_n594), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n477), .A2(new_n468), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(G2100), .ZN(new_n614));
  OAI221_X1 g189(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n480), .A2(G135), .ZN(new_n616));
  INV_X1    g191(.A(G123), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n478), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(G156));
  XOR2_X1   g195(.A(G1341), .B(G1348), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT74), .ZN(new_n622));
  XOR2_X1   g197(.A(G2451), .B(G2454), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n622), .B(new_n624), .Z(new_n625));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n625), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(G14), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT75), .Z(G401));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT76), .ZN(new_n639));
  NOR2_X1   g214(.A1(G2072), .A2(G2078), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n442), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n639), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT18), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n641), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n641), .B(KEYINPUT17), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n646), .B(new_n643), .C1(new_n639), .C2(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n639), .A3(new_n642), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT77), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(KEYINPUT78), .B(KEYINPUT19), .Z(new_n654));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT79), .Z(new_n661));
  AND2_X1   g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n656), .A2(new_n662), .A3(new_n659), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  MUX2_X1   g247(.A(G23), .B(G288), .S(G16), .Z(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT33), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G22), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G166), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G1971), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n578), .B2(G16), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n677), .A2(new_n678), .A3(new_n683), .A4(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT82), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT82), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(KEYINPUT34), .A3(new_n690), .ZN(new_n694));
  INV_X1    g269(.A(G24), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n695), .A2(KEYINPUT80), .A3(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT80), .B1(new_n695), .B2(G16), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n696), .B(new_n697), .C1(new_n585), .C2(new_n679), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1986), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n479), .A2(G119), .B1(new_n480), .B2(G131), .ZN(new_n700));
  OAI221_X1 g275(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  AOI211_X1 g280(.A(new_n699), .B(new_n705), .C1(KEYINPUT83), .C2(KEYINPUT36), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n693), .A2(new_n694), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G21), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G168), .B2(G16), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT94), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT95), .B(G1966), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT96), .Z(new_n715));
  NOR2_X1   g290(.A1(G171), .A2(new_n679), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G5), .B2(new_n679), .ZN(new_n717));
  INV_X1    g292(.A(G1961), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT97), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n618), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT30), .B(G28), .ZN(new_n723));
  OR2_X1    g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  NAND2_X1  g299(.A1(KEYINPUT31), .A2(G11), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n723), .A2(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n712), .B2(new_n713), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n715), .A2(new_n720), .A3(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT98), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n707), .A2(new_n708), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n721), .A2(G26), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n479), .A2(G128), .ZN(new_n734));
  OR2_X1    g309(.A1(G104), .A2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n467), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n737), .B1(new_n736), .B2(new_n735), .C1(G116), .C2(new_n466), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n480), .A2(G140), .ZN(new_n739));
  AND3_X1   g314(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2067), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n721), .B1(new_n745), .B2(G34), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(KEYINPUT89), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(KEYINPUT89), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n475), .A2(new_n721), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n602), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G4), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n468), .A2(G105), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT91), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G141), .B2(new_n480), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n479), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(new_n721), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n721), .B2(G32), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT92), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n752), .B1(new_n754), .B2(new_n755), .C1(new_n765), .C2(new_n768), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n744), .B(new_n769), .C1(new_n755), .C2(new_n754), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n721), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n721), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT29), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G2090), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT99), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n548), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT84), .B(G1341), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n717), .A2(new_n718), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n779), .B(new_n780), .C1(G2090), .C2(new_n773), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n679), .A2(G20), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT23), .Z(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n721), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n721), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2078), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n770), .A2(new_n775), .A3(new_n781), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n750), .A2(new_n751), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT90), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n765), .A2(new_n768), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n480), .A2(G139), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n797), .B(new_n798), .C1(new_n466), .C2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT86), .ZN(new_n801));
  MUX2_X1   g376(.A(G33), .B(new_n801), .S(G29), .Z(new_n802));
  AOI211_X1 g377(.A(new_n793), .B(new_n794), .C1(G2072), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(G2072), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT87), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n803), .A2(KEYINPUT93), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(KEYINPUT93), .B1(new_n803), .B2(new_n805), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n791), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AND4_X1   g383(.A1(new_n709), .A2(new_n730), .A3(new_n731), .A4(new_n808), .ZN(G311));
  NAND4_X1  g384(.A1(new_n730), .A2(new_n808), .A3(new_n709), .A4(new_n731), .ZN(G150));
  NAND2_X1  g385(.A1(new_n602), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT38), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n545), .A2(G93), .B1(new_n499), .B2(G55), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n509), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n547), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n547), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n812), .B(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n821), .A2(new_n822), .A3(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n815), .A2(G860), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n823), .A2(new_n825), .ZN(G145));
  INV_X1    g401(.A(G37), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n801), .B(new_n763), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n740), .B(G164), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n479), .A2(G130), .B1(new_n480), .B2(G142), .ZN(new_n833));
  OAI221_X1 g408(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n610), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n702), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT100), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n618), .B(new_n475), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n483), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n837), .A2(KEYINPUT100), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n830), .A2(new_n842), .A3(new_n831), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n839), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n841), .B1(new_n839), .B2(new_n843), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g422(.A(KEYINPUT101), .B(new_n841), .C1(new_n839), .C2(new_n843), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n827), .B(new_n844), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(G395));
  NAND2_X1  g426(.A1(new_n815), .A2(new_n595), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n557), .A2(new_n561), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g430(.A1(G299), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n602), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n594), .A2(new_n855), .A3(G299), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n857), .A2(KEYINPUT41), .A3(new_n858), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n818), .B(new_n605), .Z(new_n864));
  MUX2_X1   g439(.A(new_n860), .B(new_n863), .S(new_n864), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT42), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n585), .B(new_n578), .ZN(new_n867));
  XNOR2_X1  g442(.A(G166), .B(G288), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n866), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n852), .B1(new_n871), .B2(new_n595), .ZN(G295));
  OAI21_X1  g447(.A(new_n852), .B1(new_n871), .B2(new_n595), .ZN(G331));
  NAND2_X1  g448(.A1(G286), .A2(G301), .ZN(new_n874));
  NAND2_X1  g449(.A1(G171), .A2(G168), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n818), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n874), .A2(new_n817), .A3(new_n816), .A4(new_n875), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(KEYINPUT104), .A3(new_n818), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n860), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(KEYINPUT105), .A3(new_n860), .ZN(new_n886));
  INV_X1    g461(.A(new_n879), .ZN(new_n887));
  INV_X1    g462(.A(new_n877), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n863), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n885), .A2(new_n870), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n888), .A2(new_n887), .A3(new_n859), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n880), .A2(new_n863), .A3(new_n881), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n880), .A2(new_n863), .A3(KEYINPUT106), .A4(new_n881), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n870), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n890), .B(new_n827), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  AOI211_X1 g474(.A(KEYINPUT107), .B(new_n870), .C1(new_n894), .C2(new_n895), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n890), .A2(new_n827), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n869), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT43), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT44), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n898), .A2(KEYINPUT43), .A3(new_n900), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n899), .B1(new_n902), .B2(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n906), .B1(new_n909), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g485(.A(new_n490), .ZN(new_n911));
  INV_X1    g486(.A(G138), .ZN(new_n912));
  OR2_X1    g487(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n913));
  NAND2_X1  g488(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n493), .B1(new_n915), .B2(new_n466), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n491), .A2(new_n473), .A3(KEYINPUT4), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(G164), .B2(G1384), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT45), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n469), .A2(G40), .A3(new_n474), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n919), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n713), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n920), .A2(new_n922), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(KEYINPUT50), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n751), .A3(new_n924), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G8), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT51), .ZN(new_n935));
  INV_X1    g510(.A(G8), .ZN(new_n936));
  NOR2_X1   g511(.A1(G168), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n928), .A2(KEYINPUT121), .A3(new_n932), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT121), .B1(new_n928), .B2(new_n932), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(G286), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n936), .B1(KEYINPUT122), .B2(new_n935), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(KEYINPUT122), .B2(new_n935), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n939), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT121), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n933), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n928), .A2(KEYINPUT121), .A3(new_n932), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n938), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n952));
  NAND3_X1  g527(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G166), .B2(new_n936), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n469), .A2(G40), .A3(new_n474), .ZN(new_n958));
  NOR2_X1   g533(.A1(G164), .A2(G1384), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n925), .A2(new_n926), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n682), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n929), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT109), .B1(new_n918), .B2(new_n919), .ZN(new_n966));
  NOR3_X1   g541(.A1(G164), .A2(new_n921), .A3(G1384), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n958), .B1(new_n959), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G2090), .B1(new_n971), .B2(KEYINPUT115), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n964), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n952), .B(new_n957), .C1(new_n975), .C2(new_n936), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n929), .B1(new_n920), .B2(new_n922), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n924), .B1(new_n925), .B2(KEYINPUT50), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT115), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2090), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n936), .B1(new_n981), .B2(new_n963), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT116), .B1(new_n982), .B2(new_n956), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n930), .A2(new_n924), .A3(new_n931), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n963), .B1(G2090), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n956), .B(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n578), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(G1981), .B1(new_n574), .B2(new_n577), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(KEYINPUT49), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n997));
  INV_X1    g572(.A(new_n577), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n545), .A2(G86), .B1(new_n499), .B2(G48), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n574), .A2(new_n577), .A3(G1981), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n992), .A2(G8), .A3(new_n996), .A4(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT113), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n569), .A2(G1976), .A3(new_n570), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT112), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(G8), .A3(new_n992), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n992), .A3(G8), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n991), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n996), .A2(new_n1002), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1014), .A2(KEYINPUT113), .A3(G8), .A4(new_n992), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1003), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT117), .A3(new_n1011), .A4(new_n1008), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n990), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n985), .A2(new_n718), .ZN(new_n1021));
  INV_X1    g596(.A(G2078), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n960), .A2(new_n1022), .A3(new_n961), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(G2078), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n474), .A2(G40), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(new_n469), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n469), .A2(new_n1029), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n961), .A2(new_n1026), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1021), .A2(new_n1025), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G171), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n718), .A2(new_n985), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1035));
  INV_X1    g610(.A(new_n923), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(new_n960), .A3(new_n1027), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(G301), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1038), .A3(KEYINPUT54), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n951), .A2(new_n984), .A3(new_n1020), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1033), .A2(G171), .ZN(new_n1042));
  AOI21_X1  g617(.A(G301), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT124), .B(new_n1041), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT125), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n984), .A2(new_n1020), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1039), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n945), .B2(new_n950), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(G299), .B(KEYINPUT57), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n960), .A2(new_n961), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1956), .B1(new_n968), .B2(new_n970), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n992), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n985), .A2(new_n755), .B1(new_n1062), .B2(new_n743), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1063), .B2(new_n594), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n785), .A2(new_n971), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1056), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT61), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT120), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n992), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n962), .B2(G1996), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n548), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT59), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1074), .B(KEYINPUT119), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1063), .A2(KEYINPUT60), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n594), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1063), .A2(KEYINPUT60), .A3(new_n602), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1082), .B(new_n1083), .C1(KEYINPUT60), .C2(new_n1063), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1061), .A2(new_n1067), .A3(KEYINPUT61), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1077), .A2(new_n1080), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1068), .B1(new_n1070), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1049), .A2(new_n1055), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n934), .A2(G286), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n984), .A2(new_n1020), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n984), .A2(new_n1020), .A3(KEYINPUT118), .A4(new_n1089), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n990), .B1(new_n957), .B2(new_n987), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(KEYINPUT63), .A3(new_n1089), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1018), .A2(new_n1009), .A3(new_n570), .A4(new_n569), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n994), .B(KEYINPUT114), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n936), .B(new_n1062), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n990), .B2(new_n1097), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n945), .A2(new_n1105), .A3(new_n950), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1050), .A2(new_n1104), .A3(new_n1106), .A4(new_n1043), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n984), .A2(new_n1020), .A3(new_n1043), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n947), .A2(G168), .A3(new_n948), .ZN(new_n1109));
  INV_X1    g684(.A(new_n944), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT62), .B(new_n949), .C1(new_n1111), .C2(new_n939), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT126), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1088), .A2(new_n1099), .A3(new_n1103), .A4(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n961), .A2(new_n958), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(G1996), .A3(new_n762), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT108), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n740), .B(G2067), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(G1996), .B2(new_n762), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1119), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1117), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n702), .B(new_n704), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(new_n585), .B(G1986), .Z(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1117), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1116), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1123), .B1(new_n1120), .B2(new_n763), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT46), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1123), .A2(G1996), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT47), .Z(new_n1134));
  NAND4_X1  g709(.A1(new_n1122), .A2(new_n704), .A3(new_n701), .A4(new_n700), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n740), .A2(new_n743), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1123), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1123), .A2(G1986), .A3(G290), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT48), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1125), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1134), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1128), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g717(.A(G319), .ZN(new_n1144));
  INV_X1    g718(.A(new_n636), .ZN(new_n1145));
  NOR4_X1   g719(.A1(G229), .A2(new_n1144), .A3(new_n1145), .A4(G227), .ZN(new_n1146));
  OAI211_X1 g720(.A(new_n849), .B(new_n1146), .C1(new_n907), .C2(new_n908), .ZN(G225));
  INV_X1    g721(.A(G225), .ZN(G308));
endmodule


