//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n209), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(new_n212), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n207), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n223), .A2(new_n226), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  XOR2_X1   g0034(.A(G226), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(G87), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n202), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n230), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT67), .A2(G58), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT8), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n207), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n252), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n216), .ZN(new_n266));
  INV_X1    g0066(.A(new_n252), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G1), .B2(new_n207), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n263), .B(new_n266), .C1(new_n216), .C2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G226), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OR2_X1    g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G222), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G223), .A2(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n291), .B(new_n277), .C1(G77), .C2(new_n287), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n281), .A2(new_n284), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G200), .B2(new_n293), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n270), .A2(new_n273), .A3(new_n274), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n276), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n298), .A2(KEYINPUT70), .A3(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(new_n269), .C1(G179), .C2(new_n293), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n288), .A2(G232), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n287), .B(new_n308), .C1(new_n213), .C2(new_n288), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n277), .C1(G107), .C2(new_n287), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n280), .A2(G244), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n310), .A2(new_n311), .A3(new_n284), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n268), .A2(new_n218), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT8), .B(G58), .Z(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT15), .B(G87), .Z(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n256), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n315), .B1(new_n320), .B2(new_n252), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G77), .B2(new_n264), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n310), .A2(new_n311), .A3(new_n284), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n304), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n314), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n307), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n268), .A2(new_n212), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT71), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n264), .A2(G68), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT12), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT72), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n330), .B2(new_n329), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n261), .A2(new_n216), .B1(new_n207), .B2(G68), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n256), .A2(new_n218), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n252), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT11), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n328), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n217), .A2(new_n288), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n287), .B(new_n339), .C1(G232), .C2(new_n288), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n277), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n278), .A2(G238), .A3(new_n279), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n345), .A3(new_n284), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT13), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n283), .B1(new_n342), .B2(new_n277), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n345), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(G190), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n349), .B1(new_n348), .B2(new_n345), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n278), .B1(new_n340), .B2(new_n341), .ZN(new_n353));
  NOR4_X1   g0153(.A1(new_n353), .A2(new_n344), .A3(KEYINPUT13), .A4(new_n283), .ZN(new_n354));
  OAI21_X1  g0154(.A(G200), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n338), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n338), .A2(new_n351), .A3(new_n355), .A4(KEYINPUT73), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(G169), .B1(new_n352), .B2(new_n354), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT14), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n347), .A2(G179), .A3(new_n350), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(G169), .C1(new_n352), .C2(new_n354), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n328), .A2(new_n333), .A3(new_n337), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n322), .B1(G190), .B2(new_n312), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n312), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n287), .A2(new_n375), .A3(G20), .ZN(new_n376));
  AND2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT3), .A2(G33), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT7), .B1(new_n379), .B2(new_n207), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n260), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n228), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n382), .A4(new_n385), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n252), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G87), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n287), .B1(G226), .B2(new_n288), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G223), .A2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n283), .B1(new_n394), .B2(new_n277), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n280), .A2(G232), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(G190), .A3(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n268), .A2(new_n255), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n255), .A2(new_n265), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n390), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n396), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n371), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n374), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n400), .A2(new_n374), .A3(new_n403), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n390), .A2(new_n398), .A3(new_n399), .ZN(new_n409));
  AOI21_X1  g0209(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(G179), .B2(new_n401), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n408), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n390), .A2(new_n398), .A3(new_n399), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n402), .B2(new_n313), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT18), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT74), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n418), .A2(KEYINPUT74), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n326), .A2(new_n373), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G283), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n379), .A2(new_n219), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(KEYINPUT4), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n287), .A2(G250), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n288), .B1(new_n427), .B2(KEYINPUT4), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n277), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT5), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(G41), .ZN(new_n431));
  INV_X1    g0231(.A(G41), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n206), .B(G45), .C1(new_n432), .C2(KEYINPUT5), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n278), .B(G257), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n277), .A2(new_n282), .A3(new_n431), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n433), .B(KEYINPUT78), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n429), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n304), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n429), .A2(new_n313), .A3(new_n434), .A4(new_n437), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n252), .B(new_n265), .C1(new_n206), .C2(G33), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT77), .B1(new_n264), .B2(G97), .ZN(new_n444));
  OR3_X1    g0244(.A1(new_n264), .A2(KEYINPUT77), .A3(G97), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n443), .A2(G97), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(G97), .B(G107), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT6), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n448), .A2(new_n202), .A3(G107), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n207), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n261), .A2(new_n218), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT75), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(G107), .B1(new_n376), .B2(new_n380), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT75), .ZN(new_n456));
  INV_X1    g0256(.A(new_n453), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n450), .B1(new_n448), .B2(new_n447), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n207), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n460), .A2(KEYINPUT76), .A3(new_n252), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT76), .B1(new_n460), .B2(new_n252), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n446), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n442), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n462), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(KEYINPUT76), .A3(new_n252), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT79), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n294), .B1(new_n468), .B2(new_n371), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n429), .A2(new_n434), .A3(new_n437), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n438), .A2(new_n468), .A3(G200), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n446), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n443), .A2(new_n318), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT19), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n256), .B2(new_n202), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n207), .B(G68), .C1(new_n377), .C2(new_n378), .ZN(new_n476));
  OR2_X1    g0276(.A1(KEYINPUT80), .A2(G87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT80), .A2(G87), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n204), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n207), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n475), .B(new_n476), .C1(new_n479), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n252), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n318), .A2(new_n264), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT81), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT81), .ZN(new_n488));
  AOI211_X1 g0288(.A(new_n488), .B(new_n485), .C1(new_n483), .C2(new_n252), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n473), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G20), .B1(new_n285), .B2(new_n286), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT80), .A2(G87), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT80), .A2(G87), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(G68), .A2(new_n493), .B1(new_n497), .B2(new_n481), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n267), .B1(new_n498), .B2(new_n475), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n488), .B1(new_n499), .B2(new_n485), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n484), .A2(KEYINPUT81), .A3(new_n486), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n473), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n213), .A2(new_n288), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n287), .B(new_n504), .C1(G244), .C2(new_n288), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n278), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G45), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n508), .A2(G1), .A3(G274), .ZN(new_n509));
  AOI21_X1  g0309(.A(G250), .B1(new_n206), .B2(G45), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n277), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G179), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n304), .B2(new_n512), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n492), .A2(new_n503), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n512), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n294), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n443), .A2(G87), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n512), .A2(new_n371), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n518), .A2(new_n502), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  AND4_X1   g0322(.A1(new_n464), .A2(new_n472), .A3(new_n515), .A4(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n207), .A2(G107), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT23), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n506), .A2(G20), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT85), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n493), .B2(G87), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n207), .B(G87), .C1(new_n377), .C2(new_n378), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n525), .B(new_n527), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT86), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n530), .B(KEYINPUT22), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(KEYINPUT86), .A3(new_n525), .A4(new_n527), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT24), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n252), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n443), .A2(G107), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n265), .A2(new_n203), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT87), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n543), .B(KEYINPUT25), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  OR2_X1    g0345(.A1(G250), .A2(G1698), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n287), .B(new_n546), .C1(G257), .C2(new_n288), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT88), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT88), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n277), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n278), .B(G264), .C1(new_n431), .C2(new_n433), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n437), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n304), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n553), .A2(new_n313), .A3(new_n437), .A4(new_n554), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n553), .A2(G190), .A3(new_n437), .A4(new_n554), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n540), .A2(new_n541), .A3(new_n544), .A4(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n555), .A2(G200), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n545), .A2(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT89), .ZN(new_n563));
  INV_X1    g0363(.A(new_n558), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT89), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n561), .C2(new_n560), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n288), .A2(G257), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G264), .A2(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n287), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g0372(.A(KEYINPUT83), .B(G303), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n277), .C1(new_n287), .C2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n278), .B(G270), .C1(new_n431), .C2(new_n433), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n436), .C2(new_n435), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT84), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n437), .A2(new_n579), .A3(new_n576), .A4(new_n575), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n443), .A2(G116), .ZN(new_n582));
  INV_X1    g0382(.A(G116), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n265), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n424), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n252), .C1(new_n207), .C2(G116), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n582), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n581), .A2(KEYINPUT21), .A3(G169), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n577), .A2(new_n313), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n590), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n578), .A2(new_n580), .A3(new_n590), .A4(G169), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n591), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n581), .A2(G200), .ZN(new_n598));
  INV_X1    g0398(.A(new_n590), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n294), .C2(new_n581), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n422), .A2(new_n523), .A3(new_n569), .A4(new_n601), .ZN(new_n602));
  XOR2_X1   g0402(.A(new_n602), .B(KEYINPUT90), .Z(G372));
  AND3_X1   g0403(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n301), .B1(new_n298), .B2(new_n302), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n407), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n366), .A2(new_n367), .B1(new_n356), .B2(new_n325), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n417), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n306), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n514), .A2(new_n490), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT91), .B1(new_n502), .B2(new_n519), .ZN(new_n615));
  OAI211_X1 g0415(.A(KEYINPUT91), .B(new_n519), .C1(new_n487), .C2(new_n489), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n521), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n517), .B1(new_n618), .B2(KEYINPUT92), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n519), .B1(new_n487), .B2(new_n489), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT91), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n520), .B1(new_n622), .B2(new_n616), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT92), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n614), .B1(new_n619), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n560), .A2(new_n561), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n597), .B2(new_n566), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n464), .A2(new_n626), .A3(new_n472), .A4(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n515), .A2(new_n442), .A3(new_n522), .A4(new_n463), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n614), .B1(new_n630), .B2(KEYINPUT26), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n441), .B1(new_n467), .B2(new_n446), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n518), .B1(new_n623), .B2(new_n624), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT92), .B(new_n520), .C1(new_n622), .C2(new_n616), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n632), .B(new_n613), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n631), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT93), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(KEYINPUT93), .B(new_n631), .C1(new_n635), .C2(KEYINPUT26), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n629), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n612), .B1(new_n421), .B2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(G13), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(G20), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n206), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n597), .B(new_n600), .C1(new_n599), .C2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n591), .A2(new_n596), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n590), .B(new_n649), .C1(new_n652), .C2(new_n592), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT94), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT94), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n651), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G330), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n566), .A2(new_n650), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n565), .A2(new_n649), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n660), .B1(new_n569), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n597), .A2(new_n649), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n569), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n564), .A2(new_n565), .A3(new_n650), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n663), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n224), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n479), .A2(new_n583), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n229), .B2(new_n671), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n626), .A2(new_n464), .A3(new_n628), .A4(new_n472), .ZN(new_n677));
  INV_X1    g0477(.A(new_n639), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n618), .A2(KEYINPUT92), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n518), .A3(new_n625), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n632), .A4(new_n613), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT93), .B1(new_n682), .B2(new_n631), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n677), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n650), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n630), .A2(new_n681), .ZN(new_n687));
  OAI211_X1 g0487(.A(KEYINPUT96), .B(new_n687), .C1(new_n635), .C2(new_n681), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT96), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n626), .A2(new_n689), .A3(KEYINPUT26), .A4(new_n632), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT97), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n471), .A2(new_n470), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n463), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n632), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n472), .A2(new_n464), .A3(KEYINPUT97), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n626), .A3(new_n628), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n688), .A2(new_n690), .A3(new_n697), .A4(new_n613), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n650), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n686), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n569), .A2(new_n523), .A3(new_n601), .A4(new_n650), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n553), .A2(new_n512), .A3(new_n554), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT95), .ZN(new_n705));
  INV_X1    g0505(.A(new_n438), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT95), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n553), .A2(new_n707), .A3(new_n512), .A4(new_n554), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n705), .A2(new_n706), .A3(new_n592), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n438), .B1(new_n704), .B2(KEYINPUT95), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n592), .A4(new_n708), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n706), .A2(G179), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n516), .A3(new_n555), .A4(new_n581), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n716), .B2(new_n649), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n702), .B1(new_n703), .B2(new_n719), .ZN(new_n720));
  OR3_X1    g0520(.A1(new_n701), .A2(KEYINPUT98), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT98), .B1(new_n701), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n676), .B1(new_n723), .B2(G1), .ZN(G364));
  NAND2_X1  g0524(.A1(new_n643), .A2(G45), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n671), .A2(G1), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n658), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n230), .B1(G20), .B2(new_n304), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT99), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n735), .A2(G190), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n207), .ZN(new_n737));
  INV_X1    g0537(.A(G294), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G326), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n207), .A2(new_n313), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n371), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n737), .A2(new_n735), .ZN(new_n745));
  INV_X1    g0545(.A(G329), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n379), .B1(new_n740), .B2(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n741), .A2(new_n294), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(KEYINPUT33), .B(G317), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n739), .B(new_n747), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n741), .A2(new_n294), .A3(new_n371), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G311), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G303), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n741), .A2(G190), .A3(new_n371), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n755), .A2(new_n294), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G322), .A2(new_n760), .B1(new_n762), .B2(G283), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n751), .A2(new_n754), .A3(new_n758), .A4(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n745), .ZN(new_n765));
  XOR2_X1   g0565(.A(KEYINPUT100), .B(G159), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT32), .Z(new_n768));
  NAND2_X1  g0568(.A1(new_n762), .A2(G107), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n769), .B(new_n287), .C1(new_n227), .C2(new_n759), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n737), .A2(new_n202), .B1(new_n212), .B2(new_n748), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(G50), .C2(new_n743), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n757), .A2(new_n477), .A3(new_n478), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n753), .A2(G77), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n768), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n764), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n730), .A2(new_n732), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n669), .A2(new_n287), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G45), .B2(new_n229), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n249), .A2(new_n508), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(G116), .B2(new_n224), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n669), .A2(new_n379), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G355), .B2(new_n783), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n731), .B1(new_n733), .B2(new_n776), .C1(new_n778), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n727), .A2(new_n702), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(new_n659), .A3(new_n726), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(G396));
  NAND3_X1  g0588(.A1(new_n314), .A2(new_n322), .A3(new_n324), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n789), .A2(KEYINPUT104), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(KEYINPUT104), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(new_n372), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n684), .A2(new_n650), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n640), .A2(new_n649), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n322), .A2(new_n649), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n372), .B(new_n796), .C1(new_n790), .C2(new_n791), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n325), .A2(new_n649), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n794), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n720), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n703), .A2(new_n719), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G330), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n803), .B(new_n794), .C1(new_n795), .C2(new_n799), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n801), .A2(new_n726), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n737), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G97), .B1(G283), .B2(new_n749), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n379), .B1(new_n756), .B2(new_n203), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(KEYINPUT101), .B2(new_n808), .C1(new_n738), .C2(new_n759), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G311), .B2(new_n765), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n743), .A2(G303), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n762), .A2(G87), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n808), .A2(KEYINPUT101), .B1(new_n753), .B2(G116), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n744), .A2(new_n815), .B1(new_n259), .B2(new_n748), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT102), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n760), .A2(G143), .B1(new_n753), .B2(new_n766), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT103), .Z(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n765), .A2(G132), .B1(G68), .B2(new_n762), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n379), .B1(new_n806), .B2(G58), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(new_n216), .C2(new_n756), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n814), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n732), .A2(new_n728), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n825), .A2(new_n732), .B1(new_n218), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n729), .B2(new_n799), .ZN(new_n828));
  INV_X1    g0628(.A(new_n726), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n805), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(KEYINPUT105), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(KEYINPUT105), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G384));
  NOR2_X1   g0635(.A1(new_n643), .A2(new_n206), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n422), .A2(new_n802), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT109), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n367), .A2(new_n649), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n360), .B2(new_n368), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n356), .A2(new_n839), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n367), .B2(new_n366), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n799), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n647), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n414), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n403), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n848), .A4(new_n397), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT107), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(new_n404), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n417), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n850), .B1(new_n849), .B2(new_n404), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT106), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n414), .B1(new_n415), .B2(new_n845), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n400), .A2(new_n403), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n855), .B(new_n856), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n859), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n856), .ZN(new_n862));
  NAND2_X1  g0662(.A1(KEYINPUT106), .A2(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n854), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n846), .B1(new_n407), .B2(new_n417), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n802), .B(new_n844), .C1(new_n867), .C2(new_n870), .ZN(new_n871));
  AOI211_X1 g0671(.A(KEYINPUT40), .B(new_n843), .C1(new_n703), .C2(new_n719), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n418), .A2(new_n847), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n869), .B1(new_n868), .B2(new_n865), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n871), .A2(KEYINPUT40), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n838), .B(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n702), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT108), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n685), .B1(new_n698), .B2(new_n650), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n795), .B2(new_n685), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n880), .B1(new_n882), .B2(new_n421), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n701), .A2(KEYINPUT108), .A3(new_n422), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n611), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n840), .A2(new_n842), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n793), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n640), .A2(new_n649), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n792), .A2(new_n649), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n876), .B(new_n887), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n853), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n417), .A3(new_n851), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n865), .B1(new_n893), .B2(new_n847), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n874), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n368), .A2(new_n649), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n874), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n417), .A2(new_n845), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n891), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n885), .B(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n836), .B1(new_n879), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT110), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n904), .B2(new_n879), .ZN(new_n907));
  INV_X1    g0707(.A(new_n458), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n583), .B1(new_n908), .B2(KEYINPUT35), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n230), .A2(new_n207), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n909), .B(new_n910), .C1(KEYINPUT35), .C2(new_n908), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n383), .A2(G77), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n229), .A2(new_n913), .B1(G50), .B2(new_n212), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n642), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n907), .A2(new_n912), .A3(new_n915), .ZN(G367));
  NAND2_X1  g0716(.A1(new_n725), .A2(G1), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n463), .A2(new_n649), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n696), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n632), .A2(new_n649), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n667), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT45), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(KEYINPUT114), .B(KEYINPUT44), .Z(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n667), .ZN(new_n927));
  INV_X1    g0727(.A(new_n921), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n667), .A3(new_n925), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n663), .B1(new_n924), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n922), .B(KEYINPUT45), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n659), .A2(new_n662), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n930), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n662), .B1(new_n597), .B2(new_n649), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n665), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT115), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(KEYINPUT115), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n659), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(G330), .A3(new_n658), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n723), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n670), .B(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n917), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT43), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n615), .A2(new_n617), .A3(new_n650), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n614), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n680), .A2(new_n613), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n951), .B1(new_n952), .B2(new_n950), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT111), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n953), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n948), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n953), .A2(new_n954), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n569), .A2(new_n664), .A3(new_n696), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  INV_X1    g0762(.A(new_n696), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n464), .B1(new_n963), .B2(new_n566), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n650), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n958), .A2(new_n960), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n959), .A2(new_n955), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT42), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n961), .B(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n969), .A2(new_n971), .A3(new_n948), .A4(new_n965), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT112), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT112), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n663), .A2(new_n928), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(KEYINPUT113), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT113), .B1(new_n976), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n976), .A2(new_n977), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT113), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n984), .A2(KEYINPUT112), .A3(new_n973), .A4(new_n978), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n730), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n959), .B2(new_n955), .ZN(new_n988));
  INV_X1    g0788(.A(new_n779), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n777), .B1(new_n224), .B2(new_n319), .C1(new_n241), .C2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(G311), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n379), .B1(new_n738), .B2(new_n748), .C1(new_n744), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G97), .B2(new_n762), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n806), .A2(G107), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G283), .A2(new_n753), .B1(new_n760), .B2(new_n574), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n757), .A2(G116), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT46), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G317), .B2(new_n765), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n756), .A2(new_n227), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n765), .A2(G137), .B1(G143), .B2(new_n743), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n806), .A2(G68), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n761), .A2(new_n218), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G50), .B2(new_n753), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n287), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1000), .B(new_n1005), .C1(G150), .C2(new_n760), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n749), .A2(new_n766), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n999), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n829), .B(new_n990), .C1(new_n1009), .C2(new_n733), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n947), .A2(new_n986), .B1(new_n988), .B2(new_n1010), .ZN(G387));
  NAND2_X1  g0811(.A1(new_n806), .A2(new_n318), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n216), .B2(new_n759), .C1(new_n255), .C2(new_n748), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n756), .A2(new_n218), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n287), .B1(new_n761), .B2(new_n202), .C1(new_n212), .C2(new_n752), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n765), .B2(G150), .ZN(new_n1017));
  INV_X1    g0817(.A(G159), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1015), .B(new_n1017), .C1(new_n1018), .C2(new_n744), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1020), .A2(new_n759), .B1(new_n752), .B2(new_n573), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT119), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n743), .A2(G322), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n991), .C2(new_n748), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  INV_X1    g0825(.A(G283), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(new_n1026), .B2(new_n737), .C1(new_n738), .C2(new_n756), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT120), .Z(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n379), .B1(new_n583), .B2(new_n761), .C1(new_n745), .C2(new_n740), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1019), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n732), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n783), .A2(new_n672), .B1(new_n203), .B2(new_n669), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT116), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n316), .A2(new_n216), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT50), .Z(new_n1036));
  OR2_X1    g0836(.A1(new_n673), .A2(KEYINPUT117), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n673), .A2(KEYINPUT117), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1036), .A2(new_n508), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n212), .A2(new_n218), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n779), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT118), .Z(new_n1042));
  NOR2_X1   g0842(.A1(new_n238), .A2(new_n508), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1034), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n777), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1032), .A2(new_n829), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n662), .B2(new_n730), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n944), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1047), .B1(new_n917), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n944), .B1(new_n721), .B2(new_n722), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n670), .B1(new_n723), .B2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n723), .A2(new_n1048), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(KEYINPUT121), .A3(new_n936), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT121), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n932), .A2(new_n935), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1057), .A3(new_n670), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1056), .A2(new_n917), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n769), .B1(new_n573), .B2(new_n748), .C1(new_n737), .C2(new_n583), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n287), .B1(new_n765), .B2(G322), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n1026), .B2(new_n756), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT52), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n744), .A2(new_n1020), .B1(new_n991), .B2(new_n759), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1061), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n1064), .B2(new_n1065), .C1(new_n738), .C2(new_n752), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G150), .A2(new_n743), .B1(new_n760), .B2(G159), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT51), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n749), .A2(G50), .B1(new_n753), .B2(new_n316), .ZN(new_n1070));
  AND4_X1   g0870(.A1(new_n287), .A2(new_n1069), .A3(new_n812), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n757), .A2(G68), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n765), .A2(G143), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n806), .A2(G77), .B1(KEYINPUT51), .B2(new_n1068), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n733), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n246), .A2(new_n779), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n778), .B1(G97), .B2(new_n669), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1079), .B(new_n829), .C1(new_n987), .C2(new_n928), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1059), .A2(new_n1060), .A3(new_n1080), .ZN(G390));
  NAND2_X1  g0881(.A1(new_n897), .A2(new_n899), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n890), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n886), .B1(new_n794), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1084), .B2(new_n898), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n898), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n698), .A2(new_n650), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n890), .B1(new_n1087), .B2(new_n793), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n895), .C1(new_n1088), .C2(new_n886), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n720), .A2(new_n799), .A3(new_n887), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1085), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n422), .A2(G330), .A3(new_n802), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n880), .B(new_n421), .C1(new_n686), .C2(new_n700), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT108), .B1(new_n701), .B2(new_n422), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n612), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n887), .B1(new_n720), .B2(new_n799), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1088), .A2(new_n1090), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1090), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n889), .A2(new_n890), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1093), .A2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1091), .A2(new_n1092), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n670), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1082), .A2(new_n728), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n806), .A2(G77), .B1(G97), .B2(new_n753), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n583), .B2(new_n759), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n744), .A2(new_n1026), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n745), .A2(new_n738), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n287), .B1(new_n757), .B2(G87), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n212), .B2(new_n761), .C1(new_n203), .C2(new_n748), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n756), .A2(new_n259), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1118), .B1(new_n1018), .B2(new_n737), .C1(new_n745), .C2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(G128), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n744), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n761), .A2(new_n216), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI21_X1  g0924(.A(new_n379), .B1(new_n753), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G132), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n759), .C1(new_n815), .C2(new_n748), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n732), .B1(new_n1116), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1109), .A2(new_n829), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n255), .B2(new_n826), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1093), .B2(new_n917), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1108), .A2(new_n1132), .ZN(G378));
  NAND2_X1  g0933(.A1(new_n270), .A2(new_n845), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT123), .Z(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n606), .B2(new_n306), .ZN(new_n1139));
  AND4_X1   g0939(.A1(new_n303), .A2(new_n300), .A3(new_n306), .A4(new_n1138), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n307), .A2(new_n1137), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n606), .A2(new_n306), .A3(new_n1138), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1135), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n728), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1002), .B1(new_n227), .B2(new_n761), .C1(new_n202), .C2(new_n748), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n379), .B1(new_n319), .B2(new_n752), .C1(new_n744), .C2(new_n583), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1147), .A2(G41), .A3(new_n1014), .A4(new_n1148), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n203), .B2(new_n759), .C1(new_n1026), .C2(new_n745), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n216), .B1(new_n377), .B2(G41), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n759), .A2(new_n1121), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n744), .A2(new_n1119), .B1(new_n815), .B2(new_n752), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n757), .C2(new_n1124), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n1126), .B2(new_n748), .C1(new_n737), .C2(new_n259), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  INV_X1    g0958(.A(G33), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n762), .A2(new_n766), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G41), .B1(new_n765), .B2(G124), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1153), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n732), .B1(new_n1152), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n826), .A2(new_n216), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1146), .A2(new_n829), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1145), .B1(new_n877), .B2(new_n702), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT40), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n843), .B1(new_n703), .B2(new_n719), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n895), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n876), .A2(new_n1172), .A3(new_n1171), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1170), .B(G330), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n903), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n901), .B1(new_n1084), .B2(new_n876), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1178), .A2(new_n900), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT124), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n903), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT124), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1168), .B1(new_n1184), .B2(new_n917), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1097), .B1(new_n1093), .B2(new_n1105), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1176), .B(new_n903), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT57), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n670), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1097), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1101), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1085), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1190), .B1(new_n1194), .B2(new_n1104), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1184), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1185), .B1(new_n1189), .B2(new_n1196), .ZN(G375));
  NAND3_X1  g0997(.A1(new_n885), .A2(new_n1094), .A3(new_n1103), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1199), .A3(new_n946), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n744), .A2(new_n738), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n765), .A2(G303), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n379), .B1(new_n756), .B2(new_n202), .C1(new_n583), .C2(new_n748), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1003), .B(new_n1203), .C1(G107), .C2(new_n753), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n760), .A2(G283), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1012), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n765), .A2(G128), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n806), .A2(G50), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n760), .A2(G137), .B1(new_n749), .B2(new_n1124), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n752), .A2(new_n259), .B1(new_n761), .B2(new_n227), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n379), .B(new_n1210), .C1(G159), .C2(new_n757), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n744), .A2(new_n1126), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1201), .A2(new_n1206), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n732), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n829), .B(new_n1215), .C1(new_n887), .C2(new_n729), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n212), .B2(new_n826), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1103), .B2(new_n917), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1200), .A2(new_n1218), .ZN(G381));
  NOR2_X1   g1019(.A1(new_n1010), .A2(new_n988), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n917), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1056), .A2(new_n1048), .B1(new_n721), .B2(new_n722), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n946), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n981), .A2(new_n985), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1226), .A2(new_n1060), .A3(new_n1080), .A4(new_n1059), .ZN(new_n1227));
  OR3_X1    g1027(.A1(G375), .A2(new_n1227), .A3(G378), .ZN(new_n1228));
  INV_X1    g1028(.A(G396), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1049), .B(new_n1229), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G384), .A2(G381), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT125), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1232), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1228), .A2(new_n1234), .A3(new_n1235), .A4(new_n1230), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1233), .A2(new_n1236), .ZN(G407));
  INV_X1    g1037(.A(G375), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1108), .A2(new_n1132), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n648), .A3(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G213), .B(new_n1240), .C1(new_n1233), .C2(new_n1236), .ZN(G409));
  NAND3_X1  g1041(.A1(new_n1195), .A2(new_n1184), .A3(new_n946), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1187), .A2(new_n917), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1167), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1239), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1185), .C1(new_n1189), .C2(new_n1196), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n648), .A2(G213), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1097), .A2(new_n1104), .A3(KEYINPUT60), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1097), .A2(new_n1104), .A3(KEYINPUT126), .A4(KEYINPUT60), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1103), .B1(new_n885), .B2(new_n1094), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n670), .B(new_n1198), .C1(new_n1254), .C2(KEYINPUT60), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1218), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(G384), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n834), .B(new_n1218), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1247), .A2(new_n1248), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n648), .A2(G213), .A3(G2897), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1258), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n671), .B1(new_n1199), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(new_n1251), .A3(new_n1198), .A4(new_n1252), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n834), .B1(new_n1268), .B2(new_n1218), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1264), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1257), .A2(new_n1258), .A3(new_n1263), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1262), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1247), .A2(new_n1275), .A3(new_n1248), .A4(new_n1259), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1261), .A2(new_n1273), .A3(new_n1274), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G390), .A2(G387), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1230), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1227), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1227), .B2(new_n1278), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1277), .A2(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1248), .A2(new_n1247), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1260), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1248), .A4(new_n1259), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1289), .A2(new_n1283), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1274), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1285), .A2(new_n1291), .ZN(G405));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1238), .A2(G378), .B1(new_n1259), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1239), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1227), .A2(new_n1278), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1280), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1227), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1298), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1298), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1296), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1283), .A2(new_n1298), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1297), .B(KEYINPUT127), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1306), .A2(new_n1307), .B1(new_n1295), .B2(new_n1294), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1305), .A2(new_n1308), .ZN(G402));
endmodule


