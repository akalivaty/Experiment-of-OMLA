//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT26), .B(G101), .Z(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT73), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n197), .B1(new_n202), .B2(new_n196), .ZN(new_n203));
  AOI21_X1  g017(.A(G137), .B1(new_n199), .B2(new_n201), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(new_n204), .B2(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(G134), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(G137), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n203), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT68), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n210), .B2(KEYINPUT67), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n214));
  AOI211_X1 g028(.A(new_n214), .B(new_n203), .C1(new_n205), .C2(new_n209), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n212), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n203), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n200), .A2(G134), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n196), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n206), .B1(new_n220), .B2(new_n207), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n204), .A2(KEYINPUT66), .A3(KEYINPUT11), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n214), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(KEYINPUT68), .A3(G131), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G143), .B(G146), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n232), .B(new_n233), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n229), .A2(G146), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n227), .A2(G143), .ZN(new_n241));
  OAI22_X1  g055(.A1(new_n240), .A2(new_n241), .B1(new_n234), .B2(new_n235), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n233), .B1(new_n242), .B2(new_n232), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n216), .A2(new_n226), .A3(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n211), .B(new_n217), .C1(new_n221), .C2(new_n222), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n228), .A2(new_n230), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n247), .A2(new_n248), .B1(KEYINPUT1), .B2(new_n241), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n237), .A2(KEYINPUT69), .A3(new_n251), .A4(G128), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n204), .B1(new_n198), .B2(G137), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n246), .B(new_n255), .C1(new_n211), .C2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n245), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n242), .A2(new_n232), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n216), .A2(new_n226), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n262), .B2(new_n257), .ZN(new_n263));
  INV_X1    g077(.A(G116), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G119), .ZN(new_n265));
  INV_X1    g079(.A(G119), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n266), .B2(G116), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n264), .A3(G119), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n265), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT2), .B(G113), .Z(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n258), .A2(new_n263), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n245), .A2(new_n273), .A3(new_n257), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n195), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(KEYINPUT28), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n245), .A2(new_n280), .A3(new_n273), .A4(new_n257), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n262), .A2(new_n257), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n272), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n284), .A3(new_n194), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n277), .A2(new_n278), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n273), .B1(new_n245), .B2(new_n257), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n279), .B2(new_n281), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n187), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n194), .B1(new_n282), .B2(new_n284), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n275), .A2(new_n194), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n274), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n283), .A2(new_n259), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n245), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n272), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n295), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(KEYINPUT31), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n293), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G472), .A2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT32), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n282), .A2(new_n284), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n195), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n299), .A2(KEYINPUT31), .A3(new_n300), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT31), .B1(new_n299), .B2(new_n300), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n303), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n292), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n315));
  AOI21_X1  g129(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n316));
  OAI21_X1  g130(.A(G131), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n190), .A2(G214), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n229), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n211), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT17), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n227), .ZN(new_n332));
  OAI211_X1 g146(.A(G146), .B(new_n326), .C1(new_n330), .C2(new_n324), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT17), .B(G131), .C1(new_n315), .C2(new_n316), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n323), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(KEYINPUT18), .B(G131), .C1(new_n315), .C2(new_n316), .ZN(new_n337));
  NAND2_X1  g151(.A1(KEYINPUT18), .A2(G131), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n319), .A2(new_n320), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n330), .A2(G146), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n329), .A3(new_n227), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT87), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n314), .B1(new_n336), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G113), .B(G122), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n346), .ZN(new_n353));
  INV_X1    g167(.A(new_n340), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n335), .A3(KEYINPUT90), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n348), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n351), .B(KEYINPUT89), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n355), .A3(new_n335), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G475), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n330), .B1(KEYINPUT88), .B2(KEYINPUT19), .ZN(new_n363));
  AND2_X1   g177(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n327), .B(new_n329), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n333), .B1(new_n367), .B2(G146), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n317), .A2(new_n321), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n352), .B1(new_n370), .B2(new_n347), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n359), .ZN(new_n372));
  NOR2_X1   g186(.A1(G475), .A2(G902), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n362), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  AOI211_X1 g189(.A(KEYINPUT20), .B(new_n375), .C1(new_n371), .C2(new_n359), .ZN(new_n376));
  OAI22_X1  g190(.A1(new_n360), .A2(new_n361), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n229), .A2(G128), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n248), .A2(G143), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n208), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n202), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g197(.A1(KEYINPUT91), .A2(G122), .ZN(new_n384));
  NOR2_X1   g198(.A1(KEYINPUT91), .A2(G122), .ZN(new_n385));
  OAI21_X1  g199(.A(G116), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n264), .A2(G122), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(KEYINPUT14), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n264), .A3(G122), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n386), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n383), .B(new_n389), .C1(new_n393), .C2(new_n387), .ZN(new_n394));
  INV_X1    g208(.A(new_n389), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n387), .B1(new_n386), .B2(new_n388), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n380), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT13), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n379), .B1(new_n378), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT92), .B1(new_n378), .B2(new_n398), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n378), .A2(KEYINPUT92), .A3(new_n398), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n198), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n394), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT77), .ZN(new_n406));
  INV_X1    g220(.A(G217), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(G953), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n408), .B(new_n394), .C1(new_n403), .C2(new_n397), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(KEYINPUT93), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G902), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT93), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n404), .A2(new_n414), .A3(new_n409), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G478), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT15), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n418), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n412), .A2(new_n413), .A3(new_n415), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(G234), .A2(G237), .ZN(new_n423));
  INV_X1    g237(.A(G953), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(G952), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(G902), .A3(G953), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(G898), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n377), .A2(new_n422), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G214), .B1(G237), .B2(G902), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G122), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT3), .B1(new_n350), .B2(G107), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT78), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n387), .A2(G104), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT78), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT3), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT3), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n387), .A3(G104), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n350), .A2(G107), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n439), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G101), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n441), .A2(new_n442), .ZN(new_n445));
  INV_X1    g259(.A(G101), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n439), .A4(new_n436), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(KEYINPUT4), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n443), .A2(new_n449), .A3(G101), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n272), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n451), .A2(KEYINPUT84), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n448), .A2(new_n453), .A3(new_n272), .A4(new_n450), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT79), .B1(new_n350), .B2(G107), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n387), .A2(G104), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G101), .B1(new_n437), .B2(KEYINPUT79), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n437), .A2(new_n442), .A3(KEYINPUT79), .ZN(new_n461));
  OR3_X1    g275(.A1(new_n350), .A2(KEYINPUT79), .A3(G107), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT80), .A4(G101), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n266), .A2(G116), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(G113), .C1(KEYINPUT5), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n270), .A2(new_n271), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n447), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n454), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n434), .B1(new_n452), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n451), .A2(KEYINPUT84), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n472), .A2(new_n433), .A3(new_n469), .A4(new_n454), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(new_n434), .C1(new_n452), .C2(new_n470), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n328), .B1(new_n242), .B2(new_n232), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n255), .B2(new_n328), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n424), .A2(G224), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n478), .B(new_n479), .Z(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(KEYINPUT86), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(KEYINPUT7), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n468), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n447), .A2(new_n463), .A3(new_n460), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n469), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n433), .B(new_n491), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n485), .A2(new_n486), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n493), .B2(new_n473), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n481), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n481), .B2(new_n494), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n431), .B(new_n432), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G221), .B1(new_n406), .B2(G902), .ZN(new_n500));
  XNOR2_X1  g314(.A(G110), .B(G140), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n424), .A2(G227), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n488), .B(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n507));
  AND4_X1   g321(.A1(new_n216), .A2(new_n226), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n448), .A2(new_n244), .A3(new_n450), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT10), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n488), .B2(new_n505), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n464), .A2(KEYINPUT10), .A3(new_n255), .A4(new_n447), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n216), .B2(new_n226), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n216), .A2(new_n226), .A3(new_n506), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n504), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n509), .A2(new_n512), .A3(new_n511), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n246), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n211), .B1(new_n223), .B2(new_n214), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n523), .B2(new_n225), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n213), .A2(new_n521), .A3(new_n215), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT82), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n513), .A2(new_n216), .A3(new_n226), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n513), .A2(new_n216), .A3(new_n226), .A4(KEYINPUT82), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n503), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n413), .B1(new_n519), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n533), .A3(G469), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n503), .A3(new_n530), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n216), .A2(new_n226), .A3(new_n506), .A4(new_n507), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n518), .A2(new_n536), .A3(new_n526), .A4(new_n504), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G469), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n533), .B1(new_n532), .B2(G469), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n499), .B(new_n500), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G234), .ZN(new_n544));
  OAI21_X1  g358(.A(G217), .B1(new_n544), .B2(G902), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n266), .A2(G128), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT76), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n248), .A2(G119), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT75), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT24), .B(G110), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n266), .B2(G128), .ZN(new_n556));
  INV_X1    g370(.A(new_n549), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n558), .A2(G110), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n333), .B(new_n342), .C1(new_n553), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n332), .A2(new_n333), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(G110), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n562), .B(new_n563), .C1(new_n552), .C2(new_n551), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT22), .B(G137), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n424), .A2(G221), .A3(G234), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n565), .B(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n569), .A2(KEYINPUT25), .A3(new_n413), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT25), .B1(new_n569), .B2(new_n413), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n546), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n544), .B2(G217), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n313), .A2(new_n543), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT94), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G3));
  INV_X1    g392(.A(new_n500), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n534), .A2(new_n540), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n529), .A2(new_n530), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n504), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n518), .A2(new_n536), .A3(new_n526), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n503), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT83), .B1(new_n585), .B2(new_n539), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n579), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n575), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n310), .A2(new_n413), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n589), .A2(G472), .B1(new_n303), .B2(new_n310), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT95), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n481), .A2(new_n494), .ZN(new_n593));
  INV_X1    g407(.A(new_n495), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n481), .A2(new_n494), .A3(new_n495), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n432), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n497), .B2(KEYINPUT96), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n377), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n412), .A2(new_n603), .A3(new_n415), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n410), .A2(KEYINPUT33), .A3(new_n411), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(G478), .A3(new_n413), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n416), .A2(new_n417), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n606), .A2(KEYINPUT97), .A3(new_n607), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n602), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n430), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n592), .A2(new_n601), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n422), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n377), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n430), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n592), .A2(new_n601), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT99), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT98), .B(KEYINPUT35), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  XNOR2_X1  g441(.A(new_n565), .B(KEYINPUT100), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n568), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n628), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n573), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n632), .A2(new_n572), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n587), .A2(new_n590), .A3(new_n499), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  NAND2_X1  g451(.A1(new_n305), .A2(new_n312), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n286), .A2(new_n291), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n633), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n586), .A2(new_n534), .A3(new_n540), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT101), .B(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n426), .B1(new_n643), .B2(new_n428), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n621), .A2(new_n644), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n500), .A2(new_n642), .A3(new_n601), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  XOR2_X1   g462(.A(new_n644), .B(KEYINPUT39), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n587), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n602), .A2(new_n619), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n633), .A2(new_n432), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n496), .A2(new_n497), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n587), .A2(new_n661), .A3(new_n649), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n195), .B1(new_n276), .B2(new_n287), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n299), .A2(new_n300), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n668), .B2(G902), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n638), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n651), .A2(new_n660), .A3(new_n662), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G143), .ZN(G45));
  AND3_X1   g486(.A1(new_n642), .A2(new_n500), .A3(new_n601), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n302), .A2(KEYINPUT32), .A3(new_n304), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n311), .B1(new_n310), .B2(new_n303), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n640), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n644), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n612), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n676), .A3(new_n634), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NOR2_X1   g495(.A1(new_n539), .A2(KEYINPUT105), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n538), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n538), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n500), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n598), .A2(new_n600), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n676), .A2(new_n588), .A3(new_n615), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND4_X1  g505(.A1(new_n676), .A2(new_n588), .A3(new_n622), .A4(new_n688), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NOR2_X1   g507(.A1(new_n538), .A2(new_n683), .ZN(new_n694));
  AOI211_X1 g508(.A(G902), .B(new_n682), .C1(new_n535), .C2(new_n537), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n694), .A2(new_n695), .A3(new_n579), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n601), .A2(KEYINPUT106), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n686), .B2(new_n687), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n431), .A3(new_n641), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NAND3_X1  g516(.A1(new_n598), .A2(new_n600), .A3(new_n652), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n686), .A2(new_n703), .A3(new_n430), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n187), .B1(new_n310), .B2(new_n413), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n296), .A2(new_n301), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n288), .A2(new_n194), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n304), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n704), .A2(new_n709), .A3(new_n588), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT107), .B(G122), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G24));
  NOR3_X1   g526(.A1(new_n705), .A2(new_n633), .A3(new_n708), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n679), .A3(new_n699), .A4(new_n697), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  NAND3_X1  g529(.A1(new_n657), .A2(new_n500), .A3(new_n432), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n519), .B1(new_n717), .B2(new_n531), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n582), .A2(KEYINPUT108), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(G469), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n539), .A2(new_n413), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n538), .B2(new_n539), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n716), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n676), .A2(new_n588), .A3(new_n679), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n575), .B1(new_n638), .B2(new_n640), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(KEYINPUT42), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(new_n679), .A3(new_n723), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NAND4_X1  g548(.A1(new_n676), .A2(new_n588), .A3(new_n645), .A4(new_n723), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NAND2_X1  g550(.A1(new_n657), .A2(new_n432), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n590), .A2(new_n633), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n377), .B(KEYINPUT110), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n610), .A2(new_n611), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n377), .A2(KEYINPUT43), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n743), .A2(KEYINPUT111), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT111), .B1(new_n743), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n738), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n737), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n718), .A2(KEYINPUT45), .A3(new_n719), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n582), .A2(new_n584), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n539), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n721), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n540), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n500), .B(new_n649), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n751), .B(new_n760), .C1(new_n750), .C2(new_n749), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  OAI21_X1  g576(.A(new_n500), .B1(new_n757), .B2(new_n758), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n765), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n676), .A2(new_n588), .A3(new_n678), .A4(new_n737), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NOR3_X1   g584(.A1(new_n742), .A2(new_n425), .A3(new_n745), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n686), .A2(new_n737), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n728), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT48), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n709), .A2(new_n771), .A3(new_n588), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n697), .A2(new_n699), .ZN(new_n780));
  OAI211_X1 g594(.A(G952), .B(new_n424), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n772), .A2(new_n588), .A3(new_n426), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n670), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n781), .B1(new_n612), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n777), .A2(KEYINPUT48), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n778), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n766), .A2(new_n767), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n694), .A2(new_n695), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n500), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n779), .A2(new_n737), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT51), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n741), .A2(new_n377), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n775), .A2(new_n713), .B1(new_n783), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n659), .A2(new_n599), .A3(new_n696), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n779), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT50), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n797), .A2(KEYINPUT50), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n786), .B1(new_n793), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n804), .A2(new_n792), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n806), .B2(KEYINPUT51), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n377), .A2(new_n422), .A3(new_n644), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n432), .A2(new_n808), .A3(new_n595), .A4(new_n597), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n500), .B(new_n809), .C1(new_n541), .C2(new_n542), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n676), .A3(new_n634), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n713), .A2(new_n679), .A3(new_n723), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n735), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n720), .A2(new_n722), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n633), .A2(new_n500), .A3(new_n677), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n816), .A2(new_n817), .A3(new_n703), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n670), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n647), .A2(new_n680), .A3(new_n714), .A4(new_n819), .ZN(new_n820));
  AOI221_X4 g634(.A(new_n814), .B1(new_n727), .B2(new_n732), .C1(new_n820), .C2(KEYINPUT52), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n589), .A2(G472), .ZN(new_n823));
  INV_X1    g637(.A(new_n708), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n588), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n601), .A2(new_n613), .A3(new_n696), .A4(new_n652), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n310), .A2(new_n303), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n302), .A2(G902), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n827), .B(new_n634), .C1(new_n828), .C2(new_n187), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n825), .A2(new_n826), .B1(new_n829), .B2(new_n543), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n576), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n612), .A2(new_n620), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n432), .B1(new_n496), .B2(new_n497), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n832), .A2(new_n833), .A3(new_n430), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n587), .A2(new_n590), .A3(new_n834), .A4(new_n588), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n728), .B(new_n688), .C1(new_n615), .C2(new_n622), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n831), .A2(new_n701), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n822), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n821), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n814), .B1(new_n727), .B2(new_n732), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n676), .A2(new_n431), .A3(new_n634), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n689), .B(new_n692), .C1(new_n841), .C2(new_n780), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n676), .A2(new_n588), .A3(new_n587), .A4(new_n499), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n635), .A3(new_n835), .A4(new_n710), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n705), .A2(new_n708), .A3(new_n633), .A4(new_n678), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n700), .A2(new_n847), .B1(new_n641), .B2(new_n646), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n680), .A4(new_n819), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n840), .A2(new_n845), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(new_n849), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(KEYINPUT53), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT54), .B1(new_n839), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n821), .A2(new_n838), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n851), .A2(new_n856), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n807), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(G952), .A2(G953), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n740), .A2(new_n741), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n588), .A2(new_n500), .A3(new_n432), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n788), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n659), .A3(new_n869), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n863), .A2(new_n864), .B1(new_n670), .B2(new_n870), .ZN(G75));
  NOR2_X1   g685(.A1(new_n424), .A2(G952), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT116), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n474), .A2(new_n476), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n480), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT55), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n858), .A2(new_n859), .ZN(new_n877));
  NAND2_X1  g691(.A1(G210), .A2(G902), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n858), .B2(new_n859), .ZN(new_n883));
  INV_X1    g697(.A(new_n876), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n873), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT117), .B(new_n873), .C1(new_n882), .C2(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(G51));
  XNOR2_X1  g704(.A(new_n721), .B(KEYINPUT57), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n860), .B1(new_n858), .B2(new_n859), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n535), .A2(new_n537), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n852), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT53), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n851), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n839), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n413), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n752), .A3(new_n755), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n872), .B1(new_n896), .B2(new_n902), .ZN(G54));
  NAND2_X1  g717(.A1(KEYINPUT58), .A2(G475), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT118), .Z(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n372), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n372), .B1(new_n901), .B2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n872), .ZN(G60));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n909));
  XOR2_X1   g723(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n910));
  NOR2_X1   g724(.A1(new_n417), .A2(new_n413), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n862), .A2(new_n912), .B1(new_n604), .B2(new_n605), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n604), .A2(new_n605), .A3(new_n912), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n892), .B2(new_n893), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n873), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n909), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n897), .A2(new_n856), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n821), .A2(new_n838), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n860), .B1(new_n919), .B2(new_n859), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n912), .B1(new_n892), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n604), .A2(new_n605), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(KEYINPUT120), .A3(new_n873), .A4(new_n915), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n924), .ZN(G63));
  INV_X1    g739(.A(new_n569), .ZN(new_n926));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n900), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n928), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n631), .B(KEYINPUT121), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n877), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n873), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G66));
  INV_X1    g749(.A(G224), .ZN(new_n936));
  OAI21_X1  g750(.A(G953), .B1(new_n429), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n845), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n874), .B1(G898), .B2(new_n424), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT122), .Z(new_n940));
  XNOR2_X1  g754(.A(new_n938), .B(new_n940), .ZN(G69));
  AND2_X1   g755(.A1(new_n761), .A2(new_n769), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n943));
  INV_X1    g757(.A(new_n728), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n703), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n760), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n647), .A2(new_n680), .A3(new_n714), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n946), .A2(new_n947), .A3(new_n735), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n942), .A2(new_n943), .A3(new_n733), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n761), .A2(new_n769), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n946), .A2(new_n947), .A3(new_n733), .A4(new_n735), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT123), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n424), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n258), .A2(new_n263), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n367), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n947), .A2(new_n671), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n761), .A3(new_n769), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n650), .A2(new_n737), .A3(new_n832), .ZN(new_n961));
  OAI22_X1  g775(.A1(new_n958), .A2(KEYINPUT62), .B1(new_n944), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n424), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n424), .B1(G227), .B2(G900), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n963), .A2(new_n955), .B1(KEYINPUT124), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n957), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G72));
  XNOR2_X1  g782(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n187), .A2(new_n413), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n277), .B2(new_n666), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n839), .B2(new_n854), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n960), .A2(new_n837), .A3(new_n962), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n274), .A2(new_n276), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n978), .A2(new_n195), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n976), .A2(new_n975), .A3(new_n972), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n974), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n872), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n949), .A2(new_n845), .A3(new_n952), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n984), .A2(new_n971), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n978), .A2(new_n195), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT127), .B(new_n983), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n984), .B2(new_n971), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n872), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n982), .B1(new_n987), .B2(new_n990), .ZN(G57));
endmodule


