//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n446, new_n451, new_n454,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(G217));
  NAND4_X1  g030(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT2), .ZN(new_n458));
  NOR4_X1   g033(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  AOI22_X1  g037(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g048(.A(KEYINPUT67), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(new_n468), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(G124), .A3(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n472), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n483), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n477), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(KEYINPUT68), .A3(new_n483), .A4(new_n485), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n490), .A2(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(new_n472), .B2(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n497), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT70), .B(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n482), .A2(new_n504), .A3(G138), .A4(new_n472), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n472), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n482), .A2(G126), .A3(G2105), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n503), .A2(new_n505), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(G651), .ZN(new_n518));
  NOR3_X1   g093(.A1(new_n514), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n513), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT71), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n516), .A2(new_n517), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(KEYINPUT72), .A3(new_n515), .A4(new_n513), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n522), .A2(G88), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n525), .A2(G543), .A3(new_n515), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G62), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n530), .A2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND3_X1  g117(.A1(new_n522), .A2(G89), .A3(new_n526), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT74), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n528), .A2(G51), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n543), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  NAND3_X1  g125(.A1(new_n522), .A2(G90), .A3(new_n526), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n514), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n528), .A2(G52), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT75), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n551), .A2(new_n557), .A3(new_n553), .A4(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(G171));
  AOI22_X1  g134(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n514), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n528), .A2(G43), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n522), .A2(new_n526), .ZN(new_n563));
  INV_X1    g138(.A(G81), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT76), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  XNOR2_X1  g145(.A(KEYINPUT77), .B(KEYINPUT8), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n572), .B(new_n573), .Z(new_n574));
  NAND2_X1  g149(.A1(new_n569), .A2(new_n574), .ZN(G188));
  NAND3_X1  g150(.A1(new_n522), .A2(G91), .A3(new_n526), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n525), .A2(G53), .A3(G543), .A4(new_n515), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n528), .A2(KEYINPUT9), .A3(G53), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n514), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n576), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  OAI21_X1  g159(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n528), .A2(G49), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n563), .C2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n536), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n528), .A2(G48), .B1(G651), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n563), .B2(new_n593), .ZN(G305));
  INV_X1    g169(.A(new_n563), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G85), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n514), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n528), .A2(G47), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n522), .A2(G92), .A3(new_n526), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT79), .B(G66), .Z(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n536), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n528), .A2(G54), .B1(new_n606), .B2(G651), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n522), .A2(new_n608), .A3(G92), .A4(new_n526), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n603), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT80), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(G860), .B2(new_n618), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g198(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n477), .A2(new_n472), .ZN(new_n629));
  AOI22_X1  g204(.A1(G123), .A2(new_n629), .B1(new_n491), .B2(G135), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G111), .C2(new_n472), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n628), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2435), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2438), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  NOR2_X1   g229(.A1(G2072), .A2(G2078), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n445), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n656), .B(KEYINPUT86), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n661), .B(new_n663), .C1(new_n665), .C2(new_n659), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n659), .A3(new_n662), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n657), .A2(new_n659), .A3(new_n663), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n637), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n627), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n680), .A3(new_n682), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(new_n684), .C2(new_n683), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT22), .B(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G4), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n611), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G1348), .ZN(new_n697));
  NOR2_X1   g272(.A1(G27), .A2(G29), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G164), .B2(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G2078), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G33), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n491), .A2(G139), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n704), .B(new_n705), .C1(new_n472), .C2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n702), .B1(new_n708), .B2(new_n701), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G2072), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n443), .B(new_n702), .C1(new_n708), .C2(new_n701), .ZN(new_n711));
  OR2_X1    g286(.A1(G16), .A2(G19), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n565), .B2(new_n694), .ZN(new_n713));
  INV_X1    g288(.A(G1341), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n701), .A2(G35), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n716), .B(new_n717), .C1(G162), .C2(new_n701), .ZN(new_n718));
  INV_X1    g293(.A(G2090), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n701), .B1(new_n490), .B2(new_n493), .ZN(new_n720));
  INV_X1    g295(.A(new_n717), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT29), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n718), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n713), .A2(new_n714), .ZN(new_n724));
  AND4_X1   g299(.A1(new_n711), .A2(new_n715), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n697), .A2(new_n700), .A3(new_n710), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n701), .A2(G26), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n629), .A2(G128), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n491), .A2(G140), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(new_n701), .ZN(new_n734));
  MUX2_X1   g309(.A(new_n727), .B(new_n734), .S(KEYINPUT28), .Z(new_n735));
  XOR2_X1   g310(.A(KEYINPUT91), .B(G2067), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n738), .A2(new_n701), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G160), .B2(new_n701), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2084), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n699), .A2(G2078), .ZN(new_n743));
  NOR4_X1   g318(.A1(new_n726), .A2(new_n737), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(KEYINPUT23), .B1(new_n694), .B2(G20), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n694), .A2(KEYINPUT23), .A3(G20), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT99), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT99), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n746), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1956), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n718), .A2(new_n722), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2090), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n749), .A2(G1956), .A3(new_n751), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT100), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n491), .A2(G141), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n629), .A2(G129), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT26), .Z(new_n766));
  NAND4_X1  g341(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT93), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  OR2_X1    g344(.A1(G29), .A2(G32), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n761), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n761), .B2(new_n769), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n744), .A2(new_n760), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n696), .A2(G1348), .ZN(new_n776));
  NOR2_X1   g351(.A1(G5), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G171), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT96), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(KEYINPUT96), .B(new_n777), .C1(G171), .C2(G16), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n780), .A2(new_n781), .A3(G1961), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n775), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT36), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  NAND2_X1  g360(.A1(G303), .A2(G16), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n694), .A2(G22), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n787), .ZN(new_n789));
  AOI211_X1 g364(.A(G1971), .B(new_n789), .C1(G303), .C2(G16), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n694), .A2(G23), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G288), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT33), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n796), .A2(G1976), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n694), .A2(G6), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n591), .A2(G651), .ZN(new_n800));
  INV_X1    g375(.A(G48), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n525), .A2(G543), .A3(new_n515), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n595), .B2(G86), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n799), .B1(new_n804), .B2(new_n694), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G1976), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n793), .A2(new_n794), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n795), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n791), .A2(new_n798), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n694), .A2(G24), .ZN(new_n813));
  INV_X1    g388(.A(G290), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n694), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(G1986), .Z(new_n816));
  INV_X1    g391(.A(KEYINPUT87), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n491), .A2(new_n817), .A3(G131), .ZN(new_n818));
  INV_X1    g393(.A(G131), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT87), .B1(new_n486), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n629), .A2(G119), .ZN(new_n821));
  OR3_X1    g396(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n472), .A2(G107), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n822), .A2(new_n823), .A3(G2104), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n818), .A2(new_n820), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT89), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G25), .B(new_n830), .S(G29), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n812), .A2(KEYINPUT90), .A3(new_n816), .A4(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n816), .B(new_n834), .C1(new_n811), .C2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT90), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n784), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n840), .ZN(new_n842));
  AOI211_X1 g417(.A(KEYINPUT36), .B(new_n842), .C1(new_n835), .C2(new_n838), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n783), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT30), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(G28), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(G28), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n846), .A2(new_n847), .A3(G29), .ZN(new_n848));
  OAI21_X1  g423(.A(G1961), .B1(new_n780), .B2(new_n781), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(KEYINPUT97), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(KEYINPUT97), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(G16), .A2(G21), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G168), .B2(G16), .ZN(new_n854));
  INV_X1    g429(.A(G1966), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n630), .A2(G29), .A3(new_n635), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT31), .B(G11), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT95), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n852), .A2(new_n856), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT98), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n844), .A2(new_n861), .ZN(G311));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n860), .B(new_n863), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(new_n783), .C1(new_n841), .C2(new_n843), .ZN(G150));
  XNOR2_X1  g440(.A(KEYINPUT101), .B(G93), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n522), .A2(new_n526), .A3(new_n866), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(new_n514), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n528), .A2(G55), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n565), .B(new_n871), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n611), .A2(G559), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n874), .B1(new_n879), .B2(G860), .ZN(G145));
  XNOR2_X1  g455(.A(G160), .B(new_n636), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n472), .A2(G118), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT104), .Z(new_n885));
  OAI211_X1 g460(.A(new_n885), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n491), .A2(G142), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n629), .A2(G130), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n828), .A2(new_n829), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n828), .B2(new_n829), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT105), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n830), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n828), .A2(new_n829), .A3(new_n889), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n892), .A2(new_n897), .A3(new_n625), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n625), .B1(new_n892), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n883), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n768), .A2(KEYINPUT103), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n768), .A2(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G164), .B(new_n732), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n906), .A3(new_n902), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n907), .A3(new_n708), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n904), .B(new_n767), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n707), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n625), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT105), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n892), .A2(new_n897), .A3(new_n625), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT106), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n900), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n911), .B1(new_n900), .B2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n882), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n900), .A2(new_n917), .ZN(new_n923));
  INV_X1    g498(.A(new_n911), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n882), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n911), .A2(new_n916), .A3(new_n915), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n921), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g505(.A1(G299), .A2(KEYINPUT107), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n577), .B(KEYINPUT9), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n932), .A2(new_n933), .A3(new_n576), .A4(new_n582), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n931), .A2(new_n610), .A3(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n610), .A2(KEYINPUT107), .A3(G299), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT41), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n603), .A2(new_n609), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n938), .A2(new_n615), .A3(new_n933), .A4(new_n607), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n931), .A2(new_n610), .A3(new_n934), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(KEYINPUT109), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n935), .A2(new_n936), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n945), .A3(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n944), .A2(KEYINPUT108), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n620), .B(new_n875), .ZN(new_n951));
  MUX2_X1   g526(.A(new_n947), .B(new_n950), .S(new_n951), .Z(new_n952));
  INV_X1    g527(.A(G288), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G305), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n804), .A2(G288), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(G290), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G290), .B1(new_n954), .B2(new_n955), .ZN(new_n958));
  OAI21_X1  g533(.A(G303), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n958), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(G166), .A3(new_n956), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT42), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n952), .A2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n871), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(G868), .B2(new_n967), .ZN(G295));
  OAI21_X1  g543(.A(new_n966), .B1(G868), .B2(new_n967), .ZN(G331));
  NAND2_X1  g544(.A1(new_n566), .A2(new_n871), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n565), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n556), .A2(G286), .A3(new_n558), .ZN(new_n973));
  AOI21_X1  g548(.A(G286), .B1(new_n556), .B2(new_n558), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G171), .A2(G168), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n556), .A2(G286), .A3(new_n558), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n875), .A3(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(new_n943), .A3(new_n946), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n978), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n944), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n962), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n922), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n962), .B1(new_n980), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n937), .A2(new_n942), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n948), .A2(new_n949), .A3(new_n981), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n979), .A2(KEYINPUT111), .A3(new_n988), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n962), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n922), .A4(new_n983), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(KEYINPUT43), .C1(new_n984), .C2(new_n985), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n997), .B1(new_n984), .B2(new_n985), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n996), .A2(new_n922), .A3(new_n983), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n997), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT44), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1007), .ZN(G397));
  XOR2_X1   g583(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n511), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n482), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT67), .B1(new_n1013), .B2(G2105), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n471), .A2(new_n464), .A3(new_n472), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(G40), .A4(new_n480), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1996), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1020), .A2(new_n768), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1021), .A2(KEYINPUT113), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(KEYINPUT113), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1017), .ZN(new_n1024));
  INV_X1    g599(.A(G2067), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n732), .B(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n767), .A2(G1996), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1022), .A2(new_n1023), .A3(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n830), .B(new_n833), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(G290), .B(G1986), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1017), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1016), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n511), .A2(new_n1010), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1035), .B(KEYINPUT118), .C1(new_n1037), .C2(KEYINPUT45), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1009), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n511), .B2(new_n1010), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1016), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G2078), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1012), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1016), .B1(new_n1011), .B2(KEYINPUT114), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1037), .A2(KEYINPUT45), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n444), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1961), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n511), .B2(new_n1010), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n1016), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n511), .A2(new_n1054), .A3(new_n1010), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1052), .A2(new_n1044), .B1(new_n1053), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1047), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G301), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT126), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n479), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT124), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(G2105), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1014), .A2(new_n1015), .A3(G40), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1064), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n475), .A2(KEYINPUT125), .A3(new_n1068), .A4(G40), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1051), .A2(new_n1012), .A3(new_n1045), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT45), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1036), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1077), .A2(new_n1011), .A3(new_n1046), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT126), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1060), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1034), .B1(new_n1062), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1077), .B1(new_n1048), .B2(new_n1012), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1050), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1059), .A2(new_n753), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(KEYINPUT57), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n576), .A2(new_n582), .ZN(new_n1092));
  OR2_X1    g667(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n932), .B2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n932), .A2(KEYINPUT120), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(G299), .A2(new_n1090), .A3(KEYINPUT57), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1016), .A2(new_n1036), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1059), .A2(new_n1100), .B1(new_n1025), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n610), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1087), .A2(new_n1088), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1085), .A2(new_n1018), .A3(new_n1050), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1016), .B2(new_n1036), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n565), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1109), .B(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1101), .A2(new_n1025), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1057), .A2(new_n1055), .A3(new_n1016), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT60), .B(new_n1113), .C1(new_n1114), .C2(G1348), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(KEYINPUT122), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(KEYINPUT122), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(new_n607), .A3(new_n938), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(KEYINPUT122), .A3(new_n610), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1112), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1105), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1981), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n804), .A2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT116), .B(G86), .Z(new_n1131));
  NAND3_X1  g706(.A1(new_n522), .A2(new_n526), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n592), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1130), .A2(KEYINPUT49), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT49), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G305), .A2(G1981), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n1133), .ZN(new_n1138));
  INV_X1    g713(.A(G8), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1101), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1140), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G288), .A2(new_n808), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT52), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT52), .B1(G288), .B2(new_n808), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1140), .B(new_n1145), .C1(new_n808), .C2(G288), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1141), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT55), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(G303), .B2(G8), .ZN(new_n1149));
  AOI211_X1 g724(.A(KEYINPUT55), .B(new_n1139), .C1(new_n530), .C2(new_n540), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT115), .B(G1971), .Z(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1085), .B2(new_n1050), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1059), .A2(G2090), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1151), .B(G8), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1153), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1059), .A2(KEYINPUT117), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1114), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1159), .A3(new_n719), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1139), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1147), .B(new_n1155), .C1(new_n1161), .C2(new_n1151), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1163), .B1(new_n1082), .B2(G171), .ZN(new_n1164));
  AOI211_X1 g739(.A(KEYINPUT127), .B(G301), .C1(new_n1081), .C2(new_n1060), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1034), .B1(new_n1061), .B2(G301), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1162), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(G286), .A2(G8), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT123), .Z(new_n1170));
  INV_X1    g745(.A(G2084), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1043), .A2(new_n855), .B1(new_n1171), .B2(new_n1114), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1172), .B2(new_n1139), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT51), .B1(new_n1172), .B2(new_n1170), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(KEYINPUT51), .B(new_n1170), .C1(new_n1172), .C2(new_n1139), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AND4_X1   g752(.A1(new_n1084), .A2(new_n1128), .A3(new_n1168), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(KEYINPUT62), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1162), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1175), .A2(new_n1181), .A3(new_n1176), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1179), .A2(new_n1180), .A3(new_n1062), .A4(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1141), .A2(new_n808), .A3(new_n953), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1142), .B1(new_n1184), .B2(new_n1130), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1172), .A2(new_n1139), .A3(G286), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1162), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(G8), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1151), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1192), .A2(new_n1155), .A3(new_n1187), .A4(new_n1147), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1185), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1155), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1147), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1183), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1033), .B1(new_n1178), .B2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1029), .A2(new_n833), .A3(new_n829), .A4(new_n828), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n733), .A2(new_n1025), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1024), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1024), .A2(G290), .A3(G1986), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT48), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1031), .A2(new_n1203), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1020), .A2(KEYINPUT46), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1020), .A2(KEYINPUT46), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1026), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1017), .B1(new_n1207), .B2(new_n767), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT47), .Z(new_n1210));
  NOR3_X1   g785(.A1(new_n1201), .A2(new_n1204), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1198), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g787(.A(new_n673), .B1(new_n652), .B2(new_n653), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n925), .A2(new_n918), .ZN(new_n1215));
  AOI21_X1  g789(.A(G37), .B1(new_n1215), .B2(new_n882), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1214), .B1(new_n1216), .B2(new_n928), .ZN(new_n1217));
  INV_X1    g791(.A(G319), .ZN(new_n1218));
  NOR2_X1   g792(.A1(G229), .A2(new_n1218), .ZN(new_n1219));
  AND3_X1   g793(.A1(new_n1217), .A2(new_n1001), .A3(new_n1219), .ZN(G308));
  NAND3_X1  g794(.A1(new_n1217), .A2(new_n1001), .A3(new_n1219), .ZN(G225));
endmodule


