//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G234));
  NAND2_X1  g027(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n464), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n471), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n468), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT68), .Z(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(new_n464), .B2(G112), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(new_n470), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n482), .A2(G2105), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n481), .B(new_n485), .C1(G136), .C2(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  OAI21_X1  g063(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT69), .A2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n492), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(KEYINPUT70), .C1(new_n490), .C2(new_n489), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n464), .A2(KEYINPUT71), .A3(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n482), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n464), .A2(KEYINPUT71), .A3(G138), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n465), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n497), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT72), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n497), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n482), .B2(new_n498), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n465), .A2(new_n500), .A3(new_n501), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n493), .A2(new_n495), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n518), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n525), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(new_n517), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n521), .A2(new_n520), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n515), .A2(new_n516), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NAND2_X1  g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n536), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(new_n524), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G90), .B1(G52), .B2(new_n517), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n528), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n517), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n524), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n528), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n524), .A2(KEYINPUT74), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n538), .A2(new_n526), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n517), .A2(G53), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n567), .B(new_n569), .C1(new_n528), .C2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  NAND2_X1  g147(.A1(new_n517), .A2(G49), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n526), .A2(G74), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n528), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n563), .A2(G87), .A3(new_n565), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n563), .A2(KEYINPUT75), .A3(G87), .A4(new_n565), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n537), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G48), .B2(new_n517), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n563), .A2(G86), .A3(new_n565), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n544), .A2(G85), .B1(G47), .B2(new_n517), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n528), .B2(new_n589), .ZN(G290));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NOR2_X1   g166(.A1(G301), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n566), .A2(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT10), .Z(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n537), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n592), .B1(new_n591), .B2(new_n599), .ZN(G284));
  AOI21_X1  g175(.A(new_n592), .B1(new_n591), .B2(new_n599), .ZN(G321));
  NAND2_X1  g176(.A1(G299), .A2(new_n591), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n591), .B2(G168), .ZN(G297));
  XOR2_X1   g178(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(new_n605), .B2(G860), .ZN(G148));
  INV_X1    g181(.A(new_n557), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n591), .ZN(new_n608));
  INV_X1    g183(.A(new_n599), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n610), .B2(new_n591), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n483), .A2(G123), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT77), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(G111), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G2105), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n486), .B2(G135), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n465), .A2(new_n474), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n620), .A2(G2096), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n621), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT78), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  OAI21_X1  g217(.A(G14), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(G401));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT79), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  NOR2_X1   g222(.A1(G2072), .A2(G2078), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n442), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(KEYINPUT17), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n646), .A2(new_n647), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n649), .B(KEYINPUT81), .ZN(new_n657));
  OAI22_X1  g232(.A1(new_n655), .A2(new_n656), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n667), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT20), .Z(new_n671));
  AOI211_X1 g246(.A(new_n669), .B(new_n671), .C1(new_n664), .C2(new_n668), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT83), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1971), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT32), .B(G1981), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n680), .A2(G6), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G305), .B2(G16), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n683), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(G23), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n580), .B2(new_n680), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT33), .B(G1976), .Z(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n687), .A2(new_n685), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n688), .A2(new_n692), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n697));
  MUX2_X1   g272(.A(G24), .B(G290), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1986), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G25), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n486), .A2(G131), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n483), .A2(G119), .ZN(new_n703));
  OR2_X1    g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  OR4_X1    g285(.A1(new_n696), .A2(new_n697), .A3(new_n699), .A4(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT85), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n713), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n700), .A2(G26), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n483), .A2(G128), .ZN(new_n720));
  INV_X1    g295(.A(new_n486), .ZN(new_n721));
  INV_X1    g296(.A(G140), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G104), .A2(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT86), .Z(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n719), .B1(new_n728), .B2(new_n700), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT88), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT87), .B(G2067), .Z(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n700), .A2(G32), .ZN(new_n733));
  AOI22_X1  g308(.A1(G129), .A2(new_n483), .B1(new_n486), .B2(G141), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n474), .A2(G105), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n700), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT93), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G35), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G162), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n732), .B(new_n744), .C1(new_n745), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G168), .A2(new_n680), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n680), .B2(G21), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G19), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n557), .B2(G16), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G1341), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n700), .B1(new_n758), .B2(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G160), .B2(G29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G2084), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n752), .A2(new_n753), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n754), .A2(new_n757), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n749), .A2(new_n745), .B1(new_n730), .B2(new_n731), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n764), .B(new_n765), .C1(new_n743), .C2(new_n742), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n700), .A2(G33), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  INV_X1    g344(.A(G139), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n721), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT89), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n464), .B1(new_n774), .B2(KEYINPUT90), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(KEYINPUT90), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT91), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n767), .B1(new_n778), .B2(new_n700), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G2072), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n750), .A2(new_n766), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n783), .A2(new_n782), .A3(G28), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n782), .B2(G28), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n700), .B1(new_n782), .B2(G28), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT31), .B(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n619), .B2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n756), .A2(G1341), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n761), .A2(G2084), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n789), .B(new_n790), .C1(KEYINPUT95), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G171), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1961), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n792), .B(new_n795), .C1(KEYINPUT95), .C2(new_n791), .ZN(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n512), .A2(new_n700), .ZN(new_n798));
  NOR2_X1   g373(.A1(G27), .A2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n798), .A2(new_n797), .A3(new_n799), .ZN(new_n801));
  NOR2_X1   g376(.A1(G4), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n599), .B2(G16), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n801), .B1(new_n803), .B2(G1348), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n680), .A2(G20), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT23), .Z(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1956), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n803), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n796), .A2(new_n800), .A3(new_n804), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n781), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n537), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n528), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n544), .A2(G93), .B1(G55), .B2(new_n517), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n557), .B1(new_n824), .B2(KEYINPUT98), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n825), .B(new_n826), .Z(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT38), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n599), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT99), .B(G860), .Z(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n822), .B2(new_n823), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n778), .B(new_n739), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n508), .A2(new_n839), .A3(new_n510), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n508), .B2(new_n510), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n838), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n483), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n464), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G142), .B2(new_n486), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n623), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n707), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n728), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n843), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G162), .B(G160), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n620), .ZN(new_n854));
  AOI21_X1  g429(.A(G37), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n852), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g432(.A1(new_n824), .A2(new_n591), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n610), .B(new_n827), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n599), .A2(G299), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n599), .B(G299), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(KEYINPUT101), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n864), .B1(new_n869), .B2(new_n859), .ZN(new_n870));
  XNOR2_X1  g445(.A(G303), .B(KEYINPUT103), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n580), .ZN(new_n872));
  XNOR2_X1  g447(.A(G290), .B(G305), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n872), .B(new_n873), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT42), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n870), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n858), .B1(new_n876), .B2(new_n591), .ZN(G295));
  OAI21_X1  g452(.A(new_n858), .B1(new_n876), .B2(new_n591), .ZN(G331));
  XNOR2_X1  g453(.A(G171), .B(G286), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n827), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n863), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n869), .B2(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n874), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n880), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n863), .B1(new_n865), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n880), .A2(new_n862), .A3(new_n867), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n874), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n882), .A2(new_n883), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(new_n884), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT44), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n891), .B1(new_n884), .B2(new_n888), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(KEYINPUT104), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n891), .A3(new_n884), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n889), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n894), .B1(new_n899), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g475(.A(KEYINPUT127), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT100), .B1(new_n496), .B2(new_n503), .ZN(new_n902));
  INV_X1    g477(.A(G1384), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n508), .A2(new_n839), .A3(new_n510), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(G160), .A2(G40), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G1996), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n739), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT105), .Z(new_n912));
  XNOR2_X1  g487(.A(new_n728), .B(G2067), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n910), .B2(new_n739), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n909), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT106), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n706), .B(new_n709), .Z(new_n918));
  NAND2_X1  g493(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(G290), .A2(G1986), .ZN(new_n920));
  AND2_X1   g495(.A1(G290), .A2(G1986), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n909), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT107), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT119), .ZN(new_n925));
  NAND2_X1  g500(.A1(G286), .A2(G8), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT117), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(KEYINPUT51), .ZN(new_n928));
  INV_X1    g503(.A(G8), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n903), .B1(new_n496), .B2(new_n503), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n908), .B1(new_n930), .B2(new_n906), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n903), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n934), .B2(new_n906), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n753), .ZN(new_n936));
  INV_X1    g511(.A(G2084), .ZN(new_n937));
  AOI21_X1  g512(.A(G1384), .B1(new_n508), .B2(new_n510), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n908), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G1384), .B1(new_n504), .B2(new_n511), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n937), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n929), .B1(new_n936), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n928), .B1(new_n944), .B2(KEYINPUT118), .ZN(new_n945));
  INV_X1    g520(.A(G40), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n468), .A2(new_n476), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n939), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n930), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(KEYINPUT50), .B2(new_n934), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n950), .A2(new_n937), .B1(new_n935), .B2(new_n753), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT118), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n951), .A2(new_n952), .A3(new_n929), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n925), .B1(new_n945), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n951), .B2(new_n929), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n944), .A2(KEYINPUT118), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT119), .A4(new_n928), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT51), .B1(new_n944), .B2(new_n927), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT62), .ZN(new_n960));
  INV_X1    g535(.A(new_n951), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n927), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n960), .B1(new_n959), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n966));
  INV_X1    g541(.A(G1961), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(G2078), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n931), .B(new_n972), .C1(new_n934), .C2(new_n906), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(KEYINPUT120), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n906), .A2(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n908), .B1(new_n842), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n934), .A2(new_n906), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n797), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n971), .ZN(new_n983));
  AOI21_X1  g558(.A(G301), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT55), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G1971), .B1(new_n980), .B2(new_n981), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n745), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(G8), .B(new_n987), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n938), .A2(new_n947), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G8), .ZN(new_n993));
  INV_X1    g568(.A(G1976), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n994), .B(new_n575), .C1(new_n578), .C2(new_n579), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n585), .A2(new_n586), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n517), .A2(G48), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT110), .B(G86), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n538), .A2(new_n526), .A3(new_n1000), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n999), .B(new_n1001), .C1(new_n1002), .C2(new_n528), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G1981), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n998), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n929), .B1(new_n938), .B2(new_n947), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n998), .A2(new_n1004), .A3(KEYINPUT49), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n996), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1012), .B(new_n1013), .C1(new_n580), .C2(G1976), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n578), .A2(new_n579), .ZN(new_n1015));
  INV_X1    g590(.A(new_n575), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(G1976), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1008), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1013), .B1(new_n580), .B2(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(KEYINPUT109), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1011), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n991), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g598(.A(G1971), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT45), .B1(new_n512), .B2(new_n903), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n902), .A2(new_n904), .A3(new_n979), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n947), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n941), .A2(new_n942), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n947), .B1(new_n938), .B2(new_n939), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n745), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n929), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1023), .B1(new_n1033), .B2(new_n987), .ZN(new_n1034));
  AOI211_X1 g609(.A(G2090), .B(new_n1030), .C1(new_n942), .C2(new_n941), .ZN(new_n1035));
  OAI21_X1  g610(.A(G8), .B1(new_n988), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT111), .A3(new_n986), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1022), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n984), .A2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n963), .A2(new_n964), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n944), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n929), .B1(new_n1028), .B2(new_n989), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n987), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1022), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1018), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1019), .A2(KEYINPUT109), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n1014), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n996), .A3(new_n1010), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n987), .B2(new_n1043), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n951), .A2(new_n929), .A3(G286), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT111), .B1(new_n1036), .B2(new_n986), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1033), .A2(new_n1023), .A3(new_n987), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1050), .B(new_n1051), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT112), .B(KEYINPUT63), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1045), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n991), .A2(new_n1049), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1010), .A2(new_n994), .A3(new_n580), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n993), .B1(new_n1058), .B2(new_n998), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1041), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1055), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1038), .B2(new_n1051), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT113), .B(new_n1060), .C1(new_n1064), .C2(new_n1045), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1038), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n959), .B2(new_n962), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n907), .A2(new_n972), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1027), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n980), .A2(KEYINPUT122), .A3(new_n972), .A4(new_n907), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1072), .A2(new_n1073), .B1(new_n971), .B2(new_n982), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n970), .A2(KEYINPUT121), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n966), .A2(new_n1076), .A3(new_n967), .A4(new_n969), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G171), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1069), .B1(new_n984), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1025), .A2(new_n1027), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1956), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1085));
  XNOR2_X1  g660(.A(G299), .B(KEYINPUT57), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  XNOR2_X1  g663(.A(G299), .B(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n808), .B1(new_n1090), .B2(new_n1030), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n980), .A2(new_n981), .A3(new_n1082), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1081), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1086), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT116), .A3(new_n1081), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n966), .A2(new_n811), .A3(new_n969), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n992), .A2(G2067), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n599), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1097), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n609), .A4(new_n1103), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n980), .A2(new_n910), .A3(new_n981), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n992), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1110), .B1(new_n1114), .B2(new_n557), .ZN(new_n1115));
  AOI211_X1 g690(.A(KEYINPUT59), .B(new_n607), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1108), .B(new_n1109), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1101), .A2(new_n1107), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n609), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1098), .B1(new_n1119), .B2(new_n1093), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT115), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1122), .B(new_n1098), .C1(new_n1119), .C2(new_n1093), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1068), .B(new_n1080), .C1(new_n1118), .C2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n970), .A2(KEYINPUT120), .A3(new_n973), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT120), .B1(new_n970), .B2(new_n973), .ZN(new_n1127));
  OAI211_X1 g702(.A(G301), .B(new_n983), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1078), .A2(G171), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT54), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT123), .A4(KEYINPUT54), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1066), .B1(new_n1125), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1040), .B1(new_n1135), .B2(KEYINPUT124), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT116), .B1(new_n1099), .B2(new_n1081), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1095), .B(KEYINPUT61), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1117), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1137), .A2(new_n1145), .A3(new_n1068), .A4(new_n1080), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1147), .A3(new_n1066), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n924), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT46), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n913), .A2(new_n739), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT47), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n909), .A2(new_n920), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT48), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n919), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n707), .A2(new_n709), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT125), .Z(new_n1160));
  INV_X1    g735(.A(G2067), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n917), .A2(new_n1160), .B1(new_n1161), .B2(new_n728), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n909), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1155), .B(new_n1158), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n901), .B1(new_n1149), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1158), .A2(new_n1155), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1164), .A2(new_n909), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1166), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1146), .A2(new_n1147), .A3(new_n1066), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1147), .B1(new_n1146), .B2(new_n1066), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1173), .A2(new_n1174), .A3(new_n1040), .ZN(new_n1175));
  OAI211_X1 g750(.A(KEYINPUT127), .B(new_n1172), .C1(new_n1175), .C2(new_n924), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1168), .A2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g752(.A1(new_n890), .A2(new_n893), .ZN(new_n1179));
  NOR4_X1   g753(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n856), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1181), .ZN(G308));
  INV_X1    g756(.A(G308), .ZN(G225));
endmodule


