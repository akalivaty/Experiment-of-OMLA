//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT70), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(G125), .B(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(KEYINPUT16), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n191), .B(G146), .C1(KEYINPUT16), .C2(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(G128), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n200), .B(new_n202), .C1(new_n203), .C2(KEYINPUT23), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  XNOR2_X1  g019(.A(G119), .B(G128), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n204), .A2(G110), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n198), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT72), .B(G110), .Z(new_n209));
  OAI22_X1  g023(.A1(new_n204), .A2(new_n209), .B1(new_n205), .B2(new_n206), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n190), .A2(new_n195), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n197), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT73), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(new_n212), .A3(new_n218), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n222), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT25), .B1(new_n222), .B2(new_n188), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n189), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n189), .A2(G902), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n222), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  OR3_X1    g051(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT65), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(G137), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n243), .A2(new_n245), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n242), .A2(G137), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n244), .A2(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n195), .A2(G143), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n199), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n195), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n195), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n254), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(KEYINPUT64), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n255), .A2(G143), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G146), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n265), .A2(new_n253), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n252), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n265), .A2(KEYINPUT0), .A3(G128), .A4(new_n253), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT0), .B(G128), .Z(new_n270));
  AOI21_X1  g084(.A(G146), .B1(new_n263), .B2(new_n264), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(new_n260), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT11), .B1(new_n244), .B2(G134), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n250), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n246), .B1(new_n274), .B2(new_n245), .ZN(new_n275));
  INV_X1    g089(.A(new_n248), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n269), .B(new_n272), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n268), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n268), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n240), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT26), .B(G101), .Z(new_n283));
  INV_X1    g097(.A(G237), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(new_n214), .A3(G210), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n290), .B(new_n240), .C1(new_n279), .C2(new_n280), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n268), .A2(new_n277), .A3(new_n238), .A4(new_n239), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n282), .A2(new_n289), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT31), .ZN(new_n294));
  INV_X1    g108(.A(new_n292), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n281), .B2(KEYINPUT66), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n289), .A4(new_n291), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n268), .A2(new_n277), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n240), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n301), .B2(new_n292), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n292), .A2(new_n299), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT68), .B1(new_n304), .B2(new_n289), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n288), .C1(new_n302), .C2(new_n303), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n294), .A2(new_n298), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G472), .A2(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT69), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n315), .A3(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G472), .ZN(new_n318));
  INV_X1    g132(.A(new_n304), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(new_n288), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(KEYINPUT29), .ZN(new_n321));
  INV_X1    g135(.A(new_n296), .ZN(new_n322));
  INV_X1    g136(.A(new_n291), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n288), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n188), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n320), .B2(KEYINPUT29), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n318), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n231), .B1(new_n317), .B2(new_n329), .ZN(new_n330));
  AOI211_X1 g144(.A(KEYINPUT71), .B(new_n328), .C1(new_n314), .C2(new_n316), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n230), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  INV_X1    g147(.A(G224), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT7), .B1(new_n334), .B2(G953), .ZN(new_n335));
  INV_X1    g149(.A(new_n254), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n271), .B2(new_n260), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n265), .A2(new_n253), .A3(new_n266), .ZN(new_n338));
  AOI21_X1  g152(.A(G125), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n272), .A2(G125), .A3(new_n269), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n272), .A2(G125), .A3(new_n269), .ZN(new_n342));
  INV_X1    g156(.A(new_n335), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n262), .A2(new_n267), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n201), .A2(G116), .ZN(new_n349));
  INV_X1    g163(.A(G116), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G119), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT5), .ZN(new_n352));
  OAI21_X1  g166(.A(G113), .B1(new_n349), .B2(KEYINPUT5), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n237), .A2(KEYINPUT5), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n350), .A2(G119), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n232), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(KEYINPUT77), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n236), .A2(new_n237), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(new_n362), .B2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G104), .ZN(new_n366));
  INV_X1    g180(.A(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(G107), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n366), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n362), .A2(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n365), .A2(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(G101), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n361), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n347), .B1(new_n360), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n363), .A2(new_n366), .A3(new_n368), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(G101), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n240), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n373), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n381), .A2(KEYINPUT78), .A3(new_n359), .A4(new_n354), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G122), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n374), .A2(new_n380), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n346), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n383), .B(KEYINPUT8), .Z(new_n386));
  OR2_X1    g200(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n353), .B1(new_n355), .B2(KEYINPUT79), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n373), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n354), .A2(new_n359), .A3(new_n361), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n369), .A2(new_n372), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n389), .B1(new_n392), .B2(KEYINPUT80), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n394), .A3(new_n391), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n386), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n333), .B1(new_n385), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT81), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n374), .A2(new_n380), .A3(new_n382), .ZN(new_n399));
  INV_X1    g213(.A(new_n383), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n384), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n339), .A2(new_n340), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n334), .A2(G953), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n409), .B(new_n333), .C1(new_n385), .C2(new_n396), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n398), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G210), .B1(G237), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n398), .A2(new_n412), .A3(new_n408), .A4(new_n410), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G214), .B1(G237), .B2(G902), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n416), .A2(new_n415), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT83), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(new_n419), .A3(new_n422), .A4(new_n418), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT9), .B(G234), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n425), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(new_n333), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT10), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n265), .A2(new_n253), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT1), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n263), .A2(new_n264), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(new_n195), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n432), .B1(new_n435), .B2(new_n199), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n267), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(KEYINPUT75), .B(new_n432), .C1(new_n435), .C2(new_n199), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n431), .B(new_n391), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n436), .A2(new_n437), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n338), .A3(new_n439), .ZN(new_n442));
  INV_X1    g256(.A(new_n391), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT76), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n430), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n275), .A2(new_n276), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n344), .A2(new_n430), .A3(new_n391), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n379), .A2(new_n377), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n272), .A2(new_n269), .ZN(new_n450));
  OR3_X1    g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n448), .B2(new_n450), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n445), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G140), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n214), .A2(G227), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT12), .ZN(new_n460));
  INV_X1    g274(.A(new_n344), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n443), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n442), .A2(new_n443), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n431), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n442), .A2(KEYINPUT76), .A3(new_n443), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n460), .B1(new_n466), .B2(new_n446), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n440), .A2(new_n444), .B1(new_n461), .B2(new_n443), .ZN(new_n468));
  INV_X1    g282(.A(new_n446), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(KEYINPUT12), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n459), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT10), .B1(new_n464), .B2(new_n465), .ZN(new_n473));
  INV_X1    g287(.A(new_n453), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n454), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n457), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n326), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n429), .B1(new_n478), .B2(new_n428), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n454), .A3(new_n458), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n473), .A2(new_n474), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n467), .A2(new_n470), .B1(new_n481), .B2(new_n446), .ZN(new_n482));
  OAI211_X1 g296(.A(G469), .B(new_n480), .C1(new_n482), .C2(new_n458), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n427), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n190), .B(new_n195), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n284), .A2(new_n214), .A3(G214), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n263), .A3(new_n264), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n284), .A2(new_n214), .A3(G143), .A4(G214), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT84), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n496), .B(new_n493), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n488), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g312(.A1(KEYINPUT85), .A2(KEYINPUT18), .A3(G131), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT85), .B1(KEYINPUT18), .B2(G131), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n490), .A2(new_n501), .A3(new_n491), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n490), .A2(new_n501), .A3(KEYINPUT86), .A4(new_n491), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n487), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n492), .A2(new_n494), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n496), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n492), .A2(KEYINPUT84), .A3(new_n494), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n504), .A2(new_n505), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n511), .A2(KEYINPUT87), .A3(new_n512), .A4(new_n488), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G125), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G140), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n193), .A2(new_n516), .A3(KEYINPUT19), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT19), .B1(new_n193), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT88), .B1(new_n519), .B2(G146), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n521), .B(new_n195), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n492), .A2(G131), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n246), .B1(new_n490), .B2(new_n491), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n197), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT89), .B1(new_n514), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G113), .B(G122), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n362), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n507), .B2(new_n513), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n198), .B1(KEYINPUT17), .B2(new_n525), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n524), .A2(new_n525), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(KEYINPUT17), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n507), .A2(new_n513), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n530), .B(KEYINPUT90), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n486), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT91), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n540), .B1(new_n528), .B2(new_n533), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n545), .B(KEYINPUT20), .C1(new_n546), .C2(new_n486), .ZN(new_n547));
  INV_X1    g361(.A(new_n546), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n485), .B(KEYINPUT92), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n537), .A2(new_n538), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n530), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n333), .B1(new_n553), .B2(new_n540), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G475), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n199), .A2(G143), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n434), .B2(new_n199), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G134), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n350), .A2(G122), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n365), .B1(new_n560), .B2(KEYINPUT14), .ZN(new_n561));
  XNOR2_X1  g375(.A(G116), .B(G122), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT14), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n561), .A2(new_n564), .B1(new_n365), .B2(new_n562), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT64), .B(G143), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(G128), .ZN(new_n569));
  OAI211_X1 g383(.A(G134), .B(new_n569), .C1(new_n558), .C2(new_n568), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n562), .B(new_n365), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n570), .B(new_n571), .C1(G134), .C2(new_n558), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n425), .A2(new_n187), .A3(G953), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT93), .Z(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT94), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n573), .B2(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n575), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n188), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n581), .B(new_n188), .C1(KEYINPUT15), .C2(new_n583), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G952), .ZN(new_n588));
  AOI211_X1 g402(.A(G953), .B(new_n588), .C1(G234), .C2(G237), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n214), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT21), .B(G898), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n424), .A2(new_n484), .A3(new_n556), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n332), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n367), .ZN(G3));
  NAND2_X1  g410(.A1(new_n454), .A2(new_n458), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n470), .B2(new_n467), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n458), .B1(new_n475), .B2(new_n454), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n428), .B(new_n188), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n429), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n483), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n426), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n308), .A2(new_n309), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n318), .B1(new_n308), .B2(new_n188), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n603), .A2(new_n229), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n551), .A2(new_n555), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n576), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n581), .A2(new_n610), .B1(new_n580), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n326), .A2(new_n583), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(KEYINPUT95), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n582), .A2(new_n583), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT95), .B1(new_n612), .B2(new_n613), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n418), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n414), .B2(new_n416), .ZN(new_n621));
  INV_X1    g435(.A(new_n592), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n608), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NAND3_X1  g440(.A1(new_n548), .A2(new_n543), .A3(new_n485), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n544), .A2(new_n547), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n555), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n608), .A2(new_n587), .A3(new_n623), .A4(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n219), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n213), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n226), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n225), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n555), .A2(new_n551), .A3(new_n593), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n424), .A2(new_n484), .A3(new_n637), .A4(new_n606), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT96), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT37), .B(G110), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  NAND4_X1  g455(.A1(new_n602), .A2(new_n426), .A3(new_n621), .A4(new_n636), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n590), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n589), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n628), .A2(new_n555), .A3(new_n587), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n330), .B2(new_n331), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n646), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n484), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT97), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n322), .A2(new_n323), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n288), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n301), .A2(new_n288), .A3(new_n292), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n333), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n317), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n417), .A2(new_n419), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT38), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n609), .A2(new_n587), .A3(new_n418), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n664), .A2(new_n636), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n655), .A2(new_n656), .A3(new_n662), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n567), .B(KEYINPUT98), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G45));
  NAND3_X1  g483(.A1(new_n609), .A2(new_n618), .A3(new_n646), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n642), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n330), .B2(new_n331), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  NAND3_X1  g487(.A1(new_n623), .A2(new_n609), .A3(new_n618), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n471), .A2(new_n459), .B1(new_n476), .B2(new_n457), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n675), .B2(new_n326), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n426), .A3(new_n600), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n678), .B(new_n230), .C1(new_n330), .C2(new_n331), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  AND4_X1   g495(.A1(new_n230), .A2(new_n629), .A3(new_n622), .A4(new_n587), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n426), .A3(new_n600), .A4(new_n621), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n682), .B(new_n684), .C1(new_n330), .C2(new_n331), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  OAI211_X1 g500(.A(new_n637), .B(new_n684), .C1(new_n330), .C2(new_n331), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  NAND2_X1  g502(.A1(new_n587), .A2(new_n418), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n414), .A2(new_n416), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n689), .B(new_n690), .C1(new_n551), .C2(new_n555), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n622), .A2(new_n676), .A3(new_n426), .A4(new_n600), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n309), .B(KEYINPUT99), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n293), .A2(KEYINPUT31), .B1(new_n319), .B2(new_n288), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n298), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n694), .B2(new_n695), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n693), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n699), .A2(new_n229), .A3(new_n605), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n691), .A2(new_n692), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  INV_X1    g516(.A(new_n670), .ZN(new_n703));
  INV_X1    g517(.A(new_n636), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n699), .A2(new_n605), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n684), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  NAND2_X1  g521(.A1(new_n313), .A2(KEYINPUT69), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT32), .B1(new_n308), .B2(new_n309), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n316), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n329), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT71), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n317), .A2(new_n231), .A3(new_n329), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n483), .A2(KEYINPUT101), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n466), .A2(new_n460), .A3(new_n446), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT12), .B1(new_n468), .B2(new_n469), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n454), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n457), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT101), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n721), .A3(G469), .A4(new_n480), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n716), .A2(new_n600), .A3(new_n722), .A4(new_n601), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n620), .B1(new_n417), .B2(new_n419), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n426), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n670), .A2(KEYINPUT42), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n715), .A2(new_n230), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n328), .A2(new_n709), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n229), .B1(new_n729), .B2(new_n313), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n703), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n731), .B2(new_n725), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(KEYINPUT102), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT102), .B1(new_n728), .B2(new_n732), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  AOI211_X1 g551(.A(new_n229), .B(new_n725), .C1(new_n713), .C2(new_n714), .ZN(new_n738));
  INV_X1    g552(.A(new_n647), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NAND3_X1  g555(.A1(new_n720), .A2(KEYINPUT45), .A3(new_n480), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT45), .B1(new_n720), .B2(new_n480), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n428), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(new_n429), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  OR3_X1    g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n747), .B1(new_n746), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n748), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n600), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(new_n426), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n651), .ZN(new_n754));
  INV_X1    g568(.A(new_n724), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n556), .A2(new_n618), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n607), .A3(new_n636), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n244), .ZN(G39));
  INV_X1    g577(.A(new_n715), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n755), .A2(new_n230), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n703), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n752), .A2(new_n426), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n766), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n192), .ZN(G42));
  NAND2_X1  g586(.A1(new_n676), .A2(new_n600), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT104), .Z(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT49), .Z(new_n775));
  NOR2_X1   g589(.A1(new_n662), .A2(new_n229), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n756), .A2(new_n620), .A3(new_n427), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n664), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n608), .A2(new_n622), .A3(new_n424), .A4(new_n619), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n332), .B2(new_n594), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n780), .B(KEYINPUT105), .C1(new_n332), .C2(new_n594), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n728), .A2(new_n732), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT102), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n685), .A2(new_n679), .A3(new_n687), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n638), .A2(new_n701), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n421), .A2(new_n423), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n604), .A2(new_n605), .A3(new_n229), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n602), .A3(new_n622), .A4(new_n426), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n587), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n585), .A2(KEYINPUT106), .A3(new_n586), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n556), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n791), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n785), .A2(new_n788), .A3(new_n801), .A4(new_n733), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n723), .A2(new_n426), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n646), .B(KEYINPUT108), .Z(new_n804));
  NAND2_X1  g618(.A1(new_n704), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT109), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n803), .A2(new_n662), .A3(new_n806), .A4(new_n691), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n649), .A2(new_n672), .A3(new_n706), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n809));
  INV_X1    g623(.A(new_n705), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n670), .A3(new_n683), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n715), .B2(new_n648), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n672), .A4(new_n807), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n725), .A2(new_n810), .A3(new_n670), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n738), .B2(new_n739), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n795), .A2(new_n796), .B1(new_n645), .B2(new_n644), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n724), .A2(new_n817), .A3(new_n555), .A4(new_n628), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n603), .A3(new_n704), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n331), .B2(new_n330), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT107), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT107), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n715), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n809), .A2(new_n814), .A3(new_n816), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n779), .B1(new_n802), .B2(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n814), .A2(new_n809), .A3(new_n824), .A4(new_n816), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n790), .A2(new_n799), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n679), .A3(new_n685), .A4(new_n687), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n783), .B2(new_n784), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n736), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  INV_X1    g647(.A(new_n786), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n834), .A4(new_n830), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n826), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n840), .A3(KEYINPUT54), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n839), .B1(new_n838), .B2(new_n841), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n755), .A2(new_n677), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n677), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT114), .B1(new_n846), .B2(new_n724), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n845), .A2(new_n645), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n757), .A3(new_n730), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT48), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n588), .A2(G953), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n700), .A2(new_n589), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n757), .A2(new_n684), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT115), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n619), .A3(new_n776), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n851), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT116), .Z(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n774), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n774), .A2(new_n858), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n427), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n767), .A2(new_n770), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n757), .A2(new_n852), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n755), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n848), .A2(new_n757), .A3(new_n705), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n609), .A2(new_n618), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n848), .A2(new_n776), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n664), .A2(new_n620), .A3(new_n846), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(KEYINPUT50), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n864), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n868), .B(new_n870), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AND4_X1   g691(.A1(KEYINPUT113), .A2(new_n866), .A3(new_n867), .A4(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n872), .B(KEYINPUT50), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n868), .A4(new_n870), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n866), .A2(new_n877), .B1(new_n881), .B2(new_n867), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n857), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n842), .A2(new_n843), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n588), .A2(new_n214), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT117), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n778), .B1(new_n884), .B2(new_n886), .ZN(G75));
  AOI21_X1  g701(.A(new_n188), .B1(new_n826), .B2(new_n835), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(new_n413), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n407), .B(KEYINPUT55), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n413), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n402), .A2(new_n404), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT118), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n214), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n891), .B2(new_n894), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(G51));
  NAND2_X1  g717(.A1(new_n826), .A2(new_n835), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n326), .A3(new_n745), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT120), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n837), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n429), .B(KEYINPUT57), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n675), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n899), .B1(new_n912), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(new_n546), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n899), .B1(new_n915), .B2(new_n546), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G60));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n908), .A2(new_n612), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n900), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n842), .B2(new_n843), .ZN(new_n926));
  INV_X1    g740(.A(new_n612), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT60), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n904), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n899), .B1(new_n931), .B2(new_n228), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT61), .B1(new_n932), .B2(KEYINPUT122), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n904), .A2(new_n634), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G66));
  NOR2_X1   g750(.A1(new_n591), .A2(new_n334), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n214), .ZN(new_n938));
  INV_X1    g752(.A(new_n830), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n214), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n896), .B1(G898), .B2(new_n214), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT123), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n940), .B(new_n942), .ZN(G69));
  AOI21_X1  g757(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n812), .A2(new_n672), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT124), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n667), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT62), .Z(new_n948));
  AOI21_X1  g762(.A(new_n619), .B1(new_n556), .B2(new_n797), .ZN(new_n949));
  OR4_X1    g763(.A1(new_n332), .A2(new_n949), .A3(new_n652), .A4(new_n755), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n754), .B2(new_n761), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT125), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n953), .B(new_n950), .C1(new_n754), .C2(new_n761), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n771), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(G953), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n279), .A2(new_n280), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n519), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(G900), .A2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n730), .A2(new_n691), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n753), .A2(new_n651), .A3(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n963), .B(new_n740), .C1(new_n754), .C2(new_n761), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n945), .B(KEYINPUT124), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n767), .A2(new_n770), .ZN(new_n967));
  INV_X1    g781(.A(new_n766), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n965), .A2(new_n736), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n961), .B1(new_n970), .B2(new_n214), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n944), .B1(new_n959), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  INV_X1    g787(.A(new_n944), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n973), .B(new_n974), .C1(new_n956), .C2(new_n958), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(new_n975), .ZN(G72));
  NAND4_X1  g790(.A1(new_n965), .A2(new_n969), .A3(new_n736), .A4(new_n830), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  XNOR2_X1  g792(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n318), .A2(new_n333), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(new_n981));
  AND3_X1   g795(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n978), .B1(new_n977), .B2(new_n981), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n288), .B(new_n657), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n948), .A2(new_n830), .A3(new_n955), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n658), .ZN(new_n987));
  INV_X1    g801(.A(new_n981), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n324), .B2(new_n293), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n899), .B1(new_n832), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n984), .A2(new_n987), .A3(new_n990), .ZN(G57));
endmodule


