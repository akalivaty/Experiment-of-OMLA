//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n567, new_n569, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n464), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n476), .B1(new_n481), .B2(G124), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT69), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(KEYINPUT4), .A2(G138), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n477), .B2(new_n478), .ZN(new_n486));
  NAND2_X1  g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n465), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n477), .B2(new_n478), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n465), .C1(new_n461), .C2(new_n462), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n489), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G62), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n501), .A2(new_n502), .B1(G75), .B2(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n500), .A2(KEYINPUT71), .A3(G62), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT70), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT5), .B(G543), .Z(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n509), .B2(new_n511), .ZN(new_n514));
  AOI22_X1  g089(.A1(G50), .A2(new_n512), .B1(new_n514), .B2(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n507), .A2(new_n515), .A3(KEYINPUT72), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n514), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n512), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(new_n525), .B1(new_n500), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n513), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(new_n506), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT73), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n514), .A2(G90), .ZN(new_n536));
  INV_X1    g111(.A(new_n512), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT74), .B(G52), .Z(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n534), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n535), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n513), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n514), .A2(G81), .B1(new_n546), .B2(new_n506), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT76), .B(G43), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n512), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT77), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n513), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n514), .A2(G91), .B1(new_n560), .B2(G651), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n512), .A2(new_n562), .A3(G53), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n562), .B1(new_n512), .B2(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT78), .ZN(G299));
  OR2_X1    g141(.A1(new_n539), .A2(new_n535), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n567), .A2(new_n541), .A3(new_n534), .ZN(G301));
  XNOR2_X1  g143(.A(new_n528), .B(KEYINPUT79), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G286));
  INV_X1    g145(.A(new_n519), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT72), .B1(new_n507), .B2(new_n515), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  NAND2_X1  g148(.A1(new_n512), .A2(G49), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n514), .A2(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n512), .A2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n514), .A2(G86), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  INV_X1    g155(.A(new_n506), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n514), .A2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n512), .A2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n581), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n514), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n513), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n512), .A2(G54), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT80), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G286), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n565), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT81), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n606), .B1(new_n609), .B2(new_n605), .ZN(G297));
  AOI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n605), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n550), .A2(new_n605), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n601), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g192(.A(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n479), .A2(new_n466), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n464), .B2(G135), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(new_n481), .B2(G123), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n618), .A2(new_n621), .B1(new_n628), .B2(G2096), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n629), .B(new_n630), .C1(new_n618), .C2(new_n621), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT83), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(KEYINPUT17), .ZN(new_n656));
  INV_X1    g231(.A(new_n650), .ZN(new_n657));
  INV_X1    g232(.A(new_n651), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n653), .A3(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(new_n652), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n655), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(new_n670), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n672), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n675));
  OAI221_X1 g250(.A(new_n671), .B1(new_n673), .B2(new_n667), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n674), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1981), .ZN(new_n678));
  INV_X1    g253(.A(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT87), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  XOR2_X1   g263(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G20), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n608), .B2(new_n690), .ZN(new_n693));
  INV_X1    g268(.A(G1956), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G35), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G162), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT29), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G2090), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n695), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT99), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n690), .A2(G4), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n602), .B2(new_n690), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT91), .B(G1348), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT25), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n464), .A2(G139), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n709), .B(new_n710), .C1(new_n465), .C2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT92), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G29), .B2(G33), .ZN(new_n715));
  INV_X1    g290(.A(G2072), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n464), .A2(G141), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n466), .A2(G105), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT26), .Z(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n481), .B2(G129), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(new_n696), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n696), .B2(G32), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT27), .B(G1996), .ZN(new_n727));
  AND2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  NOR2_X1   g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n696), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G160), .B2(G29), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n726), .A2(new_n727), .B1(G2084), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n717), .A2(new_n718), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n707), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n690), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n690), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT30), .B(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  NAND2_X1  g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n741), .A2(new_n696), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n628), .B2(new_n696), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT95), .Z(new_n746));
  NOR2_X1   g321(.A1(G171), .A2(new_n690), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G5), .B2(new_n690), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n740), .B(new_n746), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n732), .A2(G2084), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT97), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n550), .A2(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n690), .A2(G19), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n753), .B1(G1341), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n748), .A2(new_n749), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  NOR2_X1   g335(.A1(G27), .A2(G29), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G164), .B2(G29), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n726), .A2(new_n727), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n760), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n696), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n464), .A2(G140), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n465), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n481), .B2(G128), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(new_n696), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2067), .ZN(new_n774));
  INV_X1    g349(.A(G1341), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n756), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n758), .A2(new_n759), .A3(new_n765), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n701), .B2(new_n700), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n736), .A2(new_n751), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n703), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(G16), .A2(G24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G290), .B2(new_n690), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(new_n679), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n696), .A2(G25), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n481), .A2(G119), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n464), .A2(G131), .ZN(new_n786));
  NOR2_X1   g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT88), .Z(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n784), .B1(new_n792), .B2(new_n696), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT35), .B(G1991), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n782), .A2(new_n679), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G6), .A2(G16), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  INV_X1    g377(.A(G1981), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n690), .A2(G22), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT89), .Z(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n690), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G1971), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(G1971), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n690), .A2(G23), .ZN(new_n810));
  INV_X1    g385(.A(G288), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n690), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT33), .B(G1976), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n804), .A2(new_n808), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n783), .B(new_n798), .C1(new_n815), .C2(KEYINPUT34), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT90), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n780), .B1(new_n820), .B2(new_n822), .ZN(G311));
  INV_X1    g398(.A(G311), .ZN(G150));
  NAND2_X1  g399(.A1(new_n514), .A2(G93), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT100), .B(G55), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n825), .B1(new_n581), .B2(new_n826), .C1(new_n537), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT101), .B(G860), .Z(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NOR2_X1   g407(.A1(new_n601), .A2(new_n612), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n828), .B(new_n550), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT39), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n829), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n832), .B1(new_n840), .B2(new_n841), .ZN(G145));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n713), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n724), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n464), .A2(G142), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n465), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n481), .B2(G130), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n620), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n772), .B(G164), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n791), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n627), .B(G160), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n483), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n857), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n859), .A2(KEYINPUT104), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(KEYINPUT104), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(G395));
  XNOR2_X1  g439(.A(G166), .B(G288), .ZN(new_n865));
  XNOR2_X1  g440(.A(G290), .B(G305), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n615), .B(new_n836), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n608), .A2(new_n596), .ZN(new_n872));
  NAND2_X1  g447(.A1(G299), .A2(new_n597), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n872), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n874), .B2(KEYINPUT41), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n877), .A2(KEYINPUT42), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n885));
  INV_X1    g460(.A(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n870), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT42), .B1(new_n877), .B2(new_n883), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n885), .A3(new_n876), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n869), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G868), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n828), .A2(new_n605), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(G295));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n896), .A3(new_n894), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n605), .B1(new_n888), .B2(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT108), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(G331));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n902));
  NAND2_X1  g477(.A1(G171), .A2(new_n569), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n528), .B1(new_n540), .B2(new_n542), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n835), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n835), .B1(new_n903), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n881), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n904), .B1(G286), .B2(G301), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n836), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n911), .A2(new_n905), .B1(new_n872), .B2(new_n873), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n869), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT109), .B1(new_n914), .B2(G37), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n912), .B1(new_n881), .B2(new_n908), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n869), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n869), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n908), .B(new_n924), .C1(new_n874), .C2(new_n879), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(new_n870), .C1(new_n875), .C2(new_n908), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n917), .A3(new_n920), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n927), .A2(new_n922), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n902), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT44), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT110), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n917), .B1(new_n918), .B2(new_n869), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n934), .A2(KEYINPUT109), .B1(new_n869), .B2(new_n918), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT43), .B1(new_n935), .B2(new_n919), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n927), .A2(new_n922), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n922), .B1(new_n935), .B2(new_n919), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n938), .B(new_n939), .C1(new_n942), .C2(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n943), .ZN(G397));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n498), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT45), .B1(new_n946), .B2(KEYINPUT111), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(KEYINPUT111), .B2(new_n946), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT112), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT46), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT46), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n772), .B(G2067), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n724), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT47), .Z(new_n960));
  NOR2_X1   g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n951), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n962), .A2(KEYINPUT48), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(KEYINPUT48), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n724), .B(G1996), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n956), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n791), .A2(new_n795), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n792), .A2(new_n794), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n951), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n963), .A2(new_n964), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n772), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n966), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n968), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n951), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT127), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n960), .A2(new_n971), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(G290), .B(G1986), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n951), .B1(new_n969), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT113), .ZN(new_n981));
  INV_X1    g556(.A(new_n485), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n461), .B2(new_n462), .ZN(new_n983));
  AOI21_X1  g558(.A(G2105), .B1(new_n983), .B2(new_n487), .ZN(new_n984));
  OAI21_X1  g559(.A(G126), .B1(new_n461), .B2(new_n462), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n465), .B1(new_n985), .B2(new_n492), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n987), .B2(new_n497), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n949), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2084), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n993), .B(new_n989), .C1(new_n498), .C2(new_n945), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n990), .B(new_n991), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n993), .B1(new_n988), .B2(new_n989), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n946), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(KEYINPUT118), .A3(new_n991), .A4(new_n990), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n946), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n739), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n997), .A2(new_n1001), .A3(G168), .A4(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT123), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n997), .A2(new_n1001), .A3(new_n1007), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1008), .A2(G8), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n995), .A2(new_n996), .B1(new_n739), .B2(new_n1006), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n1001), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(KEYINPUT51), .C1(new_n1010), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n528), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT62), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1014), .A2(new_n1019), .A3(new_n1023), .A4(new_n1020), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n803), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(KEYINPUT49), .A3(new_n1026), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1016), .B1(new_n988), .B2(new_n1004), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1033), .B2(G288), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1033), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1031), .B(new_n1036), .C1(new_n1033), .C2(G288), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(G166), .B2(new_n1016), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1000), .A2(new_n701), .A3(new_n990), .ZN(new_n1043));
  INV_X1    g618(.A(G1971), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1006), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1016), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n946), .A2(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n990), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n990), .A2(KEYINPUT117), .A3(new_n1048), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n701), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1016), .B1(new_n1053), .B2(new_n1045), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1038), .B(new_n1047), .C1(new_n1054), .C2(new_n1042), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n990), .B1(new_n992), .B2(new_n994), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n749), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1006), .B2(G2078), .ZN(new_n1059));
  AND4_X1   g634(.A1(KEYINPUT53), .A2(new_n1005), .A3(new_n1004), .A4(new_n760), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1003), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G171), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1055), .A2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1022), .A2(new_n1024), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1038), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G288), .A2(G1976), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1067), .B(KEYINPUT115), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1032), .A2(new_n1068), .B1(new_n803), .B2(new_n800), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1031), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1066), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1018), .A2(new_n569), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1055), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1075), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n1074), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(new_n1079), .A3(new_n1047), .A4(new_n1038), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1073), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1049), .A2(new_n694), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n565), .B(KEYINPUT57), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n988), .A2(new_n1004), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(G2067), .ZN(new_n1092));
  INV_X1    g667(.A(G1348), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n1056), .B2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1094), .A2(new_n596), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n597), .B1(new_n1094), .B2(KEYINPUT60), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT122), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n597), .C1(new_n1094), .C2(KEYINPUT60), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1091), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT120), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1091), .A2(new_n1109), .A3(new_n1106), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1108), .B(new_n1110), .C1(G1996), .C2(new_n1006), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1111), .A2(new_n551), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1111), .B2(new_n551), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1089), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n1085), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT61), .B1(new_n1118), .B2(new_n1090), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1116), .A3(new_n1085), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1096), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1115), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1097), .B1(new_n1105), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n948), .A2(new_n1060), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1057), .A2(new_n1059), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G171), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1057), .A2(G301), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(KEYINPUT54), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1127), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1128), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1057), .A2(new_n1125), .A3(new_n1059), .A4(G301), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT54), .B1(new_n1063), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1055), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1021), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1081), .B1(new_n1124), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1065), .B1(new_n1138), .B2(KEYINPUT125), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1081), .B(new_n1140), .C1(new_n1124), .C2(new_n1137), .ZN(new_n1141));
  AOI211_X1 g716(.A(KEYINPUT126), .B(new_n981), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1138), .A2(KEYINPUT125), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1065), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n981), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n978), .B1(new_n1142), .B2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g724(.A(G319), .ZN(new_n1151));
  NOR3_X1   g725(.A1(G401), .A2(new_n1151), .A3(G227), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n862), .A2(new_n687), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n1153), .A2(new_n942), .ZN(G308));
  INV_X1    g728(.A(G308), .ZN(G225));
endmodule


