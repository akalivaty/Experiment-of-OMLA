

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U550 ( .A1(n738), .A2(G2084), .ZN(n737) );
  XNOR2_X2 U551 ( .A(n737), .B(n736), .ZN(n762) );
  INV_X2 U552 ( .A(n738), .ZN(n717) );
  XNOR2_X2 U553 ( .A(n710), .B(KEYINPUT64), .ZN(n738) );
  AND2_X1 U554 ( .A1(n516), .A2(n849), .ZN(n850) );
  AND2_X1 U555 ( .A1(n518), .A2(n839), .ZN(n517) );
  OR2_X1 U556 ( .A1(n722), .A2(n527), .ZN(n526) );
  INV_X1 U557 ( .A(KEYINPUT105), .ZN(n532) );
  NOR2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n548) );
  NAND2_X1 U559 ( .A1(n519), .A2(n517), .ZN(n516) );
  AND2_X1 U560 ( .A1(n775), .A2(n788), .ZN(n789) );
  XNOR2_X1 U561 ( .A(n770), .B(n532), .ZN(n775) );
  NOR2_X1 U562 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U563 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U564 ( .A1(n528), .A2(n726), .ZN(n531) );
  XNOR2_X1 U565 ( .A(n715), .B(n529), .ZN(n528) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n815) );
  OR2_X1 U567 ( .A1(G2090), .A2(n787), .ZN(n788) );
  INV_X1 U568 ( .A(n562), .ZN(n524) );
  NOR2_X1 U569 ( .A1(n562), .A2(n521), .ZN(n520) );
  INV_X1 U570 ( .A(n525), .ZN(n522) );
  AND2_X1 U571 ( .A1(n910), .A2(G137), .ZN(n525) );
  NOR2_X2 U572 ( .A1(G2105), .A2(n550), .ZN(n557) );
  INV_X1 U573 ( .A(KEYINPUT101), .ZN(n529) );
  NAND2_X1 U574 ( .A1(n790), .A2(n795), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n786), .A2(n988), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n522), .A2(n520), .ZN(n814) );
  NAND2_X1 U577 ( .A1(n559), .A2(G40), .ZN(n521) );
  NOR2_X1 U578 ( .A1(n523), .A2(n525), .ZN(G160) );
  NAND2_X1 U579 ( .A1(n524), .A2(n559), .ZN(n523) );
  AND2_X1 U580 ( .A1(n729), .A2(n526), .ZN(n530) );
  INV_X1 U581 ( .A(n726), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n730) );
  INV_X1 U583 ( .A(KEYINPUT106), .ZN(n784) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n673) );
  XOR2_X1 U585 ( .A(KEYINPUT32), .B(KEYINPUT104), .Z(n533) );
  NOR2_X1 U586 ( .A1(n996), .A2(n714), .ZN(n716) );
  AND2_X1 U587 ( .A1(n742), .A2(n741), .ZN(n745) );
  NOR2_X1 U588 ( .A1(n745), .A2(n744), .ZN(n746) );
  INV_X1 U589 ( .A(KEYINPUT103), .ZN(n750) );
  XNOR2_X1 U590 ( .A(n761), .B(n533), .ZN(n769) );
  INV_X1 U591 ( .A(KEYINPUT5), .ZN(n542) );
  XNOR2_X1 U592 ( .A(n542), .B(KEYINPUT74), .ZN(n543) );
  NOR2_X1 U593 ( .A1(n661), .A2(n539), .ZN(n674) );
  AND2_X1 U594 ( .A1(n550), .A2(G2105), .ZN(n905) );
  XNOR2_X1 U595 ( .A(n544), .B(n543), .ZN(n545) );
  AND2_X1 U596 ( .A1(n556), .A2(n555), .ZN(G164) );
  XOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .Z(n661) );
  NOR2_X1 U598 ( .A1(G651), .A2(n661), .ZN(n668) );
  NAND2_X1 U599 ( .A1(G51), .A2(n668), .ZN(n536) );
  INV_X1 U600 ( .A(G651), .ZN(n539) );
  NOR2_X1 U601 ( .A1(G543), .A2(n539), .ZN(n534) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n534), .Z(n669) );
  NAND2_X1 U603 ( .A1(G63), .A2(n669), .ZN(n535) );
  NAND2_X1 U604 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U605 ( .A(KEYINPUT6), .B(n537), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n673), .A2(G89), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n538), .B(KEYINPUT4), .ZN(n541) );
  NAND2_X1 U608 ( .A1(G76), .A2(n674), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U611 ( .A(KEYINPUT7), .B(n547), .Z(G168) );
  XOR2_X2 U612 ( .A(KEYINPUT17), .B(n548), .Z(n910) );
  NAND2_X1 U613 ( .A1(n910), .A2(G138), .ZN(n556) );
  INV_X1 U614 ( .A(G2104), .ZN(n550) );
  NAND2_X1 U615 ( .A1(G126), .A2(n905), .ZN(n549) );
  XNOR2_X1 U616 ( .A(KEYINPUT89), .B(n549), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G102), .A2(n557), .ZN(n552) );
  AND2_X1 U618 ( .A1(G2104), .A2(G2105), .ZN(n906) );
  NAND2_X1 U619 ( .A1(G114), .A2(n906), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U622 ( .A1(G101), .A2(n557), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT23), .B(n558), .Z(n559) );
  NAND2_X1 U624 ( .A1(G125), .A2(n905), .ZN(n561) );
  NAND2_X1 U625 ( .A1(G113), .A2(n906), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G90), .A2(n673), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G77), .A2(n674), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT9), .B(n565), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G52), .A2(n668), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G64), .A2(n669), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT66), .B(n568), .Z(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(G301) );
  INV_X1 U636 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U637 ( .A(G2451), .B(G2446), .ZN(n580) );
  XOR2_X1 U638 ( .A(G2430), .B(KEYINPUT110), .Z(n572) );
  XNOR2_X1 U639 ( .A(G2454), .B(G2435), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n572), .B(n571), .ZN(n576) );
  XOR2_X1 U641 ( .A(G2438), .B(KEYINPUT109), .Z(n574) );
  XNOR2_X1 U642 ( .A(G1348), .B(G1341), .ZN(n573) );
  XNOR2_X1 U643 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U644 ( .A(n576), .B(n575), .Z(n578) );
  XNOR2_X1 U645 ( .A(G2443), .B(G2427), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n581) );
  AND2_X1 U648 ( .A1(n581), .A2(G14), .ZN(G401) );
  INV_X1 U649 ( .A(G57), .ZN(G237) );
  NAND2_X1 U650 ( .A1(G88), .A2(n673), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G75), .A2(n674), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G50), .A2(n668), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G62), .A2(n669), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT83), .B(n586), .Z(n587) );
  NOR2_X1 U657 ( .A1(n588), .A2(n587), .ZN(G166) );
  XOR2_X1 U658 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U659 ( .A1(G94), .A2(G452), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U661 ( .A1(G7), .A2(G661), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U663 ( .A(G223), .ZN(n851) );
  NAND2_X1 U664 ( .A1(n851), .A2(G567), .ZN(n591) );
  XOR2_X1 U665 ( .A(KEYINPUT11), .B(n591), .Z(G234) );
  NAND2_X1 U666 ( .A1(n673), .A2(G81), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G68), .A2(n674), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n595), .B(KEYINPUT13), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G43), .A2(n668), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n669), .A2(G56), .ZN(n598) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n598), .Z(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U676 ( .A(KEYINPUT71), .B(n601), .ZN(n996) );
  INV_X1 U677 ( .A(G860), .ZN(n625) );
  OR2_X1 U678 ( .A1(n996), .A2(n625), .ZN(G153) );
  NAND2_X1 U679 ( .A1(G868), .A2(G171), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G79), .A2(n674), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G54), .A2(n668), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G66), .A2(n669), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n673), .A2(G92), .ZN(n604) );
  XOR2_X1 U685 ( .A(KEYINPUT72), .B(n604), .Z(n605) );
  NOR2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT15), .ZN(n980) );
  INV_X1 U689 ( .A(G868), .ZN(n689) );
  NAND2_X1 U690 ( .A1(n980), .A2(n689), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT73), .ZN(G284) );
  NAND2_X1 U693 ( .A1(n668), .A2(G53), .ZN(n613) );
  XNOR2_X1 U694 ( .A(KEYINPUT69), .B(n613), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n669), .A2(G65), .ZN(n614) );
  XOR2_X1 U696 ( .A(KEYINPUT68), .B(n614), .Z(n615) );
  NOR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U698 ( .A(KEYINPUT70), .B(n617), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G91), .A2(n673), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G78), .A2(n674), .ZN(n618) );
  AND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(G299) );
  NOR2_X1 U703 ( .A1(G286), .A2(n689), .ZN(n622) );
  XOR2_X1 U704 ( .A(KEYINPUT75), .B(n622), .Z(n624) );
  NOR2_X1 U705 ( .A1(G868), .A2(G299), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n624), .A2(n623), .ZN(G297) );
  NAND2_X1 U707 ( .A1(n625), .A2(G559), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n626), .A2(n980), .ZN(n627) );
  XNOR2_X1 U709 ( .A(n627), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U710 ( .A1(n980), .A2(G868), .ZN(n628) );
  NOR2_X1 U711 ( .A1(G559), .A2(n628), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT76), .ZN(n631) );
  NOR2_X1 U713 ( .A1(n996), .A2(G868), .ZN(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(G282) );
  XOR2_X1 U715 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n633) );
  NAND2_X1 U716 ( .A1(G123), .A2(n905), .ZN(n632) );
  XNOR2_X1 U717 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n634), .B(KEYINPUT77), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n906), .A2(G111), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G135), .A2(n910), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G99), .A2(n557), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n954) );
  XNOR2_X1 U725 ( .A(n954), .B(G2096), .ZN(n642) );
  INV_X1 U726 ( .A(G2100), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(G156) );
  NAND2_X1 U728 ( .A1(n980), .A2(G559), .ZN(n685) );
  XNOR2_X1 U729 ( .A(n996), .B(n685), .ZN(n643) );
  NOR2_X1 U730 ( .A1(n643), .A2(G860), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G93), .A2(n673), .ZN(n645) );
  NAND2_X1 U732 ( .A1(G80), .A2(n674), .ZN(n644) );
  NAND2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G55), .A2(n668), .ZN(n647) );
  NAND2_X1 U735 ( .A1(G67), .A2(n669), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n647), .A2(n646), .ZN(n648) );
  OR2_X1 U737 ( .A1(n649), .A2(n648), .ZN(n688) );
  XOR2_X1 U738 ( .A(n650), .B(n688), .Z(G145) );
  NAND2_X1 U739 ( .A1(G48), .A2(n668), .ZN(n652) );
  NAND2_X1 U740 ( .A1(G61), .A2(n669), .ZN(n651) );
  NAND2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n673), .A2(G86), .ZN(n653) );
  XOR2_X1 U743 ( .A(KEYINPUT80), .B(n653), .Z(n654) );
  NOR2_X1 U744 ( .A1(n655), .A2(n654), .ZN(n659) );
  XOR2_X1 U745 ( .A(KEYINPUT81), .B(KEYINPUT2), .Z(n657) );
  NAND2_X1 U746 ( .A1(G73), .A2(n674), .ZN(n656) );
  XNOR2_X1 U747 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U748 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U749 ( .A(n660), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U750 ( .A1(G49), .A2(n668), .ZN(n663) );
  NAND2_X1 U751 ( .A1(G87), .A2(n661), .ZN(n662) );
  NAND2_X1 U752 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U753 ( .A1(n669), .A2(n664), .ZN(n667) );
  NAND2_X1 U754 ( .A1(G74), .A2(G651), .ZN(n665) );
  XOR2_X1 U755 ( .A(KEYINPUT79), .B(n665), .Z(n666) );
  NAND2_X1 U756 ( .A1(n667), .A2(n666), .ZN(G288) );
  NAND2_X1 U757 ( .A1(G47), .A2(n668), .ZN(n671) );
  NAND2_X1 U758 ( .A1(G60), .A2(n669), .ZN(n670) );
  NAND2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U760 ( .A(KEYINPUT65), .B(n672), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G85), .A2(n673), .ZN(n676) );
  NAND2_X1 U762 ( .A1(G72), .A2(n674), .ZN(n675) );
  AND2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(G290) );
  XNOR2_X1 U765 ( .A(n688), .B(KEYINPUT19), .ZN(n679) );
  XNOR2_X1 U766 ( .A(G288), .B(n679), .ZN(n680) );
  XNOR2_X1 U767 ( .A(G305), .B(n680), .ZN(n683) );
  XNOR2_X1 U768 ( .A(G166), .B(G290), .ZN(n681) );
  XNOR2_X1 U769 ( .A(n681), .B(G299), .ZN(n682) );
  XNOR2_X1 U770 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n684), .B(n996), .ZN(n876) );
  XNOR2_X1 U772 ( .A(n876), .B(n685), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n686), .A2(G868), .ZN(n687) );
  XNOR2_X1 U774 ( .A(n687), .B(KEYINPUT84), .ZN(n691) );
  NAND2_X1 U775 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n691), .A2(n690), .ZN(G295) );
  NAND2_X1 U777 ( .A1(G2084), .A2(G2078), .ZN(n692) );
  XOR2_X1 U778 ( .A(KEYINPUT20), .B(n692), .Z(n693) );
  NAND2_X1 U779 ( .A1(G2090), .A2(n693), .ZN(n694) );
  XNOR2_X1 U780 ( .A(KEYINPUT21), .B(n694), .ZN(n695) );
  NAND2_X1 U781 ( .A1(n695), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U782 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U783 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n697) );
  NAND2_X1 U784 ( .A1(G132), .A2(G82), .ZN(n696) );
  XNOR2_X1 U785 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U786 ( .A1(n698), .A2(G218), .ZN(n699) );
  XNOR2_X1 U787 ( .A(KEYINPUT86), .B(n699), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n700), .A2(G96), .ZN(n701) );
  XOR2_X1 U789 ( .A(n701), .B(KEYINPUT87), .Z(n856) );
  AND2_X1 U790 ( .A1(n856), .A2(G2106), .ZN(n706) );
  NAND2_X1 U791 ( .A1(G120), .A2(G108), .ZN(n702) );
  NOR2_X1 U792 ( .A1(G237), .A2(n702), .ZN(n703) );
  NAND2_X1 U793 ( .A1(G69), .A2(n703), .ZN(n855) );
  NAND2_X1 U794 ( .A1(G567), .A2(n855), .ZN(n704) );
  XOR2_X1 U795 ( .A(KEYINPUT88), .B(n704), .Z(n705) );
  NOR2_X1 U796 ( .A1(n706), .A2(n705), .ZN(G319) );
  INV_X1 U797 ( .A(G319), .ZN(n708) );
  NAND2_X1 U798 ( .A1(G483), .A2(G661), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n854) );
  NAND2_X1 U800 ( .A1(n854), .A2(G36), .ZN(G176) );
  INV_X1 U801 ( .A(G166), .ZN(G303) );
  INV_X1 U802 ( .A(n814), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n709), .A2(n815), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n717), .A2(G1996), .ZN(n711) );
  XNOR2_X1 U805 ( .A(n711), .B(KEYINPUT26), .ZN(n713) );
  INV_X1 U806 ( .A(n717), .ZN(n753) );
  NAND2_X1 U807 ( .A1(n753), .A2(G1341), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U809 ( .A1(n716), .A2(n980), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n980), .ZN(n721) );
  NOR2_X1 U811 ( .A1(G2067), .A2(n753), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n717), .A2(G1348), .ZN(n718) );
  NOR2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  INV_X1 U815 ( .A(G299), .ZN(n987) );
  NAND2_X1 U816 ( .A1(G2072), .A2(n717), .ZN(n723) );
  XNOR2_X1 U817 ( .A(n723), .B(KEYINPUT27), .ZN(n725) );
  AND2_X1 U818 ( .A1(n753), .A2(G1956), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n987), .A2(n727), .ZN(n726) );
  NOR2_X1 U821 ( .A1(n987), .A2(n727), .ZN(n728) );
  XOR2_X1 U822 ( .A(n728), .B(KEYINPUT28), .Z(n729) );
  XNOR2_X1 U823 ( .A(n730), .B(KEYINPUT29), .ZN(n735) );
  XOR2_X1 U824 ( .A(KEYINPUT25), .B(G2078), .Z(n932) );
  NAND2_X1 U825 ( .A1(n932), .A2(n717), .ZN(n732) );
  NAND2_X1 U826 ( .A1(n753), .A2(G1961), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U828 ( .A(KEYINPUT100), .B(n733), .Z(n743) );
  AND2_X1 U829 ( .A1(G171), .A2(n743), .ZN(n734) );
  NOR2_X1 U830 ( .A1(n735), .A2(n734), .ZN(n749) );
  INV_X1 U831 ( .A(KEYINPUT99), .ZN(n736) );
  NAND2_X1 U832 ( .A1(G8), .A2(n762), .ZN(n739) );
  NAND2_X1 U833 ( .A1(G8), .A2(n738), .ZN(n795) );
  NOR2_X1 U834 ( .A1(G1966), .A2(n795), .ZN(n765) );
  NOR2_X1 U835 ( .A1(n739), .A2(n765), .ZN(n740) );
  XNOR2_X1 U836 ( .A(n740), .B(KEYINPUT30), .ZN(n742) );
  INV_X1 U837 ( .A(G168), .ZN(n741) );
  NOR2_X1 U838 ( .A1(G171), .A2(n743), .ZN(n744) );
  XNOR2_X1 U839 ( .A(KEYINPUT31), .B(n746), .ZN(n747) );
  XNOR2_X1 U840 ( .A(n747), .B(KEYINPUT102), .ZN(n748) );
  NOR2_X1 U841 ( .A1(n749), .A2(n748), .ZN(n751) );
  XNOR2_X1 U842 ( .A(n751), .B(n750), .ZN(n764) );
  INV_X1 U843 ( .A(n764), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n752), .A2(G286), .ZN(n760) );
  INV_X1 U845 ( .A(G8), .ZN(n758) );
  NOR2_X1 U846 ( .A1(n753), .A2(G2090), .ZN(n755) );
  NOR2_X1 U847 ( .A1(G1971), .A2(n795), .ZN(n754) );
  NOR2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U849 ( .A1(n756), .A2(G303), .ZN(n757) );
  OR2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  INV_X1 U852 ( .A(n762), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n763), .A2(G8), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n772) );
  NOR2_X1 U858 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n986) );
  INV_X1 U860 ( .A(n795), .ZN(n778) );
  NAND2_X1 U861 ( .A1(n772), .A2(n778), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n773), .A2(KEYINPUT33), .ZN(n776) );
  AND2_X1 U863 ( .A1(n986), .A2(n776), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n783) );
  INV_X1 U865 ( .A(n776), .ZN(n781) );
  INV_X1 U866 ( .A(KEYINPUT33), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n979) );
  AND2_X1 U868 ( .A1(n777), .A2(n979), .ZN(n779) );
  AND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  OR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(n784), .ZN(n786) );
  XOR2_X1 U873 ( .A(G1981), .B(G305), .Z(n988) );
  NAND2_X1 U874 ( .A1(G8), .A2(G166), .ZN(n787) );
  XNOR2_X1 U875 ( .A(n789), .B(KEYINPUT107), .ZN(n790) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n793) );
  XNOR2_X1 U877 ( .A(KEYINPUT97), .B(KEYINPUT24), .ZN(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(KEYINPUT98), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n793), .B(n792), .ZN(n794) );
  NOR2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n838) );
  NAND2_X1 U881 ( .A1(n557), .A2(G105), .ZN(n797) );
  XNOR2_X1 U882 ( .A(KEYINPUT38), .B(KEYINPUT94), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n797), .B(n796), .ZN(n804) );
  NAND2_X1 U884 ( .A1(G129), .A2(n905), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G117), .A2(n906), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U887 ( .A1(G141), .A2(n910), .ZN(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT95), .B(n800), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n894) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n894), .ZN(n960) );
  NAND2_X1 U892 ( .A1(G119), .A2(n905), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G107), .A2(n906), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U895 ( .A1(G131), .A2(n910), .ZN(n807) );
  XNOR2_X1 U896 ( .A(KEYINPUT93), .B(n807), .ZN(n808) );
  NOR2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U898 ( .A1(n557), .A2(G95), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n892) );
  NAND2_X1 U900 ( .A1(G1991), .A2(n892), .ZN(n813) );
  NAND2_X1 U901 ( .A1(G1996), .A2(n894), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n955) );
  NOR2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n841) );
  NAND2_X1 U904 ( .A1(n955), .A2(n841), .ZN(n816) );
  XOR2_X1 U905 ( .A(KEYINPUT96), .B(n816), .Z(n842) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n892), .ZN(n956) );
  NOR2_X1 U908 ( .A1(n817), .A2(n956), .ZN(n818) );
  NOR2_X1 U909 ( .A1(n842), .A2(n818), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n819), .B(KEYINPUT108), .ZN(n820) );
  NOR2_X1 U911 ( .A1(n960), .A2(n820), .ZN(n821) );
  XNOR2_X1 U912 ( .A(KEYINPUT39), .B(n821), .ZN(n833) );
  XNOR2_X1 U913 ( .A(G2067), .B(KEYINPUT37), .ZN(n834) );
  NAND2_X1 U914 ( .A1(G128), .A2(n905), .ZN(n823) );
  NAND2_X1 U915 ( .A1(G116), .A2(n906), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U917 ( .A(KEYINPUT35), .B(n824), .Z(n831) );
  XNOR2_X1 U918 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT34), .ZN(n829) );
  NAND2_X1 U920 ( .A1(G140), .A2(n910), .ZN(n827) );
  NAND2_X1 U921 ( .A1(G104), .A2(n557), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U923 ( .A(n829), .B(n828), .Z(n830) );
  NOR2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U925 ( .A(KEYINPUT36), .B(n832), .ZN(n918) );
  NOR2_X1 U926 ( .A1(n834), .A2(n918), .ZN(n968) );
  NAND2_X1 U927 ( .A1(n841), .A2(n968), .ZN(n843) );
  NAND2_X1 U928 ( .A1(n833), .A2(n843), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n834), .A2(n918), .ZN(n965) );
  NAND2_X1 U930 ( .A1(n835), .A2(n965), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n836), .A2(n841), .ZN(n848) );
  INV_X1 U932 ( .A(n848), .ZN(n837) );
  XNOR2_X1 U933 ( .A(KEYINPUT90), .B(G1986), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n840), .B(G290), .ZN(n1000) );
  AND2_X1 U935 ( .A1(n1000), .A2(n841), .ZN(n846) );
  INV_X1 U936 ( .A(n842), .ZN(n844) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n845) );
  OR2_X1 U938 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U939 ( .A(n850), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n851), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U942 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U944 ( .A1(n854), .A2(n853), .ZN(G188) );
  XNOR2_X1 U945 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U947 ( .A(G132), .ZN(G219) );
  INV_X1 U948 ( .A(G120), .ZN(G236) );
  INV_X1 U949 ( .A(G96), .ZN(G221) );
  INV_X1 U950 ( .A(G82), .ZN(G220) );
  NOR2_X1 U951 ( .A1(n856), .A2(n855), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XOR2_X1 U953 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(G2072), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U960 ( .A(G2084), .B(G2078), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(G227) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1981), .Z(n866) );
  XNOR2_X1 U963 ( .A(G1966), .B(G1956), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U965 ( .A(n867), .B(KEYINPUT111), .Z(n869) );
  XNOR2_X1 U966 ( .A(G1991), .B(G1996), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U968 ( .A(G1976), .B(G1961), .Z(n871) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1971), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U971 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U972 ( .A(KEYINPUT112), .B(G2474), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(G229) );
  XOR2_X1 U974 ( .A(n876), .B(n980), .Z(n878) );
  XNOR2_X1 U975 ( .A(G286), .B(G171), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n879) );
  NOR2_X1 U977 ( .A1(G37), .A2(n879), .ZN(G397) );
  NAND2_X1 U978 ( .A1(n905), .A2(G124), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n880), .B(KEYINPUT44), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G112), .A2(n906), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U982 ( .A1(G136), .A2(n910), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G100), .A2(n557), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(G162) );
  XOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n888) );
  XNOR2_X1 U987 ( .A(KEYINPUT115), .B(KEYINPUT114), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n889), .B(G162), .Z(n891) );
  XNOR2_X1 U990 ( .A(G164), .B(G160), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n904) );
  NAND2_X1 U994 ( .A1(G130), .A2(n905), .ZN(n897) );
  NAND2_X1 U995 ( .A1(G118), .A2(n906), .ZN(n896) );
  NAND2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n902) );
  NAND2_X1 U997 ( .A1(G142), .A2(n910), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G106), .A2(n557), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(KEYINPUT45), .B(n900), .Z(n901) );
  NOR2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(n904), .B(n903), .Z(n917) );
  NAND2_X1 U1003 ( .A1(G127), .A2(n905), .ZN(n908) );
  NAND2_X1 U1004 ( .A1(G115), .A2(n906), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n909), .B(KEYINPUT47), .ZN(n912) );
  NAND2_X1 U1007 ( .A1(G139), .A2(n910), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n915) );
  NAND2_X1 U1009 ( .A1(G103), .A2(n557), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT113), .B(n913), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n949) );
  XNOR2_X1 U1012 ( .A(n949), .B(n954), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n920), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT116), .B(n921), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n923), .ZN(n924) );
  AND2_X1 U1020 ( .A1(G319), .A2(n924), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G397), .A2(G395), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1025 ( .A(G29), .B(KEYINPUT123), .ZN(n948) );
  XOR2_X1 U1026 ( .A(G2090), .B(G35), .Z(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n927) );
  XNOR2_X1 U1028 ( .A(G34), .B(n927), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(n928), .B(G2084), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n945) );
  XOR2_X1 U1031 ( .A(G1991), .B(G25), .Z(n931) );
  NAND2_X1 U1032 ( .A1(n931), .A2(G28), .ZN(n941) );
  XNOR2_X1 U1033 ( .A(G1996), .B(G32), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(n932), .B(G27), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(KEYINPUT120), .B(n935), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G2067), .B(G26), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(G33), .B(G2072), .ZN(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1042 ( .A(KEYINPUT121), .B(n942), .Z(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT53), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(KEYINPUT55), .B(n946), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n977) );
  XOR2_X1 U1047 ( .A(G2072), .B(n949), .Z(n951) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1050 ( .A(KEYINPUT50), .B(n952), .Z(n971) );
  XOR2_X1 U1051 ( .A(G2084), .B(G160), .Z(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1055 ( .A(G2090), .B(G162), .Z(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT118), .B(n961), .Z(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT51), .B(n962), .Z(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT119), .B(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n972), .B(KEYINPUT52), .ZN(n974) );
  INV_X1 U1065 ( .A(KEYINPUT55), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(G29), .A2(n975), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n1030) );
  XOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .Z(n1002) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1348), .B(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G171), .B(G1961), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n994) );
  XNOR2_X1 U1077 ( .A(n987), .B(G1956), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G168), .B(G1966), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(n990), .B(KEYINPUT57), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n998) );
  XOR2_X1 U1083 ( .A(G1341), .B(KEYINPUT124), .Z(n995) );
  XNOR2_X1 U1084 ( .A(n996), .B(n995), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1027) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(n1003), .B(G4), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G6), .B(G1981), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(KEYINPUT125), .B(G1956), .Z(n1008) );
  XNOR2_X1 U1095 ( .A(G20), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1011), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(n1012), .B(KEYINPUT126), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G21), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1103 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G23), .B(G1976), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1024), .Z(n1025) );
  NOR2_X1 U1111 ( .A1(G16), .A2(n1025), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(G11), .ZN(n1032) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

