//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  AND3_X1   g0031(.A1(new_n217), .A2(new_n230), .A3(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n205), .A2(G20), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT68), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(new_n213), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n252), .B1(new_n258), .B2(G50), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n201), .A2(new_n206), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n206), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n263), .A2(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n259), .B1(new_n269), .B2(new_n256), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  AND2_X1   g0072(.A1(G1), .A2(G13), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(new_n274), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n276), .ZN(new_n280));
  INV_X1    g0080(.A(G226), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G222), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G223), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(G77), .B2(new_n283), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n279), .B1(new_n288), .B2(KEYINPUT66), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT71), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(G200), .B1(new_n293), .B2(KEYINPUT10), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(G190), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n271), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G232), .A2(G1698), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n285), .A2(G238), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n283), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G107), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G107), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n301), .B1(new_n306), .B2(new_n283), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT70), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n279), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n278), .B1(new_n280), .B2(new_n219), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G20), .A2(G77), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT15), .B(G87), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n317), .B1(new_n318), .B2(new_n264), .C1(new_n267), .C2(new_n263), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n255), .A2(new_n213), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n258), .A2(G77), .ZN(new_n322));
  INV_X1    g0122(.A(new_n251), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n202), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n312), .B1(new_n309), .B2(new_n310), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n314), .A2(G200), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n326), .B2(G190), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n316), .A2(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n297), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n271), .A2(new_n294), .A3(new_n333), .A4(new_n295), .ZN(new_n334));
  INV_X1    g0134(.A(new_n270), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n327), .B2(new_n291), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(G169), .B2(new_n291), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n298), .A2(new_n332), .A3(new_n334), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n226), .A2(G20), .ZN(new_n339));
  INV_X1    g0139(.A(G50), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(new_n264), .B2(new_n202), .C1(new_n267), .C2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT11), .A3(new_n320), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n250), .A2(KEYINPUT12), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n342), .B1(KEYINPUT12), .B2(new_n323), .C1(new_n339), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT11), .B1(new_n341), .B2(new_n320), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n258), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n226), .B1(new_n347), .B2(KEYINPUT12), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n281), .A2(new_n285), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n225), .A2(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n283), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT72), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(KEYINPUT72), .A3(new_n354), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n278), .B1(new_n280), .B2(new_n227), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT13), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n279), .B1(new_n355), .B2(new_n356), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n359), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  INV_X1    g0165(.A(new_n361), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n362), .A2(G179), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n369));
  AOI211_X1 g0169(.A(KEYINPUT13), .B(new_n361), .C1(new_n363), .C2(new_n359), .ZN(new_n370));
  OAI21_X1  g0170(.A(G169), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n368), .B1(new_n371), .B2(KEYINPUT14), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT14), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n362), .A2(new_n367), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(G169), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n350), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n350), .B1(new_n374), .B2(G200), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n374), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n338), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n263), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n251), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n258), .B2(new_n383), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n358), .A2(new_n272), .A3(new_n276), .ZN(new_n386));
  INV_X1    g0186(.A(new_n280), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n386), .B1(G232), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G33), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G223), .A2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n281), .B2(G1698), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n393), .A2(new_n395), .B1(G33), .B2(G87), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n388), .B1(new_n279), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n388), .B(new_n378), .C1(new_n279), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT77), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT3), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT77), .A3(G33), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT74), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n405), .A2(KEYINPUT74), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n389), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n411), .B2(KEYINPUT76), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(new_n389), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n402), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n405), .A2(G33), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n390), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n206), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(G68), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(G58), .B(G68), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(G20), .B1(G159), .B2(new_n266), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT16), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n405), .A2(KEYINPUT74), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(G33), .ZN(new_n426));
  AOI21_X1  g0226(.A(G20), .B1(new_n426), .B2(new_n390), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT7), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI211_X1 g0229(.A(G20), .B(new_n416), .C1(new_n426), .C2(new_n390), .ZN(new_n430));
  OAI211_X1 g0230(.A(KEYINPUT16), .B(new_n422), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n320), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n385), .B(new_n401), .C1(new_n423), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n433), .B(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n385), .B1(new_n423), .B2(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n397), .A2(G169), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n388), .B(G179), .C1(new_n279), .C2(new_n396), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT18), .B1(new_n436), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(KEYINPUT78), .ZN(new_n442));
  INV_X1    g0242(.A(new_n385), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT76), .B1(new_n392), .B2(G33), .ZN(new_n444));
  INV_X1    g0244(.A(new_n407), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n414), .ZN(new_n446));
  INV_X1    g0246(.A(new_n402), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n419), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n422), .B1(new_n448), .B2(new_n226), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT16), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n431), .A2(new_n320), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n443), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n439), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT18), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT78), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n435), .B1(new_n442), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n376), .A2(new_n379), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT73), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n382), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  OR3_X1    g0261(.A1(new_n251), .A2(KEYINPUT25), .A3(G107), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT25), .B1(new_n251), .B2(G107), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n256), .B(new_n251), .C1(G1), .C2(new_n389), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n462), .B(new_n463), .C1(new_n302), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT85), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n303), .A2(new_n305), .A3(G20), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n468), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT83), .B1(new_n468), .B2(KEYINPUT23), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n206), .A2(G87), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT22), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n426), .A2(new_n474), .A3(new_n390), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n418), .B2(new_n472), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G20), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n475), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT24), .B1(new_n471), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n475), .A2(new_n476), .A3(new_n480), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n468), .A2(KEYINPUT23), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n468), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n256), .B1(new_n482), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n467), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI211_X1 g0293(.A(KEYINPUT84), .B(new_n256), .C1(new_n482), .C2(new_n490), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(G41), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g0299(.A(G45), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G1), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n275), .A2(new_n497), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n497), .A3(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n279), .ZN(new_n504));
  INV_X1    g0304(.A(G264), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(G257), .A2(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n426), .A2(new_n390), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT86), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n426), .A2(new_n511), .A3(new_n390), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n426), .A2(G250), .A3(new_n285), .A4(new_n390), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n510), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(new_n516), .A3(new_n358), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n515), .B2(new_n358), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n507), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n506), .B1(new_n515), .B2(new_n358), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n519), .A2(G190), .B1(G200), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n495), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n519), .A2(G169), .B1(G179), .B2(new_n520), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n495), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT88), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n491), .A2(new_n492), .ZN(new_n526));
  INV_X1    g0326(.A(new_n494), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(new_n467), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(G169), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n520), .A2(G179), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n495), .A2(new_n521), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT88), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n537), .A2(new_n219), .A3(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n283), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n283), .B2(G250), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n536), .B(new_n539), .C1(new_n540), .C2(new_n285), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT4), .B1(new_n393), .B2(G244), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n358), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n503), .A2(G257), .A3(new_n279), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n502), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n315), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n543), .A2(new_n327), .A3(new_n502), .A4(new_n544), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n306), .B1(new_n415), .B2(new_n419), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n302), .A2(KEYINPUT6), .A3(G97), .ZN(new_n549));
  INV_X1    g0349(.A(G97), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n302), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n553), .B2(KEYINPUT6), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n256), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n464), .A2(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n251), .A2(new_n550), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n557), .A2(KEYINPUT79), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT79), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n546), .B(new_n547), .C1(new_n556), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n545), .A2(G200), .ZN(new_n563));
  INV_X1    g0363(.A(new_n306), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n555), .B1(new_n448), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n320), .ZN(new_n566));
  INV_X1    g0366(.A(new_n561), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n543), .A2(G190), .A3(new_n502), .A4(new_n544), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n563), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n323), .A2(new_n318), .ZN(new_n570));
  INV_X1    g0370(.A(new_n464), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n318), .B(KEYINPUT81), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n303), .A2(new_n305), .A3(new_n220), .A4(new_n550), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n354), .B2(new_n206), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n206), .A2(G33), .A3(G97), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n574), .A2(new_n576), .B1(new_n577), .B2(new_n575), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n426), .A2(new_n206), .A3(G68), .A4(new_n390), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n570), .B(new_n573), .C1(new_n580), .C2(new_n256), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n358), .A2(new_n221), .A3(new_n501), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n279), .A2(G274), .A3(new_n501), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT80), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n275), .A2(KEYINPUT80), .A3(new_n501), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G238), .A2(G1698), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n219), .B2(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(new_n426), .A3(new_n390), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n590), .A2(new_n478), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n587), .B(new_n327), .C1(new_n591), .C2(new_n279), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n279), .B(G250), .C1(G1), .C2(new_n500), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n275), .A2(KEYINPUT80), .A3(new_n501), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT80), .B1(new_n275), .B2(new_n501), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n279), .B1(new_n590), .B2(new_n478), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n315), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n581), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n256), .B1(new_n578), .B2(new_n579), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n464), .A2(new_n220), .ZN(new_n601));
  INV_X1    g0401(.A(new_n570), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n587), .B(G190), .C1(new_n591), .C2(new_n279), .ZN(new_n604));
  OAI21_X1  g0404(.A(G200), .B1(new_n596), .B2(new_n597), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n562), .A2(new_n569), .A3(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n536), .B(new_n206), .C1(G33), .C2(new_n550), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n609), .B(new_n320), .C1(new_n206), .C2(G116), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT20), .ZN(new_n611));
  INV_X1    g0411(.A(G116), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n323), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n464), .B2(new_n612), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G257), .A2(G1698), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n505), .B2(G1698), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n426), .A3(new_n390), .ZN(new_n618));
  XOR2_X1   g0418(.A(KEYINPUT82), .B(G303), .Z(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n418), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n279), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G270), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n502), .B1(new_n504), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n615), .A2(KEYINPUT21), .A3(G169), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(G190), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n611), .A2(new_n614), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n628), .C1(new_n398), .C2(new_n624), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT21), .ZN(new_n630));
  OAI21_X1  g0430(.A(G169), .B1(new_n611), .B2(new_n614), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n624), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n621), .A2(new_n623), .A3(new_n327), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n626), .A2(new_n629), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n608), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n461), .A2(new_n525), .A3(new_n535), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT89), .Z(G372));
  OAI21_X1  g0438(.A(new_n455), .B1(new_n453), .B2(new_n454), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n440), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n372), .A2(new_n375), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n328), .A2(new_n316), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(new_n350), .B1(new_n379), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n435), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT91), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n298), .A2(new_n334), .ZN(new_n647));
  OAI211_X1 g0447(.A(KEYINPUT91), .B(new_n640), .C1(new_n643), .C2(new_n435), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(new_n337), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n626), .A2(new_n632), .A3(new_n634), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n495), .B2(new_n523), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n608), .A3(new_n533), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n599), .B(KEYINPUT90), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n599), .A2(new_n606), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n562), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n546), .A2(new_n547), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n566), .A2(new_n567), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n607), .A3(KEYINPUT26), .A4(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n654), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n461), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n650), .A2(new_n663), .ZN(G369));
  NAND2_X1  g0464(.A1(new_n250), .A2(new_n206), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n528), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n525), .A2(new_n535), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT92), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT92), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n525), .A2(new_n675), .A3(new_n535), .A4(new_n672), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n651), .A2(new_n671), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n670), .B(KEYINPUT93), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n524), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT94), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n674), .A2(new_n676), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n532), .A2(new_n670), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n635), .B1(new_n628), .B2(new_n670), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n615), .A2(new_n671), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n651), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n685), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n209), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n574), .A2(G116), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n698), .A2(new_n205), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n698), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n701), .A2(KEYINPUT95), .B1(new_n215), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(KEYINPUT95), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  INV_X1    g0505(.A(G330), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n596), .A2(new_n597), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(new_n543), .A3(new_n544), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n520), .A4(new_n633), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n633), .A2(new_n708), .A3(new_n543), .A4(new_n544), .ZN(new_n712));
  INV_X1    g0512(.A(new_n520), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT30), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR4_X1   g0514(.A1(new_n520), .A2(new_n708), .A3(G179), .A4(new_n624), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n711), .A2(new_n714), .B1(new_n545), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n671), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n714), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n545), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n719), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n707), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n716), .A2(new_n707), .A3(new_n679), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n525), .A2(new_n636), .A3(new_n535), .A4(new_n679), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n706), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n662), .A2(new_n679), .ZN(new_n727));
  XNOR2_X1  g0527(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n671), .B1(new_n653), .B2(new_n661), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(KEYINPUT29), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n705), .B1(new_n731), .B2(G1), .ZN(G364));
  NOR2_X1   g0532(.A1(new_n249), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n205), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n698), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n694), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G330), .B2(new_n692), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n736), .B(KEYINPUT98), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n213), .B1(G20), .B2(new_n315), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n327), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n206), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G159), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n283), .B1(new_n202), .B2(new_n745), .C1(new_n749), .C2(KEYINPUT32), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n206), .A2(new_n378), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n398), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n220), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n743), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n744), .A2(new_n752), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n224), .B1(new_n756), .B2(new_n302), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n750), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n378), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n749), .A2(KEYINPUT32), .B1(new_n760), .B2(G50), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n206), .B1(new_n746), .B2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n550), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n759), .A2(G190), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(G68), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n758), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G322), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n418), .B1(new_n755), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(G326), .B2(new_n760), .ZN(new_n769));
  INV_X1    g0569(.A(new_n756), .ZN(new_n770));
  INV_X1    g0570(.A(new_n745), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G283), .A2(new_n770), .B1(new_n771), .B2(G311), .ZN(new_n772));
  INV_X1    g0572(.A(new_n753), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G303), .A2(new_n773), .B1(new_n748), .B2(G329), .ZN(new_n774));
  INV_X1    g0574(.A(new_n762), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n775), .A2(G294), .B1(new_n764), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n769), .A2(new_n772), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n742), .B1(new_n766), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n741), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n697), .A2(new_n393), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n216), .A2(new_n500), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n244), .C2(new_n500), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n697), .A2(new_n418), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n787), .A2(G355), .B1(new_n612), .B2(new_n697), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n740), .B(new_n779), .C1(new_n783), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n782), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n692), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n738), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n642), .A2(new_n670), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n329), .A2(new_n331), .B1(new_n330), .B2(new_n671), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n642), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n662), .B2(new_n679), .ZN(new_n799));
  INV_X1    g0599(.A(new_n679), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n800), .B(new_n797), .C1(new_n653), .C2(new_n661), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n726), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n736), .B1(new_n726), .B2(new_n802), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n755), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT99), .B(G143), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n808), .A2(new_n809), .B1(new_n771), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(new_n760), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  INV_X1    g0612(.A(new_n764), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n810), .B1(new_n811), .B2(new_n812), .C1(new_n265), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT34), .ZN(new_n815));
  INV_X1    g0615(.A(new_n393), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n756), .A2(new_n226), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G132), .B2(new_n748), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n340), .B2(new_n753), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n816), .B(new_n819), .C1(G58), .C2(new_n775), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n283), .B(new_n763), .C1(G107), .C2(new_n773), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n756), .A2(new_n220), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G311), .B2(new_n748), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G294), .A2(new_n808), .B1(new_n771), .B2(G116), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G283), .A2(new_n764), .B1(new_n760), .B2(G303), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n742), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n741), .A2(new_n780), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n740), .B(new_n828), .C1(new_n202), .C2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n798), .B2(new_n781), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n807), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  OR2_X1    g0633(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n834), .A2(G116), .A3(new_n214), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT36), .Z(new_n837));
  OAI211_X1 g0637(.A(new_n216), .B(G77), .C1(new_n224), .C2(new_n226), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n340), .A2(G68), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n205), .B(G13), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n641), .A2(new_n350), .A3(new_n671), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n350), .A2(new_n671), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n376), .A2(new_n379), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n795), .B(KEYINPUT101), .Z(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n801), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n429), .A2(new_n430), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n848), .B2(new_n422), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n385), .B1(new_n849), .B2(new_n432), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n669), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n439), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(new_n433), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT102), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n453), .B2(new_n454), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n436), .A2(KEYINPUT102), .A3(new_n439), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n433), .B(new_n859), .C1(new_n453), .C2(new_n668), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n854), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT38), .B(new_n861), .C1(new_n458), .C2(new_n851), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n442), .A2(new_n457), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n433), .B(KEYINPUT17), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n851), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n854), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n860), .B1(new_n857), .B2(new_n856), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n863), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n847), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n640), .A2(new_n669), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT103), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  INV_X1    g0674(.A(new_n872), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n870), .A2(new_n862), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n847), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n641), .A2(new_n350), .A3(new_n670), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n433), .B1(new_n453), .B2(new_n454), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT105), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n436), .A2(new_n669), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT105), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n433), .B(new_n884), .C1(new_n453), .C2(new_n454), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n868), .B1(new_n886), .B2(KEYINPUT37), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n865), .B2(new_n640), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n880), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n890), .A3(new_n862), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n870), .B2(new_n862), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n879), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n873), .A2(new_n877), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n649), .A2(new_n337), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n461), .A2(new_n730), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT106), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT106), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n461), .A2(new_n730), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n896), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n895), .B(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n903));
  OR3_X1    g0703(.A1(new_n718), .A2(new_n721), .A3(new_n707), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n707), .C1(new_n718), .C2(new_n721), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n903), .A2(new_n725), .A3(new_n904), .A4(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n845), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n797), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n453), .A2(new_n455), .A3(new_n454), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT78), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n639), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n865), .B1(new_n912), .B2(new_n456), .ZN(new_n913));
  INV_X1    g0713(.A(new_n851), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n915), .B2(new_n861), .ZN(new_n916));
  INV_X1    g0716(.A(new_n862), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n907), .B(new_n909), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n907), .A2(new_n909), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n889), .B2(new_n862), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n918), .A2(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n922), .A2(new_n461), .A3(new_n907), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n461), .B2(new_n907), .ZN(new_n924));
  OR3_X1    g0724(.A1(new_n923), .A2(new_n924), .A3(new_n706), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n902), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n205), .B2(new_n733), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n902), .A2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n841), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT108), .Z(G367));
  INV_X1    g0730(.A(new_n569), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n659), .B2(new_n800), .ZN(new_n932));
  INV_X1    g0732(.A(new_n562), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n679), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(KEYINPUT42), .B2(new_n680), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n681), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n934), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT42), .B1(new_n678), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n935), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT43), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n603), .A2(new_n670), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT109), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n656), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n654), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n941), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n942), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n695), .ZN(new_n950));
  INV_X1    g0750(.A(new_n936), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n949), .B(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n954));
  XOR2_X1   g0754(.A(new_n698), .B(new_n954), .Z(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT45), .B1(new_n685), .B2(new_n951), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n678), .A2(new_n683), .A3(new_n680), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n683), .B1(new_n678), .B2(new_n680), .ZN(new_n959));
  OAI211_X1 g0759(.A(KEYINPUT45), .B(new_n951), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n682), .A2(new_n684), .A3(new_n936), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n682), .A2(new_n965), .A3(new_n684), .A4(new_n936), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n950), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n960), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n972), .A2(new_n695), .A3(new_n964), .A4(new_n966), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n689), .A2(new_n677), .ZN(new_n974));
  INV_X1    g0774(.A(new_n678), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n694), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n693), .B(new_n678), .C1(new_n689), .C2(new_n677), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(new_n731), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n968), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n956), .B1(new_n980), .B2(new_n731), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n953), .B1(new_n981), .B2(new_n735), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n946), .A2(new_n782), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n784), .A2(new_n240), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n783), .C1(new_n209), .C2(new_n318), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n739), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT111), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n753), .A2(new_n612), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT46), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT112), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n756), .A2(new_n550), .ZN(new_n991));
  INV_X1    g0791(.A(G283), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n745), .A2(new_n992), .B1(new_n747), .B2(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n991), .B(new_n994), .C1(new_n619), .C2(new_n808), .ZN(new_n995));
  INV_X1    g0795(.A(G294), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n988), .A2(KEYINPUT46), .B1(new_n996), .B2(new_n813), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G311), .B2(new_n760), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n393), .B1(new_n306), .B2(new_n775), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n990), .A2(new_n995), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n762), .A2(new_n226), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n418), .B(new_n1001), .C1(G50), .C2(new_n771), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G58), .A2(new_n773), .B1(new_n748), .B2(G137), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n756), .A2(new_n202), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G150), .B2(new_n808), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n760), .A2(new_n809), .B1(new_n764), .B2(G159), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1000), .A2(KEYINPUT47), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT47), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n742), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n987), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n983), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT113), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n982), .A2(new_n1013), .ZN(G387));
  INV_X1    g0814(.A(KEYINPUT116), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n979), .B2(new_n702), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n978), .A2(new_n731), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(KEYINPUT116), .A3(new_n698), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(new_n731), .C2(new_n978), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n978), .A2(new_n735), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n784), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n237), .B2(G45), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n700), .C1(G68), .C2(G77), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(KEYINPUT114), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n263), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1026));
  OAI21_X1  g0826(.A(KEYINPUT50), .B1(new_n263), .B2(G50), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT114), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1027), .C1(new_n1023), .C2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1022), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n787), .A2(new_n700), .B1(new_n302), .B2(new_n697), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n740), .B1(new_n1032), .B2(new_n783), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n572), .A2(new_n775), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G68), .A2(new_n771), .B1(new_n748), .B2(G150), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n340), .C2(new_n755), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n991), .B1(G77), .B2(new_n773), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n383), .A2(new_n764), .B1(G159), .B2(new_n760), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n393), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n753), .A2(new_n996), .B1(new_n762), .B2(new_n992), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n808), .A2(G317), .B1(new_n771), .B2(new_n619), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n764), .A2(G311), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n767), .C2(new_n811), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT49), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT115), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n748), .A2(G326), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n816), .C1(new_n612), .C2(new_n756), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1048), .B2(KEYINPUT115), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1040), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1033), .B1(new_n742), .B2(new_n1053), .C1(new_n689), .C2(new_n791), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1020), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1019), .A2(new_n1055), .ZN(G393));
  NAND3_X1  g0856(.A1(new_n968), .A2(new_n973), .A3(new_n735), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n783), .B1(new_n550), .B2(new_n209), .C1(new_n1021), .C2(new_n247), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n739), .A2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n808), .A2(G159), .B1(G150), .B2(new_n760), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT51), .Z(new_n1061));
  OAI22_X1  g0861(.A1(new_n753), .A2(new_n226), .B1(new_n745), .B2(new_n263), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n823), .B(new_n1062), .C1(new_n748), .C2(new_n809), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n762), .A2(new_n202), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1064), .B(new_n816), .C1(G50), .C2(new_n764), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n771), .A2(G294), .B1(new_n619), .B2(new_n764), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n612), .B2(new_n762), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT118), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n808), .A2(G311), .B1(G317), .B2(new_n760), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n283), .B1(new_n770), .B2(G107), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G283), .A2(new_n773), .B1(new_n748), .B2(G322), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1066), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1059), .B1(new_n1077), .B2(new_n741), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n951), .B2(new_n791), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1057), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n980), .A2(new_n698), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n968), .A2(new_n973), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1017), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(G390));
  AOI21_X1  g0885(.A(new_n740), .B1(new_n263), .B2(new_n829), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT54), .B(G143), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n283), .B1(new_n745), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G132), .A2(new_n808), .B1(new_n748), .B2(G125), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n340), .B2(new_n756), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(G159), .C2(new_n775), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n773), .B2(G150), .ZN(new_n1094));
  INV_X1    g0894(.A(G128), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n813), .A2(new_n812), .B1(new_n811), .B2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n753), .A2(new_n1092), .A3(new_n265), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n755), .A2(new_n612), .B1(new_n747), .B2(new_n996), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n817), .B(new_n1099), .C1(G97), .C2(new_n771), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n564), .A2(new_n813), .B1(new_n811), .B2(new_n992), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1101), .A2(new_n283), .A3(new_n754), .A4(new_n1064), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1091), .A2(new_n1098), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1086), .B1(new_n742), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n892), .A2(new_n893), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n780), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n847), .A2(new_n878), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n891), .B(new_n1108), .C1(new_n876), .C2(new_n890), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n796), .A2(new_n642), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n729), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n795), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n845), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n889), .A2(new_n862), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n878), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n907), .A2(KEYINPUT119), .A3(G330), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1117), .A2(new_n726), .A3(new_n909), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1109), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n907), .A2(G330), .A3(new_n909), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1109), .A2(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1107), .B1(new_n1123), .B2(new_n734), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n845), .B1(new_n726), .B2(new_n798), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1125), .A2(new_n1121), .B1(new_n801), .B2(new_n846), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n907), .A2(G330), .A3(new_n798), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n908), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT120), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1113), .B1(new_n726), .B2(new_n909), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1126), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n461), .A2(G330), .A3(new_n907), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n900), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n899), .B1(new_n461), .B2(new_n730), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n650), .B(new_n1134), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n702), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1123), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1124), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(G378));
  NAND2_X1  g0945(.A1(new_n647), .A2(new_n337), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n335), .A2(new_n668), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1148), .B(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n907), .A2(new_n909), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n919), .B1(new_n876), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n920), .A2(new_n921), .ZN(new_n1154));
  AND4_X1   g0954(.A1(G330), .A2(new_n1151), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1151), .B1(new_n922), .B2(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT122), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n895), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n873), .A2(new_n877), .A3(new_n894), .ZN(new_n1159));
  OAI211_X1 g0959(.A(KEYINPUT122), .B(new_n1159), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n734), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n760), .A2(G125), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n265), .B2(new_n762), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1087), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G128), .A2(new_n808), .B1(new_n773), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n812), .B2(new_n745), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1163), .B(new_n1166), .C1(G132), .C2(new_n764), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n770), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n748), .C2(G124), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n813), .A2(new_n550), .B1(new_n226), .B2(new_n762), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n572), .A2(new_n771), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n393), .A2(G41), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G77), .A2(new_n773), .B1(new_n770), .B2(G58), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G107), .A2(new_n808), .B1(new_n748), .B2(G283), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1174), .B(new_n1179), .C1(G116), .C2(new_n760), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1176), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n340), .C1(G33), .C2(G41), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1173), .A2(new_n1181), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n741), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n735), .B(new_n698), .C1(new_n340), .C2(new_n829), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n1151), .C2(new_n781), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1161), .A2(KEYINPUT123), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT123), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1160), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1153), .A2(G330), .A3(new_n1154), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1151), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n922), .A2(G330), .A3(new_n1151), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1159), .B1(new_n1197), .B2(KEYINPUT122), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n735), .B1(new_n1192), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1191), .B1(new_n1199), .B2(new_n1188), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1190), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1159), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n895), .A2(new_n1196), .A3(new_n1195), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT124), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1137), .B(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1142), .B2(new_n1123), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n702), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1133), .B(new_n1138), .C1(new_n1122), .C2(new_n1119), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1158), .A2(new_n1160), .B1(new_n1210), .B2(new_n1207), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1209), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1201), .A2(new_n1212), .ZN(G375));
  NAND2_X1  g1013(.A1(new_n1133), .A2(new_n735), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n740), .B1(new_n226), .B2(new_n829), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n771), .A2(new_n306), .B1(G294), .B2(new_n760), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n612), .B2(new_n813), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT125), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1004), .A2(new_n283), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n808), .A2(G283), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G97), .A2(new_n773), .B1(new_n748), .B2(G303), .ZN(new_n1221));
  AND4_X1   g1021(.A1(new_n1034), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G159), .A2(new_n773), .B1(new_n771), .B2(G150), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1095), .B2(new_n747), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n755), .A2(new_n812), .B1(new_n756), .B2(new_n224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1224), .A2(new_n816), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n760), .A2(G132), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n340), .B2(new_n762), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n764), .B2(new_n1164), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1218), .A2(new_n1222), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1215), .B1(new_n742), .B2(new_n1230), .C1(new_n845), .C2(new_n781), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1214), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1137), .B(new_n1126), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1142), .A2(new_n955), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(G381));
  NAND3_X1  g1036(.A1(new_n1201), .A2(new_n1144), .A3(new_n1212), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1084), .A2(new_n982), .A3(new_n1013), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1239), .A2(new_n832), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1240));
  OR3_X1    g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(G407));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G343), .C2(new_n1237), .ZN(G409));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(G343), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1208), .B(new_n955), .C1(new_n1192), .C2(new_n1198), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1248), .A2(KEYINPUT126), .A3(new_n955), .A4(new_n1208), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1189), .B1(new_n1250), .B2(new_n735), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1247), .A2(new_n1249), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1144), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1212), .C1(new_n1190), .C2(new_n1200), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1244), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1234), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n698), .A3(new_n1142), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT127), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1234), .B2(new_n1257), .ZN(new_n1261));
  OR3_X1    g1061(.A1(new_n1234), .A2(new_n1260), .A3(new_n1257), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n832), .B1(new_n1263), .B2(new_n1232), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1261), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1259), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(G384), .A3(new_n1233), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1244), .A2(G2897), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1264), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1084), .A2(new_n982), .A3(new_n1013), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1080), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n982), .A2(new_n1013), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n793), .B1(new_n1019), .B2(new_n1055), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1239), .A2(new_n1281), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1277), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1239), .A2(new_n1281), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(G390), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1285), .B2(new_n1238), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1269), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1255), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1288), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1276), .A2(new_n1287), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1255), .A2(new_n1294), .A3(new_n1288), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1255), .B2(new_n1274), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1294), .B1(new_n1255), .B2(new_n1288), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1295), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1293), .B1(new_n1299), .B2(new_n1287), .ZN(G405));
  AOI21_X1  g1100(.A(G378), .B1(new_n1201), .B2(new_n1212), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1254), .ZN(new_n1302));
  OR3_X1    g1102(.A1(new_n1301), .A2(new_n1288), .A3(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1288), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1287), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1287), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(G402));
endmodule


