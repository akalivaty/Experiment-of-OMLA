

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(n668), .ZN(n696) );
  INV_X1 U549 ( .A(n696), .ZN(n702) );
  XOR2_X1 U550 ( .A(KEYINPUT65), .B(n524), .Z(n615) );
  XNOR2_X1 U551 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U552 ( .A1(n544), .A2(n543), .ZN(n546) );
  NOR2_X1 U553 ( .A1(G651), .A2(n629), .ZN(n624) );
  NOR2_X2 U554 ( .A1(G2104), .A2(G2105), .ZN(n512) );
  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n757) );
  NOR2_X2 U556 ( .A1(n663), .A2(n662), .ZN(G164) );
  XOR2_X2 U557 ( .A(KEYINPUT17), .B(n512), .Z(n869) );
  INV_X1 U558 ( .A(KEYINPUT26), .ZN(n669) );
  NOR2_X1 U559 ( .A1(n673), .A2(n969), .ZN(n674) );
  INV_X1 U560 ( .A(KEYINPUT93), .ZN(n713) );
  NAND2_X1 U561 ( .A1(n712), .A2(n711), .ZN(n721) );
  INV_X1 U562 ( .A(KEYINPUT97), .ZN(n730) );
  XNOR2_X1 U563 ( .A(n731), .B(n730), .ZN(n732) );
  INV_X1 U564 ( .A(KEYINPUT13), .ZN(n540) );
  AND2_X2 U565 ( .A1(n517), .A2(G2104), .ZN(n866) );
  XNOR2_X1 U566 ( .A(n541), .B(n540), .ZN(n544) );
  NAND2_X1 U567 ( .A1(n546), .A2(n545), .ZN(n969) );
  NAND2_X1 U568 ( .A1(n869), .A2(G137), .ZN(n515) );
  INV_X1 U569 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U570 ( .A1(G101), .A2(n866), .ZN(n513) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n513), .Z(n514) );
  NAND2_X1 U572 ( .A1(n515), .A2(n514), .ZN(n522) );
  INV_X1 U573 ( .A(G2104), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n516), .A2(n517), .ZN(n861) );
  NAND2_X1 U575 ( .A1(n861), .A2(G113), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n517), .A2(G2104), .ZN(n518) );
  XNOR2_X1 U577 ( .A(n518), .B(KEYINPUT66), .ZN(n580) );
  NAND2_X1 U578 ( .A1(G125), .A2(n580), .ZN(n519) );
  NAND2_X1 U579 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X2 U580 ( .A1(n522), .A2(n521), .ZN(G160) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n629) );
  NAND2_X1 U582 ( .A1(G52), .A2(n624), .ZN(n523) );
  XOR2_X1 U583 ( .A(KEYINPUT68), .B(n523), .Z(n533) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n524) );
  NAND2_X1 U585 ( .A1(G90), .A2(n615), .ZN(n526) );
  XNOR2_X1 U586 ( .A(G651), .B(KEYINPUT67), .ZN(n528) );
  NOR2_X1 U587 ( .A1(n629), .A2(n528), .ZN(n618) );
  NAND2_X1 U588 ( .A1(G77), .A2(n618), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT9), .ZN(n531) );
  NOR2_X1 U591 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X2 U592 ( .A(KEYINPUT1), .B(n529), .Z(n628) );
  NAND2_X1 U593 ( .A1(G64), .A2(n628), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(G171) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U597 ( .A(G132), .ZN(G219) );
  INV_X1 U598 ( .A(G82), .ZN(G220) );
  NAND2_X1 U599 ( .A1(G7), .A2(G661), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U601 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n536) );
  INV_X1 U602 ( .A(G223), .ZN(n817) );
  NAND2_X1 U603 ( .A1(G567), .A2(n817), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G234) );
  NAND2_X1 U605 ( .A1(n615), .A2(G81), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n537), .B(KEYINPUT12), .ZN(n539) );
  NAND2_X1 U607 ( .A1(G68), .A2(n618), .ZN(n538) );
  NAND2_X1 U608 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U609 ( .A1(G56), .A2(n628), .ZN(n542) );
  XOR2_X1 U610 ( .A(KEYINPUT14), .B(n542), .Z(n543) );
  NAND2_X1 U611 ( .A1(n624), .A2(G43), .ZN(n545) );
  INV_X1 U612 ( .A(G860), .ZN(n574) );
  OR2_X1 U613 ( .A1(n969), .A2(n574), .ZN(G153) );
  INV_X1 U614 ( .A(G171), .ZN(G301) );
  NAND2_X1 U615 ( .A1(G868), .A2(G301), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G66), .A2(n628), .ZN(n548) );
  NAND2_X1 U617 ( .A1(G92), .A2(n615), .ZN(n547) );
  NAND2_X1 U618 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U619 ( .A1(G79), .A2(n618), .ZN(n550) );
  NAND2_X1 U620 ( .A1(G54), .A2(n624), .ZN(n549) );
  NAND2_X1 U621 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U622 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U623 ( .A(KEYINPUT15), .B(n553), .Z(n891) );
  INV_X1 U624 ( .A(n891), .ZN(n974) );
  INV_X1 U625 ( .A(G868), .ZN(n639) );
  NAND2_X1 U626 ( .A1(n974), .A2(n639), .ZN(n554) );
  NAND2_X1 U627 ( .A1(n555), .A2(n554), .ZN(G284) );
  NAND2_X1 U628 ( .A1(n615), .A2(G89), .ZN(n556) );
  XNOR2_X1 U629 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U630 ( .A1(G76), .A2(n618), .ZN(n557) );
  NAND2_X1 U631 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U632 ( .A(n559), .B(KEYINPUT5), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G63), .A2(n628), .ZN(n561) );
  NAND2_X1 U634 ( .A1(G51), .A2(n624), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U636 ( .A(KEYINPUT6), .B(n562), .Z(n563) );
  NAND2_X1 U637 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U638 ( .A(n565), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G65), .A2(n628), .ZN(n567) );
  NAND2_X1 U641 ( .A1(G53), .A2(n624), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U643 ( .A1(G91), .A2(n615), .ZN(n569) );
  NAND2_X1 U644 ( .A1(G78), .A2(n618), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U646 ( .A1(n571), .A2(n570), .ZN(n966) );
  INV_X1 U647 ( .A(n966), .ZN(G299) );
  NOR2_X1 U648 ( .A1(G286), .A2(n639), .ZN(n573) );
  NOR2_X1 U649 ( .A1(G868), .A2(G299), .ZN(n572) );
  NOR2_X1 U650 ( .A1(n573), .A2(n572), .ZN(G297) );
  NAND2_X1 U651 ( .A1(n574), .A2(G559), .ZN(n575) );
  NAND2_X1 U652 ( .A1(n575), .A2(n891), .ZN(n576) );
  XNOR2_X1 U653 ( .A(n576), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U654 ( .A1(G868), .A2(n969), .ZN(n579) );
  NAND2_X1 U655 ( .A1(G868), .A2(n891), .ZN(n577) );
  NOR2_X1 U656 ( .A1(G559), .A2(n577), .ZN(n578) );
  NOR2_X1 U657 ( .A1(n579), .A2(n578), .ZN(G282) );
  BUF_X1 U658 ( .A(n580), .Z(n862) );
  NAND2_X1 U659 ( .A1(n862), .A2(G123), .ZN(n581) );
  XNOR2_X1 U660 ( .A(n581), .B(KEYINPUT18), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G135), .A2(n869), .ZN(n583) );
  NAND2_X1 U662 ( .A1(G111), .A2(n861), .ZN(n582) );
  NAND2_X1 U663 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U664 ( .A1(G99), .A2(n866), .ZN(n584) );
  XNOR2_X1 U665 ( .A(KEYINPUT71), .B(n584), .ZN(n585) );
  NOR2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U668 ( .A(KEYINPUT72), .B(n589), .Z(n914) );
  XNOR2_X1 U669 ( .A(n914), .B(G2096), .ZN(n591) );
  INV_X1 U670 ( .A(G2100), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(G156) );
  XNOR2_X1 U672 ( .A(n969), .B(KEYINPUT73), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n891), .A2(G559), .ZN(n592) );
  XOR2_X1 U674 ( .A(n593), .B(n592), .Z(n637) );
  NOR2_X1 U675 ( .A1(n637), .A2(G860), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G67), .A2(n628), .ZN(n595) );
  NAND2_X1 U677 ( .A1(G55), .A2(n624), .ZN(n594) );
  NAND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U679 ( .A1(G93), .A2(n615), .ZN(n597) );
  NAND2_X1 U680 ( .A1(G80), .A2(n618), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U682 ( .A1(n599), .A2(n598), .ZN(n640) );
  XNOR2_X1 U683 ( .A(n600), .B(n640), .ZN(G145) );
  AND2_X1 U684 ( .A1(n615), .A2(G85), .ZN(n604) );
  NAND2_X1 U685 ( .A1(G60), .A2(n628), .ZN(n602) );
  NAND2_X1 U686 ( .A1(G47), .A2(n624), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n618), .A2(G72), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(G290) );
  NAND2_X1 U691 ( .A1(G62), .A2(n628), .ZN(n608) );
  NAND2_X1 U692 ( .A1(G50), .A2(n624), .ZN(n607) );
  NAND2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U694 ( .A(KEYINPUT74), .B(n609), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G88), .A2(n615), .ZN(n611) );
  NAND2_X1 U696 ( .A1(G75), .A2(n618), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U699 ( .A(KEYINPUT75), .B(n614), .Z(G166) );
  NAND2_X1 U700 ( .A1(G86), .A2(n615), .ZN(n617) );
  NAND2_X1 U701 ( .A1(G48), .A2(n624), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n618), .A2(G73), .ZN(n619) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n619), .Z(n620) );
  NOR2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n628), .A2(G61), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G49), .A2(n624), .ZN(n626) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(G288) );
  XNOR2_X1 U714 ( .A(n966), .B(G290), .ZN(n634) );
  XNOR2_X1 U715 ( .A(G166), .B(n640), .ZN(n632) );
  XNOR2_X1 U716 ( .A(n632), .B(G305), .ZN(n633) );
  XNOR2_X1 U717 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U718 ( .A(KEYINPUT19), .B(n635), .ZN(n636) );
  XNOR2_X1 U719 ( .A(n636), .B(G288), .ZN(n889) );
  XOR2_X1 U720 ( .A(n889), .B(n637), .Z(n638) );
  NAND2_X1 U721 ( .A1(n638), .A2(G868), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U724 ( .A(KEYINPUT76), .B(n643), .Z(G295) );
  NAND2_X1 U725 ( .A1(G2084), .A2(G2078), .ZN(n644) );
  XOR2_X1 U726 ( .A(KEYINPUT20), .B(n644), .Z(n645) );
  NAND2_X1 U727 ( .A1(G2090), .A2(n645), .ZN(n647) );
  XOR2_X1 U728 ( .A(KEYINPUT21), .B(KEYINPUT77), .Z(n646) );
  XNOR2_X1 U729 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U730 ( .A1(G2072), .A2(n648), .ZN(G158) );
  XNOR2_X1 U731 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U732 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U733 ( .A1(G108), .A2(G120), .ZN(n649) );
  NOR2_X1 U734 ( .A1(G237), .A2(n649), .ZN(n650) );
  NAND2_X1 U735 ( .A1(G69), .A2(n650), .ZN(n822) );
  NAND2_X1 U736 ( .A1(G567), .A2(n822), .ZN(n655) );
  NOR2_X1 U737 ( .A1(G220), .A2(G219), .ZN(n651) );
  XOR2_X1 U738 ( .A(KEYINPUT22), .B(n651), .Z(n652) );
  NOR2_X1 U739 ( .A1(G218), .A2(n652), .ZN(n653) );
  NAND2_X1 U740 ( .A1(G96), .A2(n653), .ZN(n823) );
  NAND2_X1 U741 ( .A1(G2106), .A2(n823), .ZN(n654) );
  NAND2_X1 U742 ( .A1(n655), .A2(n654), .ZN(n843) );
  NAND2_X1 U743 ( .A1(G661), .A2(G483), .ZN(n656) );
  NOR2_X1 U744 ( .A1(n843), .A2(n656), .ZN(n821) );
  NAND2_X1 U745 ( .A1(n821), .A2(G36), .ZN(G176) );
  NAND2_X1 U746 ( .A1(G138), .A2(n869), .ZN(n658) );
  NAND2_X1 U747 ( .A1(G102), .A2(n866), .ZN(n657) );
  NAND2_X1 U748 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U749 ( .A(n659), .B(KEYINPUT78), .ZN(n663) );
  NAND2_X1 U750 ( .A1(n861), .A2(G114), .ZN(n661) );
  NAND2_X1 U751 ( .A1(G126), .A2(n862), .ZN(n660) );
  NAND2_X1 U752 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U753 ( .A(KEYINPUT79), .B(G166), .ZN(G303) );
  NAND2_X1 U754 ( .A1(G160), .A2(G40), .ZN(n756) );
  XNOR2_X1 U755 ( .A(KEYINPUT85), .B(n756), .ZN(n664) );
  NAND2_X1 U756 ( .A1(n664), .A2(n757), .ZN(n668) );
  NAND2_X1 U757 ( .A1(G8), .A2(n668), .ZN(n749) );
  NOR2_X1 U758 ( .A1(G1971), .A2(n749), .ZN(n666) );
  NOR2_X1 U759 ( .A1(G2090), .A2(n702), .ZN(n665) );
  NOR2_X1 U760 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U761 ( .A1(G303), .A2(n667), .ZN(n716) );
  NAND2_X1 U762 ( .A1(n702), .A2(G1341), .ZN(n672) );
  INV_X1 U763 ( .A(G1996), .ZN(n794) );
  NOR2_X1 U764 ( .A1(n668), .A2(n794), .ZN(n670) );
  XNOR2_X1 U765 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U766 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U767 ( .A(n674), .B(KEYINPUT64), .Z(n680) );
  OR2_X1 U768 ( .A1(n680), .A2(n974), .ZN(n679) );
  AND2_X1 U769 ( .A1(n696), .A2(G2067), .ZN(n675) );
  XOR2_X1 U770 ( .A(n675), .B(KEYINPUT90), .Z(n677) );
  NAND2_X1 U771 ( .A1(n702), .A2(G1348), .ZN(n676) );
  NAND2_X1 U772 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U773 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n680), .A2(n974), .ZN(n681) );
  NAND2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n689) );
  XOR2_X1 U776 ( .A(KEYINPUT89), .B(KEYINPUT27), .Z(n684) );
  NAND2_X1 U777 ( .A1(G2072), .A2(n696), .ZN(n683) );
  XNOR2_X1 U778 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U779 ( .A(KEYINPUT88), .B(n685), .ZN(n687) );
  INV_X1 U780 ( .A(G1956), .ZN(n988) );
  NOR2_X1 U781 ( .A1(n696), .A2(n988), .ZN(n686) );
  NOR2_X1 U782 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n966), .A2(n690), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n693) );
  NOR2_X1 U785 ( .A1(n966), .A2(n690), .ZN(n691) );
  XOR2_X1 U786 ( .A(n691), .B(KEYINPUT28), .Z(n692) );
  NAND2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n695) );
  XNOR2_X1 U788 ( .A(KEYINPUT91), .B(KEYINPUT29), .ZN(n694) );
  XNOR2_X1 U789 ( .A(n695), .B(n694), .ZN(n700) );
  OR2_X1 U790 ( .A1(n696), .A2(G1961), .ZN(n698) );
  XNOR2_X1 U791 ( .A(KEYINPUT25), .B(G2078), .ZN(n933) );
  NAND2_X1 U792 ( .A1(n696), .A2(n933), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n707), .A2(G171), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n712) );
  NOR2_X1 U796 ( .A1(n749), .A2(G1966), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n701), .B(KEYINPUT87), .ZN(n720) );
  INV_X1 U798 ( .A(G8), .ZN(n703) );
  NOR2_X1 U799 ( .A1(G2084), .A2(n702), .ZN(n719) );
  NOR2_X1 U800 ( .A1(n703), .A2(n719), .ZN(n704) );
  AND2_X1 U801 ( .A1(n720), .A2(n704), .ZN(n705) );
  XOR2_X1 U802 ( .A(KEYINPUT30), .B(n705), .Z(n706) );
  NOR2_X1 U803 ( .A1(G168), .A2(n706), .ZN(n709) );
  NOR2_X1 U804 ( .A1(G171), .A2(n707), .ZN(n708) );
  NOR2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U806 ( .A(KEYINPUT31), .B(n710), .Z(n711) );
  NAND2_X1 U807 ( .A1(G286), .A2(n721), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n717), .A2(G8), .ZN(n718) );
  XNOR2_X1 U810 ( .A(n718), .B(KEYINPUT32), .ZN(n727) );
  NAND2_X1 U811 ( .A1(G8), .A2(n719), .ZN(n725) );
  INV_X1 U812 ( .A(n720), .ZN(n723) );
  XOR2_X1 U813 ( .A(n721), .B(KEYINPUT92), .Z(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n740) );
  NOR2_X1 U817 ( .A1(G2090), .A2(G303), .ZN(n728) );
  NAND2_X1 U818 ( .A1(G8), .A2(n728), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n740), .A2(n729), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n749), .ZN(n733) );
  XNOR2_X1 U821 ( .A(n733), .B(KEYINPUT98), .ZN(n738) );
  NOR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n734) );
  XOR2_X1 U823 ( .A(n734), .B(KEYINPUT86), .Z(n735) );
  XNOR2_X1 U824 ( .A(KEYINPUT24), .B(n735), .ZN(n736) );
  OR2_X1 U825 ( .A1(n749), .A2(n736), .ZN(n737) );
  AND2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n755) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n746) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n746), .A2(n739), .ZN(n977) );
  NAND2_X1 U830 ( .A1(n977), .A2(n740), .ZN(n741) );
  XNOR2_X1 U831 ( .A(n741), .B(KEYINPUT94), .ZN(n744) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n967) );
  INV_X1 U833 ( .A(n967), .ZN(n742) );
  NOR2_X1 U834 ( .A1(n749), .A2(n742), .ZN(n743) );
  AND2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(n745), .ZN(n752) );
  NAND2_X1 U837 ( .A1(KEYINPUT33), .A2(n746), .ZN(n747) );
  XOR2_X1 U838 ( .A(KEYINPUT95), .B(n747), .Z(n748) );
  NOR2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U840 ( .A(n750), .B(KEYINPUT96), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n958) );
  NAND2_X1 U843 ( .A1(n753), .A2(n958), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n788) );
  XNOR2_X1 U845 ( .A(G1986), .B(G290), .ZN(n965) );
  NOR2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n802) );
  AND2_X1 U847 ( .A1(n965), .A2(n802), .ZN(n786) );
  XOR2_X1 U848 ( .A(KEYINPUT83), .B(G1991), .Z(n934) );
  NAND2_X1 U849 ( .A1(G95), .A2(n866), .ZN(n759) );
  NAND2_X1 U850 ( .A1(G107), .A2(n861), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U852 ( .A1(G131), .A2(n869), .ZN(n761) );
  NAND2_X1 U853 ( .A1(G119), .A2(n862), .ZN(n760) );
  NAND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U856 ( .A(n764), .B(KEYINPUT82), .Z(n875) );
  AND2_X1 U857 ( .A1(n934), .A2(n875), .ZN(n919) );
  NAND2_X1 U858 ( .A1(G105), .A2(n866), .ZN(n765) );
  XNOR2_X1 U859 ( .A(n765), .B(KEYINPUT38), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G141), .A2(n869), .ZN(n766) );
  XNOR2_X1 U861 ( .A(n766), .B(KEYINPUT84), .ZN(n767) );
  NAND2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n861), .A2(G117), .ZN(n770) );
  NAND2_X1 U864 ( .A1(G129), .A2(n862), .ZN(n769) );
  NAND2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n876) );
  NOR2_X1 U867 ( .A1(n876), .A2(n794), .ZN(n913) );
  OR2_X1 U868 ( .A1(n919), .A2(n913), .ZN(n773) );
  NAND2_X1 U869 ( .A1(n802), .A2(n773), .ZN(n790) );
  XNOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .ZN(n789) );
  XNOR2_X1 U871 ( .A(KEYINPUT81), .B(KEYINPUT36), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n861), .A2(G116), .ZN(n775) );
  NAND2_X1 U873 ( .A1(G128), .A2(n862), .ZN(n774) );
  NAND2_X1 U874 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U875 ( .A(KEYINPUT35), .B(n776), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n869), .A2(G140), .ZN(n777) );
  XNOR2_X1 U877 ( .A(n777), .B(KEYINPUT80), .ZN(n779) );
  NAND2_X1 U878 ( .A1(G104), .A2(n866), .ZN(n778) );
  NAND2_X1 U879 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U880 ( .A(KEYINPUT34), .B(n780), .Z(n781) );
  NAND2_X1 U881 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U882 ( .A(n784), .B(n783), .ZN(n885) );
  NOR2_X1 U883 ( .A1(n789), .A2(n885), .ZN(n923) );
  NAND2_X1 U884 ( .A1(n802), .A2(n923), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n790), .A2(n799), .ZN(n785) );
  NOR2_X1 U886 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U887 ( .A1(n788), .A2(n787), .ZN(n805) );
  NAND2_X1 U888 ( .A1(n789), .A2(n885), .ZN(n924) );
  INV_X1 U889 ( .A(n790), .ZN(n793) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n791) );
  NOR2_X1 U891 ( .A1(n934), .A2(n875), .ZN(n915) );
  NOR2_X1 U892 ( .A1(n791), .A2(n915), .ZN(n792) );
  NOR2_X1 U893 ( .A1(n793), .A2(n792), .ZN(n795) );
  AND2_X1 U894 ( .A1(n794), .A2(n876), .ZN(n908) );
  NOR2_X1 U895 ( .A1(n795), .A2(n908), .ZN(n797) );
  XOR2_X1 U896 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n796) );
  XNOR2_X1 U897 ( .A(n797), .B(n796), .ZN(n798) );
  NAND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n924), .A2(n800), .ZN(n801) );
  XNOR2_X1 U900 ( .A(KEYINPUT100), .B(n801), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U903 ( .A(n806), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U904 ( .A(KEYINPUT101), .B(G2446), .Z(n808) );
  XNOR2_X1 U905 ( .A(G2435), .B(G2438), .ZN(n807) );
  XNOR2_X1 U906 ( .A(n808), .B(n807), .ZN(n815) );
  XOR2_X1 U907 ( .A(G2451), .B(G2430), .Z(n810) );
  XNOR2_X1 U908 ( .A(G2454), .B(G2427), .ZN(n809) );
  XNOR2_X1 U909 ( .A(n810), .B(n809), .ZN(n811) );
  XOR2_X1 U910 ( .A(n811), .B(G2443), .Z(n813) );
  XNOR2_X1 U911 ( .A(G1341), .B(G1348), .ZN(n812) );
  XNOR2_X1 U912 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U913 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n816), .A2(G14), .ZN(n898) );
  XOR2_X1 U915 ( .A(KEYINPUT102), .B(n898), .Z(G401) );
  NAND2_X1 U916 ( .A1(n817), .A2(G2106), .ZN(n818) );
  XOR2_X1 U917 ( .A(KEYINPUT103), .B(n818), .Z(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U919 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U921 ( .A1(n821), .A2(n820), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n823), .A2(n822), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XOR2_X1 U929 ( .A(G2100), .B(G2096), .Z(n825) );
  XNOR2_X1 U930 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n824) );
  XNOR2_X1 U931 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U932 ( .A(G2678), .B(G2090), .Z(n827) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n826) );
  XNOR2_X1 U934 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U935 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U936 ( .A(G2084), .B(G2078), .ZN(n830) );
  XNOR2_X1 U937 ( .A(n831), .B(n830), .ZN(G227) );
  XOR2_X1 U938 ( .A(KEYINPUT106), .B(G1956), .Z(n833) );
  XNOR2_X1 U939 ( .A(G1981), .B(G1966), .ZN(n832) );
  XNOR2_X1 U940 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U941 ( .A(n834), .B(KEYINPUT41), .Z(n836) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U943 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U944 ( .A(G1961), .B(G1971), .Z(n838) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1976), .ZN(n837) );
  XNOR2_X1 U946 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U947 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U948 ( .A(KEYINPUT105), .B(G2474), .ZN(n841) );
  XNOR2_X1 U949 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U950 ( .A(KEYINPUT104), .B(n843), .Z(G319) );
  NAND2_X1 U951 ( .A1(G136), .A2(n869), .ZN(n845) );
  NAND2_X1 U952 ( .A1(G112), .A2(n861), .ZN(n844) );
  NAND2_X1 U953 ( .A1(n845), .A2(n844), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n862), .A2(G124), .ZN(n846) );
  XNOR2_X1 U955 ( .A(n846), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U956 ( .A1(G100), .A2(n866), .ZN(n847) );
  XOR2_X1 U957 ( .A(KEYINPUT107), .B(n847), .Z(n848) );
  NAND2_X1 U958 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U959 ( .A1(n851), .A2(n850), .ZN(G162) );
  NAND2_X1 U960 ( .A1(G142), .A2(n869), .ZN(n853) );
  NAND2_X1 U961 ( .A1(G106), .A2(n866), .ZN(n852) );
  NAND2_X1 U962 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U963 ( .A(n854), .B(KEYINPUT45), .ZN(n856) );
  NAND2_X1 U964 ( .A1(G118), .A2(n861), .ZN(n855) );
  NAND2_X1 U965 ( .A1(n856), .A2(n855), .ZN(n859) );
  NAND2_X1 U966 ( .A1(n862), .A2(G130), .ZN(n857) );
  XOR2_X1 U967 ( .A(KEYINPUT108), .B(n857), .Z(n858) );
  NOR2_X1 U968 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U969 ( .A(n914), .B(n860), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n861), .A2(G115), .ZN(n864) );
  NAND2_X1 U971 ( .A1(G127), .A2(n862), .ZN(n863) );
  NAND2_X1 U972 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U973 ( .A(n865), .B(KEYINPUT47), .ZN(n868) );
  NAND2_X1 U974 ( .A1(G103), .A2(n866), .ZN(n867) );
  NAND2_X1 U975 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n869), .A2(G139), .ZN(n870) );
  XOR2_X1 U977 ( .A(KEYINPUT110), .B(n870), .Z(n871) );
  NOR2_X1 U978 ( .A1(n872), .A2(n871), .ZN(n903) );
  XNOR2_X1 U979 ( .A(G164), .B(n903), .ZN(n873) );
  XNOR2_X1 U980 ( .A(n874), .B(n873), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT109), .B(KEYINPUT111), .Z(n878) );
  XNOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n877) );
  XNOR2_X1 U984 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U985 ( .A(n879), .B(KEYINPUT46), .Z(n881) );
  XNOR2_X1 U986 ( .A(G160), .B(G162), .ZN(n880) );
  XNOR2_X1 U987 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U988 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U989 ( .A(n885), .B(n884), .Z(n886) );
  XNOR2_X1 U990 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U991 ( .A1(G37), .A2(n888), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(n969), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n893) );
  XOR2_X1 U994 ( .A(G171), .B(n891), .Z(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U996 ( .A1(G37), .A2(n894), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(n895), .Z(G397) );
  XNOR2_X1 U998 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n897) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n896) );
  XNOR2_X1 U1000 ( .A(n897), .B(n896), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n898), .ZN(n899) );
  NOR2_X1 U1002 ( .A1(n900), .A2(n899), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n901) );
  NAND2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(KEYINPUT55), .ZN(n954) );
  XOR2_X1 U1007 ( .A(G2072), .B(n903), .Z(n905) );
  XOR2_X1 U1008 ( .A(G164), .B(G2078), .Z(n904) );
  NOR2_X1 U1009 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(KEYINPUT50), .B(n906), .ZN(n928) );
  XOR2_X1 U1011 ( .A(G2090), .B(G162), .Z(n907) );
  NOR2_X1 U1012 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1013 ( .A(KEYINPUT51), .B(n909), .Z(n910) );
  XNOR2_X1 U1014 ( .A(KEYINPUT116), .B(n910), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G160), .B(G2084), .ZN(n911) );
  XNOR2_X1 U1016 ( .A(n911), .B(KEYINPUT115), .ZN(n912) );
  NOR2_X1 U1017 ( .A1(n913), .A2(n912), .ZN(n917) );
  NOR2_X1 U1018 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT117), .B(n926), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n929), .B(KEYINPUT52), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT118), .B(n930), .Z(n931) );
  NAND2_X1 U1028 ( .A1(n954), .A2(n931), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n932), .A2(G29), .ZN(n987) );
  XOR2_X1 U1030 ( .A(n933), .B(G27), .Z(n936) );
  XNOR2_X1 U1031 ( .A(n934), .B(G25), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(G1996), .B(G32), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(G33), .B(G2072), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(G28), .A2(n939), .ZN(n942) );
  XOR2_X1 U1037 ( .A(G26), .B(G2067), .Z(n940) );
  XNOR2_X1 U1038 ( .A(KEYINPUT119), .B(n940), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT53), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT120), .B(n946), .ZN(n952) );
  XOR2_X1 U1043 ( .A(KEYINPUT121), .B(G34), .Z(n948) );
  XNOR2_X1 U1044 ( .A(G2084), .B(KEYINPUT54), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(n948), .B(n947), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G35), .B(G2090), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n954), .B(n953), .ZN(n956) );
  INV_X1 U1050 ( .A(G29), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n957), .ZN(n985) );
  XOR2_X1 U1053 ( .A(G16), .B(KEYINPUT56), .Z(n982) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(n960), .B(KEYINPUT122), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(KEYINPUT57), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n980) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G301), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(G1956), .B(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G1341), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n974), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1072 ( .A(KEYINPUT123), .B(n983), .Z(n984) );
  NOR2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n1015) );
  XNOR2_X1 U1075 ( .A(n988), .B(G20), .ZN(n997) );
  XOR2_X1 U1076 ( .A(G4), .B(KEYINPUT126), .Z(n990) );
  XNOR2_X1 U1077 ( .A(G1348), .B(KEYINPUT59), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n990), .B(n989), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(G1981), .B(G6), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G19), .B(G1341), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n993), .B(KEYINPUT125), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(n998), .B(KEYINPUT60), .ZN(n1010) );
  XOR2_X1 U1086 ( .A(G1986), .B(G24), .Z(n1002) );
  XNOR2_X1 U1087 ( .A(G1976), .B(G23), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1004), .B(n1003), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G5), .B(G1961), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1011), .Z(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT124), .B(G16), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1016), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

