//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n438, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n438), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT69), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n459), .A2(G101), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NOR3_X1   g045(.A1(new_n468), .A2(G2105), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n471), .B2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n469), .A2(new_n473), .A3(G125), .ZN(new_n474));
  AND3_X1   g049(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n466), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(new_n460), .A3(new_n469), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(G2105), .B(new_n469), .C1(new_n459), .C2(new_n463), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(G124), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT70), .ZN(G162));
  NAND2_X1  g066(.A1(new_n469), .A2(new_n473), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(new_n460), .A3(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n482), .A2(G138), .A3(new_n460), .A4(new_n469), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  NOR2_X1   g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(new_n460), .B2(G114), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n488), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT71), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n520), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n514), .B1(new_n522), .B2(new_n523), .C1(new_n524), .C2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  INV_X1    g103(.A(new_n522), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  INV_X1    g105(.A(new_n526), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n530), .A2(new_n532), .A3(new_n535), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(new_n531), .A2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n529), .A2(G52), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n515), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n511), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n529), .A2(G43), .B1(G651), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n531), .A2(G81), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n529), .A2(G53), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT73), .B(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n522), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT74), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n511), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n531), .A2(G91), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  OAI21_X1  g143(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n569));
  INV_X1    g144(.A(G49), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI221_X1 g146(.A(new_n569), .B1(new_n522), .B2(new_n570), .C1(new_n571), .C2(new_n526), .ZN(G288));
  NAND3_X1  g147(.A1(new_n508), .A2(new_n510), .A3(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n521), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n520), .A2(G86), .A3(new_n521), .A4(new_n525), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT75), .ZN(G305));
  NAND2_X1  g155(.A1(new_n531), .A2(G85), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n529), .A2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n581), .B(new_n582), .C1(new_n515), .C2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n531), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(new_n529), .A2(G54), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n515), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  XNOR2_X1  g173(.A(KEYINPUT76), .B(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(G860), .B2(new_n599), .ZN(G148));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n465), .A2(new_n467), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G2105), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n606), .A2(new_n469), .A3(new_n473), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n471), .A2(G135), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(KEYINPUT77), .B1(G123), .B2(new_n489), .ZN(new_n612));
  NOR2_X1   g187(.A1(G99), .A2(G2105), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n614));
  OAI221_X1 g189(.A(new_n612), .B1(KEYINPUT77), .B2(new_n611), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G2096), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT78), .Z(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2443), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G14), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2067), .B(G2678), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n641), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT83), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n638), .A2(new_n639), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(KEYINPUT83), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n647), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n652));
  NAND4_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n640), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n644), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n616), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n662), .A2(KEYINPUT20), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n658), .A3(new_n661), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n665), .B(new_n667), .C1(KEYINPUT20), .C2(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(G229));
  INV_X1    g249(.A(G29), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G26), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n489), .A2(G128), .ZN(new_n677));
  INV_X1    g252(.A(G140), .ZN(new_n678));
  NOR2_X1   g253(.A1(G104), .A2(G2105), .ZN(new_n679));
  OAI21_X1  g254(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n680));
  OAI22_X1  g255(.A1(new_n483), .A2(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n676), .B1(new_n683), .B2(new_n675), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n676), .B(new_n684), .S(KEYINPUT28), .Z(new_n685));
  INV_X1    g260(.A(G2067), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(G160), .A2(G29), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G34), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n688), .B1(G29), .B2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G2084), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(G171), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G5), .B2(G16), .ZN(new_n695));
  INV_X1    g270(.A(G1961), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(G29), .A2(G32), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n489), .A2(G129), .B1(G105), .B2(new_n606), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT26), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n471), .A2(G141), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n698), .B1(new_n703), .B2(new_n675), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n687), .A2(new_n693), .A3(new_n697), .A4(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n691), .A2(new_n692), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(KEYINPUT90), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT85), .B(G16), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n550), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G19), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n715), .B2(G1341), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G1341), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n471), .A2(G139), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT87), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT25), .Z(new_n721));
  AND2_X1   g296(.A1(new_n469), .A2(new_n473), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n722), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n719), .B(new_n721), .C1(new_n460), .C2(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G33), .B(new_n724), .S(G29), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT88), .B(G2072), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n707), .A2(new_n708), .A3(new_n717), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G35), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G162), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2090), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n712), .A2(KEYINPUT23), .A3(G20), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT23), .ZN(new_n734));
  INV_X1    g309(.A(G20), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n711), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n733), .B(new_n736), .C1(new_n596), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT97), .B(G1956), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n695), .A2(new_n696), .ZN(new_n742));
  NAND2_X1  g317(.A1(G168), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G16), .B2(G21), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n615), .A2(new_n675), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n675), .B1(new_n748), .B2(G28), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(G28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AND4_X1   g328(.A1(new_n742), .A2(new_n746), .A3(new_n747), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n744), .A2(new_n745), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT92), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT93), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n737), .A2(G4), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n592), .B2(new_n737), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G1348), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n675), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n675), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n765), .B(new_n766), .S(KEYINPUT94), .Z(new_n767));
  XOR2_X1   g342(.A(KEYINPUT95), .B(G2078), .Z(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT96), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n767), .B(new_n769), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n764), .B(new_n770), .C1(KEYINPUT90), .C2(new_n709), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n728), .A2(new_n741), .A3(new_n759), .A4(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G24), .B(G290), .S(new_n711), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1986), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n737), .A2(G23), .ZN(new_n775));
  INV_X1    g350(.A(G288), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n737), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT33), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1976), .ZN(new_n779));
  MUX2_X1   g354(.A(G6), .B(G305), .S(G16), .Z(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n712), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n712), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT86), .B(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n779), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n774), .B1(new_n787), .B2(KEYINPUT34), .ZN(new_n788));
  OR2_X1    g363(.A1(G95), .A2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n789), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n790));
  INV_X1    g365(.A(G119), .ZN(new_n791));
  INV_X1    g366(.A(G131), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n790), .B1(new_n488), .B2(new_n791), .C1(new_n483), .C2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT84), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT35), .B(G1991), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n788), .B(new_n797), .C1(KEYINPUT34), .C2(new_n787), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT36), .Z(new_n799));
  AOI211_X1 g374(.A(new_n772), .B(new_n799), .C1(new_n763), .C2(new_n762), .ZN(G311));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n772), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G1348), .B2(new_n761), .ZN(G150));
  NAND2_X1  g377(.A1(new_n531), .A2(G93), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n529), .A2(G55), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n803), .B(new_n804), .C1(new_n515), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G860), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n592), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n550), .B(new_n806), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT99), .Z(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT100), .Z(new_n819));
  OAI21_X1  g394(.A(new_n809), .B1(new_n817), .B2(new_n819), .ZN(G145));
  XNOR2_X1  g395(.A(new_n682), .B(new_n504), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n703), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n724), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n724), .A2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n824), .B2(new_n822), .ZN(new_n827));
  XNOR2_X1  g402(.A(G162), .B(G160), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n489), .A2(G130), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT103), .Z(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT104), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(KEYINPUT104), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n833), .B(new_n834), .C1(G118), .C2(new_n460), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n471), .A2(G142), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n793), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT105), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n615), .B(new_n608), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n829), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n829), .A2(new_n841), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g421(.A1(new_n596), .A2(new_n591), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n592), .A2(G299), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(KEYINPUT41), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n601), .B(new_n813), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n849), .B2(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT108), .ZN(new_n857));
  XNOR2_X1  g432(.A(G303), .B(G288), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G305), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(G290), .Z(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n859), .B(G290), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT42), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n857), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT108), .B1(new_n860), .B2(new_n861), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n856), .A2(new_n867), .ZN(new_n868));
  OAI221_X1 g443(.A(new_n855), .B1(new_n849), .B2(new_n854), .C1(new_n865), .C2(new_n866), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n869), .A3(G868), .ZN(new_n870));
  INV_X1    g445(.A(G868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n806), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  MUX2_X1   g448(.A(new_n870), .B(new_n873), .S(KEYINPUT109), .Z(G295));
  MUX2_X1   g449(.A(new_n870), .B(new_n873), .S(KEYINPUT109), .Z(G331));
  XNOR2_X1  g450(.A(G171), .B(G286), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n813), .B(new_n876), .Z(new_n877));
  INV_X1    g452(.A(KEYINPUT111), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n813), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n877), .B2(KEYINPUT111), .ZN(new_n880));
  OAI22_X1  g455(.A1(new_n853), .A2(new_n877), .B1(new_n880), .B2(new_n850), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n860), .ZN(new_n882));
  OAI221_X1 g457(.A(new_n863), .B1(new_n880), .B2(new_n850), .C1(new_n853), .C2(new_n877), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n843), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n849), .A2(new_n852), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n880), .B(new_n886), .C1(KEYINPUT41), .C2(new_n849), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n877), .A2(new_n849), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n863), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n883), .A2(new_n890), .A3(new_n891), .A4(new_n843), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n883), .A2(new_n890), .A3(new_n843), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT43), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n884), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(G397));
  INV_X1    g474(.A(KEYINPUT121), .ZN(new_n900));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n497), .B2(new_n502), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n472), .A2(KEYINPUT112), .A3(G40), .A4(new_n478), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n482), .A2(G137), .A3(new_n460), .A4(new_n469), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n906), .A2(new_n478), .A3(G40), .A4(new_n461), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT112), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(KEYINPUT45), .B(new_n901), .C1(new_n497), .C2(new_n502), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G1971), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n915));
  INV_X1    g490(.A(G2090), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT50), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(new_n901), .C1(new_n497), .C2(new_n502), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n915), .A2(new_n910), .A3(new_n916), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(G303), .A2(G8), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(G8), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT114), .ZN(new_n925));
  INV_X1    g500(.A(G8), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n914), .B2(new_n919), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT114), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n923), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n912), .A2(new_n745), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n915), .A2(new_n910), .A3(new_n692), .A4(new_n918), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(G8), .A3(G168), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT119), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT119), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n933), .A2(new_n936), .A3(G8), .A4(G168), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT117), .B1(new_n927), .B2(new_n923), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT117), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n915), .A2(new_n910), .A3(new_n918), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n941), .A2(new_n916), .B1(new_n912), .B2(new_n913), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n940), .B(new_n922), .C1(new_n942), .C2(new_n926), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n579), .A2(G1981), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1981), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n576), .A2(new_n947), .A3(new_n577), .A4(new_n578), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT115), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n902), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n910), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(new_n949), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT49), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n945), .A3(new_n951), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n956), .A3(new_n959), .A4(G8), .ZN(new_n960));
  INV_X1    g535(.A(G1976), .ZN(new_n961));
  NOR2_X1   g536(.A1(G288), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(G288), .B2(new_n961), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n956), .A2(G8), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI211_X1 g540(.A(new_n926), .B(new_n962), .C1(new_n910), .C2(new_n955), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n960), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT118), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n956), .A2(G8), .A3(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT118), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n960), .A4(new_n965), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n930), .A2(new_n938), .A3(new_n944), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT120), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT63), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  INV_X1    g554(.A(new_n968), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n927), .A2(new_n923), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(new_n977), .ZN(new_n982));
  AND4_X1   g557(.A1(new_n930), .A2(new_n938), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n978), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n925), .A2(new_n929), .A3(new_n980), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n960), .A2(new_n961), .A3(new_n776), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n948), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(G8), .A3(new_n956), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n989), .A2(KEYINPUT116), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(KEYINPUT116), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n900), .B1(new_n984), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n994));
  NAND2_X1  g569(.A1(G286), .A2(G8), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n941), .A2(new_n692), .B1(new_n912), .B2(new_n745), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n994), .B(new_n995), .C1(new_n996), .C2(new_n926), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT51), .B(G8), .C1(new_n933), .C2(G286), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n933), .A2(G8), .A3(G286), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT62), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT62), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1003), .A3(new_n1000), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n930), .A2(new_n944), .A3(new_n974), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n912), .A2(G2078), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n915), .A2(new_n910), .A3(new_n918), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1007), .A2(new_n1008), .B1(new_n696), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(G171), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1005), .A2(KEYINPUT125), .A3(new_n1006), .A4(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1006), .A2(new_n1002), .A3(new_n1012), .A4(new_n1004), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT125), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n907), .B(KEYINPUT112), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(new_n902), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n686), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1009), .A2(new_n763), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n592), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n591), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT60), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1021), .A2(KEYINPUT60), .A3(new_n591), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT58), .B(G1341), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n912), .A2(G1996), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n550), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT123), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(KEYINPUT123), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1024), .A2(new_n1025), .A3(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT56), .B(G2072), .Z(new_n1036));
  OR2_X1    g611(.A1(new_n912), .A2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n941), .A2(KEYINPUT122), .A3(G1956), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  INV_X1    g614(.A(G1956), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1009), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1037), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n562), .A2(new_n1043), .A3(new_n567), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT61), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1045), .B(new_n1037), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1034), .B(new_n1035), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1023), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n1047), .ZN(new_n1054));
  XOR2_X1   g629(.A(G301), .B(KEYINPUT54), .Z(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1011), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n904), .A2(new_n911), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n472), .A2(G40), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1058), .A2(G2078), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n474), .A2(new_n477), .ZN(new_n1061));
  XOR2_X1   g636(.A(new_n1061), .B(KEYINPUT124), .Z(new_n1062));
  OAI211_X1 g637(.A(new_n1060), .B(KEYINPUT53), .C1(new_n460), .C2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1010), .A2(new_n1055), .A3(new_n1063), .ZN(new_n1064));
  AND4_X1   g639(.A1(new_n1057), .A2(new_n1006), .A3(new_n1001), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1013), .A2(new_n1016), .B1(new_n1054), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n990), .A2(new_n991), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n975), .A2(new_n977), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT120), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT121), .B(new_n1067), .C1(new_n1071), .C2(new_n983), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n993), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1017), .A2(new_n904), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n682), .B(G2067), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n703), .B(G1996), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT113), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n793), .A2(new_n796), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n793), .A2(new_n796), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(G290), .B(G1986), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1074), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1073), .A2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1017), .A2(new_n904), .A3(G1996), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1086), .A2(KEYINPUT46), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1074), .B1(new_n1075), .B2(new_n703), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(KEYINPUT46), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n1090), .B(KEYINPUT47), .Z(new_n1091));
  NOR2_X1   g666(.A1(G290), .A2(G1986), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT48), .B1(new_n1074), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1074), .A2(KEYINPUT48), .A3(new_n1092), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1082), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1080), .B(KEYINPUT126), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1078), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(G2067), .B2(new_n682), .ZN(new_n1098));
  AOI211_X1 g673(.A(new_n1091), .B(new_n1095), .C1(new_n1074), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1085), .A2(new_n1099), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g675(.A(G229), .ZN(new_n1102));
  AND2_X1   g676(.A1(new_n845), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g677(.A(G319), .ZN(new_n1104));
  OR2_X1    g678(.A1(G227), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g679(.A(new_n635), .B1(KEYINPUT127), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g680(.A(new_n1106), .B1(KEYINPUT127), .B2(new_n1105), .ZN(new_n1107));
  AND3_X1   g681(.A1(new_n1103), .A2(new_n893), .A3(new_n1107), .ZN(G308));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n893), .A3(new_n1107), .ZN(G225));
endmodule


