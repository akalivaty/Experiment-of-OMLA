//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT70), .Z(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n195), .A2(KEYINPUT65), .A3(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT65), .B1(new_n195), .B2(G146), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n192), .B(new_n194), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(G143), .B2(new_n191), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n202), .B2(new_n193), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(G137), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n211), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n206), .A2(G137), .ZN(new_n214));
  OAI21_X1  g028(.A(G131), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n212), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n195), .A2(G146), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n191), .B2(G143), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n195), .A2(KEYINPUT65), .A3(G146), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n224), .A2(new_n225), .B1(new_n200), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT2), .B(G113), .Z(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G116), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT67), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n234), .A2(new_n241), .B1(new_n239), .B2(new_n240), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n230), .A2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n216), .A2(new_n229), .A3(KEYINPUT30), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n219), .A2(new_n228), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n219), .B2(new_n228), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n216), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n244), .B1(new_n251), .B2(new_n243), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT31), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n245), .ZN(new_n259));
  INV_X1    g073(.A(new_n216), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n229), .A2(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n219), .A2(new_n228), .A3(new_n246), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n250), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n259), .B(new_n243), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n244), .ZN(new_n266));
  AND4_X1   g080(.A1(KEYINPUT31), .A2(new_n265), .A3(new_n266), .A4(new_n257), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n249), .A2(new_n269), .A3(new_n243), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n266), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n249), .B2(new_n243), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT28), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n244), .A2(KEYINPUT28), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n257), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n268), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n257), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n261), .A2(new_n262), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n242), .B1(new_n281), .B2(new_n216), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n244), .B1(new_n282), .B2(new_n269), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT68), .B1(new_n263), .B2(new_n242), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n279), .B1(new_n285), .B2(new_n274), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n265), .A2(new_n266), .A3(new_n257), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n252), .A2(KEYINPUT31), .A3(new_n257), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT69), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n190), .B1(new_n278), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n230), .A2(new_n243), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n266), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n230), .A2(KEYINPUT71), .A3(new_n243), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n274), .B1(new_n298), .B2(KEYINPUT28), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n279), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n273), .A2(new_n275), .A3(new_n257), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n252), .A2(new_n257), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G472), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n277), .B1(new_n268), .B2(new_n276), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n291), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n188), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n293), .B(new_n307), .C1(new_n310), .C2(KEYINPUT32), .ZN(new_n311));
  INV_X1    g125(.A(G469), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  INV_X1    g127(.A(G104), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n314), .B2(G107), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G104), .ZN(new_n318));
  INV_X1    g132(.A(G101), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(G107), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n315), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n314), .A2(G107), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n317), .A2(G104), .ZN(new_n323));
  OAI21_X1  g137(.A(G101), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n204), .A3(KEYINPUT10), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT78), .ZN(new_n327));
  INV_X1    g141(.A(new_n219), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n315), .A2(new_n318), .A3(new_n320), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G101), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n332), .A3(G101), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n228), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n224), .A2(new_n335), .A3(new_n194), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n198), .A2(KEYINPUT77), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n202), .A2(new_n193), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n224), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n325), .B(new_n336), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n327), .A2(new_n328), .A3(new_n334), .A4(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G140), .ZN(new_n344));
  INV_X1    g158(.A(G953), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G227), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n321), .A2(new_n324), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n198), .A3(new_n203), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT12), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n328), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n350), .B(new_n353), .C1(new_n351), .C2(new_n352), .ZN(new_n357));
  AND4_X1   g171(.A1(new_n343), .A2(new_n347), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n326), .B(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n342), .A2(new_n334), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n219), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n347), .B1(new_n362), .B2(new_n343), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n312), .B(new_n313), .C1(new_n358), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(G469), .A2(G902), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n343), .A2(new_n356), .A3(new_n357), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n347), .B(KEYINPUT76), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n343), .A3(new_n347), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(G469), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n364), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G221), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT9), .B(G234), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n372), .B1(new_n374), .B2(new_n313), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G125), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT73), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT73), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n191), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(G146), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT18), .A2(G131), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n392));
  AOI21_X1  g206(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n253), .A2(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n195), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n390), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n378), .B1(new_n389), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n394), .A2(new_n398), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n387), .A2(new_n388), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT84), .ZN(new_n403));
  OAI21_X1  g217(.A(G131), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n210), .A3(new_n397), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n379), .A3(G125), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n383), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n191), .ZN(new_n411));
  OAI211_X1 g225(.A(G146), .B(new_n409), .C1(new_n383), .C2(new_n408), .ZN(new_n412));
  OAI211_X1 g226(.A(KEYINPUT17), .B(G131), .C1(new_n392), .C2(new_n393), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n400), .A2(new_n403), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT86), .B(G104), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT88), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT87), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n407), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n401), .A2(KEYINPUT84), .A3(new_n402), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT84), .B1(new_n401), .B2(new_n402), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(KEYINPUT87), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n420), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(KEYINPUT87), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n400), .A2(new_n403), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n421), .A3(new_n423), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n429), .A2(new_n431), .A3(KEYINPUT88), .A4(new_n418), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n313), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G475), .ZN(new_n434));
  NOR2_X1   g248(.A1(G475), .A2(G902), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n385), .A2(new_n436), .A3(new_n386), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n383), .A2(KEYINPUT19), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n191), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n412), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT85), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n404), .A2(new_n405), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n443), .A3(new_n412), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n419), .B1(new_n445), .B2(new_n430), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n426), .A2(new_n418), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n435), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(new_n435), .C1(new_n446), .C2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n434), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT13), .B1(new_n193), .B2(G143), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(new_n206), .ZN(new_n455));
  XNOR2_X1  g269(.A(G128), .B(G143), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G116), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n237), .A2(G122), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n461), .A2(new_n317), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n317), .B1(new_n461), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n457), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n459), .B(KEYINPUT89), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n462), .B(KEYINPUT14), .ZN(new_n467));
  OAI21_X1  g281(.A(G107), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n461), .A2(new_n317), .A3(new_n462), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n456), .B(new_n206), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n374), .A2(G217), .A3(new_n345), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G478), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT15), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n453), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(G234), .A2(G237), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(G952), .A3(new_n345), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(G902), .A3(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT21), .B(G898), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G214), .B1(G237), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT80), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n234), .A2(new_n241), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n236), .A2(new_n238), .A3(KEYINPUT5), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(G113), .C1(KEYINPUT5), .C2(new_n236), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n348), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G113), .B1(new_n236), .B2(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT81), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n233), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(G113), .C1(new_n236), .C2(KEYINPUT5), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n503), .A2(new_n504), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n497), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n348), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n497), .A3(KEYINPUT83), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n501), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n497), .A2(new_n325), .A3(new_n499), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n331), .A2(new_n333), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(new_n494), .C1(new_n516), .C2(new_n242), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI22_X1  g332(.A1(new_n514), .A2(new_n518), .B1(new_n495), .B2(new_n494), .ZN(new_n519));
  MUX2_X1   g333(.A(new_n204), .B(new_n228), .S(G125), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n345), .A2(G224), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n520), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n515), .B1(new_n516), .B2(new_n242), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n493), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n517), .A3(KEYINPUT6), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n528), .A3(new_n493), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n520), .B(new_n521), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n313), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G210), .B1(G237), .B2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n519), .B2(new_n523), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n533), .A3(new_n531), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n489), .B(new_n491), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n377), .A2(new_n482), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G234), .ZN(new_n540));
  OAI21_X1  g354(.A(G217), .B1(new_n540), .B2(G902), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT72), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n235), .B2(G128), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n545), .B(new_n546), .C1(G119), .C2(new_n193), .ZN(new_n547));
  XNOR2_X1  g361(.A(G119), .B(G128), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT24), .B(G110), .Z(new_n549));
  OAI22_X1  g363(.A1(new_n547), .A2(G110), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n412), .A3(new_n387), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT74), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n550), .A2(KEYINPUT74), .A3(new_n412), .A4(new_n387), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n411), .A2(new_n412), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n547), .A2(G110), .B1(new_n548), .B2(new_n549), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n372), .A2(new_n540), .A3(G953), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  NAND3_X1  g375(.A1(new_n555), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n555), .B2(new_n558), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT25), .A3(new_n313), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n555), .A2(new_n558), .ZN(new_n567));
  INV_X1    g381(.A(new_n561), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n313), .A3(new_n562), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT25), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n543), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n542), .A2(G902), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT75), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n311), .A2(new_n539), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT90), .B(G101), .Z(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(G3));
  OAI21_X1  g394(.A(new_n313), .B1(new_n278), .B2(new_n292), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n310), .B1(new_n581), .B2(G472), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n377), .A2(new_n577), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n536), .A2(KEYINPUT91), .A3(new_n533), .A4(new_n531), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n586), .A2(new_n490), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n535), .A2(new_n588), .A3(new_n537), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n489), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n433), .A2(G475), .B1(new_n449), .B2(new_n451), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n478), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n476), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n475), .B1(new_n465), .B2(new_n471), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n597), .A2(KEYINPUT33), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n474), .B2(new_n476), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n595), .B(new_n596), .C1(new_n599), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n596), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT33), .B1(new_n597), .B2(new_n598), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n474), .A2(new_n600), .A3(new_n476), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT92), .B1(new_n477), .B2(G478), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n593), .A2(new_n594), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n585), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  AOI22_X1  g426(.A1(new_n452), .A2(KEYINPUT93), .B1(new_n433), .B2(G475), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n449), .A2(new_n614), .A3(new_n451), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n593), .A2(new_n480), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n585), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G107), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n555), .A2(new_n621), .A3(new_n558), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n555), .B2(new_n558), .ZN(new_n624));
  OAI22_X1  g438(.A1(new_n623), .A2(new_n624), .B1(KEYINPUT36), .B2(new_n568), .ZN(new_n625));
  INV_X1    g439(.A(new_n624), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n568), .A2(KEYINPUT36), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n622), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n625), .A2(new_n628), .A3(new_n575), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n566), .A2(new_n572), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n630), .B1(new_n631), .B2(new_n543), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n582), .A2(new_n539), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n485), .B1(new_n487), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n613), .A2(new_n481), .A3(new_n615), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n632), .A2(new_n589), .A3(new_n587), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n311), .A2(new_n641), .A3(new_n377), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT95), .B(G128), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G30));
  NAND2_X1  g458(.A1(new_n535), .A2(new_n537), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n632), .A2(new_n594), .A3(new_n480), .A4(new_n491), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(KEYINPUT98), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n637), .B(KEYINPUT39), .Z(new_n650));
  NAND3_X1  g464(.A1(new_n371), .A2(new_n376), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n649), .B(new_n653), .C1(KEYINPUT98), .C2(new_n648), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n296), .A2(new_n279), .A3(new_n297), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n287), .A3(G472), .ZN(new_n656));
  NAND2_X1  g470(.A1(G472), .A2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT96), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n293), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n308), .A2(new_n309), .ZN(new_n661));
  INV_X1    g475(.A(new_n188), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT32), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT97), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  OR3_X1    g478(.A1(new_n660), .A2(new_n663), .A3(KEYINPUT97), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n654), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n195), .ZN(G45));
  INV_X1    g481(.A(new_n608), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n449), .A2(new_n451), .ZN(new_n669));
  INV_X1    g483(.A(G475), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n429), .A2(new_n431), .A3(new_n418), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n671), .B2(new_n420), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n672), .B2(new_n432), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n668), .B(new_n638), .C1(new_n669), .C2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n640), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n311), .A2(new_n377), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  INV_X1    g491(.A(new_n577), .ZN(new_n678));
  INV_X1    g492(.A(G472), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n302), .B2(new_n305), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n662), .B1(new_n278), .B2(new_n292), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n681), .B2(new_n189), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n678), .B1(new_n682), .B2(new_n293), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n358), .A2(new_n363), .ZN(new_n684));
  OAI21_X1  g498(.A(G469), .B1(new_n684), .B2(G902), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n376), .A3(new_n364), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n609), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND3_X1  g505(.A1(new_n683), .A2(new_n617), .A3(new_n688), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NAND2_X1  g507(.A1(new_n482), .A2(new_n592), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n640), .A3(new_n686), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n311), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND4_X1  g511(.A1(new_n591), .A2(new_n453), .A3(new_n481), .A4(new_n592), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n687), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT100), .B(G472), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n581), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n291), .B1(new_n299), .B2(new_n257), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n662), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n577), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NOR3_X1   g520(.A1(new_n590), .A2(new_n674), .A3(new_n686), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n632), .A3(new_n701), .A4(new_n703), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  AND2_X1   g523(.A1(new_n535), .A2(new_n537), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n369), .A2(KEYINPUT101), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n362), .A2(new_n343), .A3(new_n712), .A4(new_n347), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n368), .A3(G469), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n364), .A3(new_n365), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n710), .A2(new_n715), .A3(new_n376), .A4(new_n490), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n674), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n661), .B2(new_n190), .ZN(new_n721));
  INV_X1    g535(.A(new_n190), .ZN(new_n722));
  AOI211_X1 g536(.A(KEYINPUT102), .B(new_n722), .C1(new_n308), .C2(new_n309), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n719), .B(new_n678), .C1(new_n724), .C2(new_n682), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n293), .A2(KEYINPUT102), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n661), .A2(new_n720), .A3(new_n190), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n682), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT103), .B1(new_n728), .B2(new_n577), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n718), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT42), .B1(new_n683), .B2(new_n717), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NOR2_X1   g548(.A1(new_n716), .A2(new_n639), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n311), .A2(new_n735), .A3(new_n577), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n311), .A2(new_n735), .A3(KEYINPUT104), .A4(new_n577), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NOR2_X1   g555(.A1(new_n453), .A2(new_n608), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT43), .B1(new_n453), .B2(new_n608), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n744), .A2(new_n632), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n582), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT44), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT106), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n711), .A2(new_n368), .A3(KEYINPUT45), .A4(new_n713), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n368), .A2(new_n369), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n750), .B(G469), .C1(new_n751), .C2(KEYINPUT45), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n365), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(KEYINPUT105), .A3(new_n364), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n752), .A2(new_n365), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n754), .B1(KEYINPUT46), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT105), .B1(new_n753), .B2(new_n364), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n376), .B(new_n650), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n535), .A2(new_n537), .A3(new_n490), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n746), .A2(new_n747), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n749), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT107), .B(G137), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G39));
  OAI21_X1  g581(.A(new_n376), .B1(new_n756), .B2(new_n757), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n376), .B(new_n769), .C1(new_n756), .C2(new_n757), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n311), .A2(new_n577), .A3(new_n674), .A4(new_n760), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  AND2_X1   g589(.A1(new_n665), .A2(new_n664), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n685), .A2(new_n364), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT49), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT109), .Z(new_n779));
  NOR3_X1   g593(.A1(new_n678), .A2(new_n375), .A3(new_n491), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(KEYINPUT49), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n647), .A2(new_n780), .A3(new_n742), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n776), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n744), .A2(new_n745), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n686), .A2(new_n760), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n485), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n632), .A3(new_n704), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n686), .A2(new_n678), .A3(new_n484), .A4(new_n760), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n776), .A2(new_n594), .A3(new_n608), .A4(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n577), .A2(new_n704), .A3(new_n485), .A4(new_n784), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n686), .A2(new_n490), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n647), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n788), .B(new_n790), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n710), .A3(new_n490), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n771), .A2(new_n772), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n685), .A2(new_n375), .A3(new_n364), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n776), .A2(new_n453), .A3(new_n668), .A4(new_n789), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n590), .A2(new_n686), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n791), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(G952), .A3(new_n345), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT113), .Z(new_n808));
  OAI21_X1  g622(.A(new_n798), .B1(new_n797), .B2(new_n802), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n307), .B1(new_n310), .B2(KEYINPUT32), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n721), .A3(new_n723), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n719), .B1(new_n811), .B2(new_n678), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n728), .A2(KEYINPUT103), .A3(new_n577), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n787), .ZN(new_n815));
  XOR2_X1   g629(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n803), .A2(new_n808), .A3(new_n809), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n731), .B1(new_n814), .B2(new_n718), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n689), .A2(new_n705), .A3(new_n692), .A4(new_n696), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT110), .B1(new_n594), .B2(new_n608), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n668), .B(new_n822), .C1(new_n669), .C2(new_n673), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n538), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n821), .A2(new_n538), .A3(new_n823), .A4(KEYINPUT111), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n538), .A2(new_n594), .A3(new_n481), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n585), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n578), .A2(new_n633), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n632), .A2(new_n480), .A3(new_n638), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n616), .A3(new_n760), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n311), .A2(new_n834), .A3(new_n377), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n717), .A2(new_n701), .A3(new_n632), .A4(new_n703), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n740), .A2(new_n831), .A3(new_n832), .A4(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n819), .A2(new_n820), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n453), .A2(new_n587), .A3(new_n589), .A4(new_n481), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n573), .A2(new_n629), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n715), .A2(new_n841), .A3(new_n376), .A4(new_n638), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n660), .B2(new_n663), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n642), .A2(new_n676), .A3(new_n708), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n838), .ZN(new_n849));
  INV_X1    g663(.A(new_n820), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n847), .A3(new_n733), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n819), .A2(new_n852), .A3(new_n820), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n838), .A2(KEYINPUT112), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n584), .B1(new_n828), .B2(new_n829), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n578), .A2(new_n633), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n740), .A4(new_n837), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(new_n847), .A3(new_n856), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n852), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n818), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n783), .B1(new_n867), .B2(new_n868), .ZN(G75));
  NOR2_X1   g683(.A1(new_n345), .A2(G952), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n847), .A2(new_n733), .A3(KEYINPUT53), .A4(new_n850), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n856), .A2(new_n861), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(G902), .B1(new_n848), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(G210), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n527), .A2(new_n529), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(new_n530), .Z(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT55), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n871), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n881), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT115), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n878), .A2(new_n885), .A3(new_n881), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n884), .B2(new_n886), .ZN(G51));
  NOR2_X1   g701(.A1(new_n876), .A2(new_n752), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT54), .B1(new_n848), .B2(new_n875), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n865), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n365), .B(KEYINPUT57), .Z(new_n891));
  AOI21_X1  g705(.A(new_n684), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n892), .B2(KEYINPUT116), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n894));
  INV_X1    g708(.A(new_n891), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n889), .B2(new_n865), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n896), .B2(new_n684), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n870), .B1(new_n893), .B2(new_n897), .ZN(G54));
  NOR2_X1   g712(.A1(new_n446), .A2(new_n447), .ZN(new_n899));
  NAND2_X1  g713(.A1(KEYINPUT58), .A2(G475), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n876), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n871), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n876), .A2(new_n899), .A3(new_n900), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(G60));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n854), .B2(new_n865), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n599), .A2(new_n601), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n871), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n890), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n912), .A2(KEYINPUT117), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(KEYINPUT117), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n862), .B2(new_n864), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n625), .A2(new_n628), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n870), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n565), .B(KEYINPUT119), .Z(new_n921));
  NOR2_X1   g735(.A1(new_n848), .A2(new_n875), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n917), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT61), .B1(new_n924), .B2(KEYINPUT118), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  AOI211_X1 g741(.A(new_n926), .B(new_n927), .C1(new_n920), .C2(new_n923), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n925), .A2(new_n928), .ZN(G66));
  INV_X1    g743(.A(G224), .ZN(new_n930));
  OAI21_X1  g744(.A(G953), .B1(new_n488), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT120), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n850), .A2(new_n859), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT121), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n879), .B1(G898), .B2(new_n345), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n936), .B(new_n937), .Z(G69));
  NAND2_X1  g752(.A1(new_n437), .A2(new_n438), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n251), .B(new_n939), .Z(new_n940));
  INV_X1    g754(.A(new_n840), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n814), .A2(new_n759), .A3(new_n941), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n733), .A2(new_n942), .A3(new_n740), .A4(new_n774), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n642), .A2(new_n708), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n676), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n765), .A2(KEYINPUT125), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT106), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n748), .B(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n759), .A3(new_n763), .ZN(new_n950));
  INV_X1    g764(.A(new_n945), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n943), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n953), .A2(new_n345), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n345), .A2(G900), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n940), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n821), .A2(new_n823), .B1(new_n594), .B2(new_n481), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n957), .A2(new_n651), .A3(new_n760), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n683), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n774), .B(new_n959), .C1(new_n749), .C2(new_n764), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n666), .A2(new_n945), .A3(KEYINPUT62), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT62), .B1(new_n666), .B2(new_n945), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT122), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(KEYINPUT62), .C1(new_n666), .C2(new_n945), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n962), .A2(new_n967), .A3(KEYINPUT123), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT123), .B1(new_n962), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n345), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n940), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n345), .B1(G227), .B2(G900), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT124), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n956), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n956), .B2(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G72));
  XNOR2_X1  g791(.A(new_n252), .B(KEYINPUT126), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n953), .A2(new_n933), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n657), .B(KEYINPUT63), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n279), .B(new_n979), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n304), .B2(new_n287), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n848), .B2(new_n853), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n871), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n979), .A2(new_n279), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n968), .A2(new_n969), .A3(new_n933), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n981), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(KEYINPUT127), .B(new_n986), .C1(new_n987), .C2(new_n981), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(G57));
endmodule


