//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  AND3_X1   g005(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT71), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT71), .A3(new_n210), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(KEYINPUT70), .B2(KEYINPUT28), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n215), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n228), .A2(new_n229), .B1(new_n230), .B2(new_n217), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n227), .B(new_n231), .C1(new_n229), .C2(new_n228), .ZN(new_n232));
  OAI22_X1  g031(.A1(new_n207), .A2(new_n208), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n233));
  INV_X1    g032(.A(G169gat), .ZN(new_n234));
  INV_X1    g033(.A(G176gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT25), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n228), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n230), .A2(new_n217), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT64), .A4(new_n228), .ZN(new_n245));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n235), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n248), .A2(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(KEYINPUT23), .A3(new_n235), .A4(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n242), .A2(new_n245), .A3(new_n252), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257));
  AOI221_X4 g056(.A(KEYINPUT69), .B1(new_n232), .B2(new_n238), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n257), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n232), .A2(new_n238), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n222), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(G127gat), .A2(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT72), .B(G127gat), .Z(new_n266));
  INV_X1    g065(.A(G134gat), .ZN(new_n267));
  OAI211_X1 g066(.A(KEYINPUT73), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n269));
  OR2_X1    g068(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n269), .B1(new_n272), .B2(new_n264), .ZN(new_n273));
  XOR2_X1   g072(.A(G113gat), .B(G120gat), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n268), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G120gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT74), .A3(G113gat), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  AND2_X1   g079(.A1(G127gat), .A2(G134gat), .ZN(new_n281));
  OAI221_X1 g080(.A(new_n280), .B1(new_n264), .B2(new_n281), .C1(new_n274), .C2(KEYINPUT74), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n283), .B(new_n222), .C1(new_n258), .C2(new_n262), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT32), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT33), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT75), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G15gat), .ZN(new_n295));
  INV_X1    g094(.A(G43gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n289), .B(KEYINPUT32), .C1(new_n291), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n287), .B1(new_n285), .B2(new_n288), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n304));
  OAI211_X1 g103(.A(KEYINPUT77), .B(KEYINPUT34), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n260), .A2(new_n261), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT69), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n256), .A2(new_n257), .B1(new_n232), .B2(new_n238), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n259), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n283), .B1(new_n311), .B2(new_n222), .ZN(new_n312));
  INV_X1    g111(.A(new_n288), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n286), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n306), .B1(new_n314), .B2(KEYINPUT76), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT34), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(new_n303), .B2(KEYINPUT77), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n305), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n202), .B1(new_n302), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n298), .A3(new_n300), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT77), .B1(new_n303), .B2(new_n304), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n306), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n301), .A2(new_n323), .A3(new_n305), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n319), .B1(new_n325), .B2(new_n202), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT35), .ZN(new_n327));
  XOR2_X1   g126(.A(G211gat), .B(G218gat), .Z(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n329), .A2(KEYINPUT80), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n329), .A2(KEYINPUT80), .B1(G211gat), .B2(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n330), .B2(new_n331), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(new_n331), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT81), .ZN(new_n339));
  INV_X1    g138(.A(new_n328), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n333), .A4(new_n334), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n219), .A2(new_n221), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n214), .B2(new_n213), .ZN(new_n344));
  INV_X1    g143(.A(G226gat), .ZN(new_n345));
  INV_X1    g144(.A(G233gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n344), .A2(new_n309), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(KEYINPUT29), .ZN(new_n350));
  AOI211_X1 g149(.A(new_n342), .B(new_n349), .C1(new_n263), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n342), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n347), .B(new_n222), .C1(new_n258), .C2(new_n262), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n350), .B1(new_n344), .B2(new_n309), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT82), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358));
  INV_X1    g157(.A(new_n349), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n344), .B1(new_n308), .B2(new_n310), .ZN(new_n360));
  INV_X1    g159(.A(new_n350), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n352), .B(new_n359), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n356), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n357), .A2(new_n362), .A3(new_n366), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n351), .A2(new_n355), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT30), .A3(new_n366), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G141gat), .B(G148gat), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n379), .A2(KEYINPUT2), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n388));
  INV_X1    g187(.A(G141gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(G148gat), .ZN(new_n390));
  INV_X1    g189(.A(G148gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT84), .A3(G141gat), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n390), .B(new_n392), .C1(G141gat), .C2(new_n391), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n379), .B1(new_n378), .B2(KEYINPUT2), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n384), .A2(new_n387), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n337), .B2(new_n341), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n397), .A2(KEYINPUT85), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n397), .B2(KEYINPUT85), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n395), .B2(new_n399), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(new_n352), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n393), .A2(new_n394), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n382), .A2(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n342), .A2(new_n412), .ZN(new_n413));
  OAI221_X1 g212(.A(new_n411), .B1(new_n404), .B2(new_n342), .C1(new_n413), .C2(new_n395), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n403), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G22gat), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n418), .B1(new_n407), .B2(new_n415), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(KEYINPUT86), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT86), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n395), .A2(new_n277), .A3(new_n282), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n395), .B1(new_n277), .B2(new_n282), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT5), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n431), .A2(KEYINPUT4), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n431), .A2(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n395), .A2(new_n399), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n283), .A3(new_n411), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n440), .B2(new_n430), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n431), .A2(KEYINPUT4), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n438), .A2(new_n283), .A3(new_n411), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n431), .A2(KEYINPUT4), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(KEYINPUT5), .A3(new_n429), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT0), .ZN(new_n449));
  XNOR2_X1  g248(.A(G57gat), .B(G85gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  AOI21_X1  g250(.A(KEYINPUT6), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n441), .A2(new_n453), .A3(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n441), .A2(new_n446), .A3(KEYINPUT89), .A4(new_n453), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n441), .A2(new_n446), .A3(KEYINPUT6), .A4(new_n453), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND4_X1   g259(.A1(new_n327), .A2(new_n375), .A3(new_n428), .A4(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n459), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n452), .B2(new_n454), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n374), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(new_n320), .A3(new_n324), .A4(new_n428), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n326), .A2(new_n461), .B1(new_n465), .B2(KEYINPUT35), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OR3_X1    g266(.A1(new_n432), .A2(new_n433), .A3(new_n430), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT39), .B(new_n468), .C1(new_n445), .C2(new_n429), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n440), .A2(new_n430), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n469), .B(new_n451), .C1(KEYINPUT39), .C2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n456), .A3(new_n457), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n366), .B1(new_n372), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n342), .B1(new_n353), .B2(new_n354), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT37), .B1(new_n480), .B2(new_n352), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(new_n459), .A3(new_n369), .A4(new_n458), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n356), .A2(new_n363), .A3(KEYINPUT37), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n478), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  OAI221_X1 g284(.A(new_n428), .B1(new_n475), .B2(new_n375), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n428), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n426), .A2(KEYINPUT87), .A3(new_n427), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n464), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT78), .B(KEYINPUT36), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT79), .B1(new_n320), .B2(new_n324), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n319), .ZN(new_n493));
  INV_X1    g292(.A(new_n325), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT36), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n486), .B1(new_n496), .B2(KEYINPUT88), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(new_n495), .ZN(new_n498));
  INV_X1    g297(.A(new_n490), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n498), .A2(KEYINPUT88), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n467), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G8gat), .ZN(new_n502));
  INV_X1    g301(.A(G1gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT16), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT92), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(G1gat), .B2(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI221_X1 g310(.A(new_n507), .B1(new_n508), .B2(new_n502), .C1(G1gat), .C2(new_n506), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n517), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n522), .A2(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  XOR2_X1   g323(.A(G43gat), .B(G50gat), .Z(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n525), .A2(new_n526), .B1(new_n521), .B2(new_n515), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n527), .B(new_n529), .C1(new_n519), .C2(new_n520), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n513), .B1(new_n514), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(KEYINPUT17), .A3(new_n530), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n532), .A2(new_n533), .B1(new_n513), .B2(new_n531), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT94), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G169gat), .B(G197gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT12), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n513), .B(new_n531), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n535), .B(KEYINPUT13), .Z(new_n547));
  AOI22_X1  g346(.A1(new_n536), .A2(new_n537), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n535), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n550), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n501), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n554), .A2(new_n463), .ZN(new_n555));
  INV_X1    g354(.A(new_n513), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT21), .ZN(new_n557));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n556), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT96), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n557), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G127gat), .B(G155gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT95), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n564), .A2(new_n570), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n571), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n531), .A2(new_n514), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n580), .A2(new_n533), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n531), .A2(new_n589), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT97), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n599), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n596), .B1(KEYINPUT97), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT98), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n562), .B1(new_n587), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n587), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT99), .B1(new_n609), .B2(KEYINPUT98), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n588), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT100), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n589), .A2(new_n562), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT101), .ZN(new_n616));
  INV_X1    g415(.A(new_n613), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT10), .B1(new_n611), .B2(new_n614), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n590), .A2(new_n562), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n616), .A2(new_n625), .A3(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n579), .A2(new_n604), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n555), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT102), .B(G1gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(G1324gat));
  NAND3_X1  g432(.A1(new_n554), .A2(new_n630), .A3(new_n374), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT42), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n634), .A2(new_n639), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n638), .B1(new_n642), .B2(new_n635), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n554), .A2(new_n374), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(KEYINPUT103), .A3(new_n630), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n634), .A2(new_n639), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(G8gat), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n643), .B1(new_n649), .B2(new_n650), .ZN(G1325gat));
  NAND2_X1  g450(.A1(new_n554), .A2(new_n630), .ZN(new_n652));
  OAI21_X1  g451(.A(G15gat), .B1(new_n652), .B2(new_n498), .ZN(new_n653));
  INV_X1    g452(.A(new_n326), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n652), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n488), .A2(new_n489), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n554), .A2(new_n630), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  NOR2_X1   g459(.A1(new_n578), .A2(new_n629), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n604), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n555), .A2(new_n519), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT45), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n498), .A2(new_n499), .A3(new_n486), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n467), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n604), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n670));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n663), .B1(new_n667), .B2(new_n467), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673));
  INV_X1    g472(.A(new_n670), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n501), .A2(new_n604), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n553), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n463), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n666), .A2(new_n684), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n644), .A2(new_n520), .A3(new_n664), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n682), .B2(new_n375), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  OAI21_X1  g489(.A(G43gat), .B1(new_n682), .B2(new_n498), .ZN(new_n691));
  INV_X1    g490(.A(new_n664), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G43gat), .A3(new_n654), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n554), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n691), .A2(KEYINPUT47), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1330gat));
  OAI21_X1  g498(.A(G50gat), .B1(new_n682), .B2(new_n428), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n692), .A2(G50gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n554), .A2(new_n657), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(KEYINPUT48), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n673), .B1(new_n672), .B2(new_n674), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n466), .B1(new_n496), .B2(new_n486), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n705), .A2(KEYINPUT106), .A3(new_n663), .A4(new_n670), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n501), .B2(new_n604), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n657), .B(new_n681), .C1(new_n707), .C2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n710), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT108), .B1(new_n710), .B2(G50gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n554), .A2(new_n714), .A3(new_n657), .A4(new_n701), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n711), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n703), .B1(new_n717), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g517(.A1(new_n680), .A2(new_n578), .A3(new_n663), .A4(new_n629), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT110), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n668), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n668), .A3(KEYINPUT111), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n683), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT112), .B(G57gat), .Z(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1332gat));
  INV_X1    g527(.A(new_n725), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n375), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n729), .B(new_n730), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT49), .ZN(new_n732));
  INV_X1    g531(.A(G64gat), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n732), .B(new_n733), .C1(new_n725), .C2(new_n375), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT113), .B(KEYINPUT114), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  XOR2_X1   g536(.A(new_n326), .B(KEYINPUT115), .Z(new_n738));
  AOI21_X1  g537(.A(G71gat), .B1(new_n729), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(G71gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n740), .A3(new_n498), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g542(.A1(new_n729), .A2(new_n657), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n553), .A2(new_n578), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n629), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n676), .B2(new_n678), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n683), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n672), .A2(new_n746), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n672), .A2(KEYINPUT51), .A3(new_n746), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n748), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n584), .A3(new_n463), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(G1336gat));
  NAND3_X1  g559(.A1(new_n679), .A2(new_n374), .A3(new_n749), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n375), .A2(G92gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n762), .A2(new_n764), .A3(new_n765), .A4(KEYINPUT52), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n585), .B1(new_n751), .B2(new_n374), .ZN(new_n769));
  INV_X1    g568(.A(new_n764), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n766), .A2(new_n771), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n752), .B2(new_n498), .ZN(new_n773));
  INV_X1    g572(.A(new_n758), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n654), .A2(G99gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(G1338gat));
  INV_X1    g575(.A(G106gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n751), .B2(new_n657), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n428), .A2(G106gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n758), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  INV_X1    g580(.A(new_n428), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n777), .B1(new_n751), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n784));
  INV_X1    g583(.A(new_n779), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(new_n786), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n680), .A2(G113gat), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n618), .A2(new_n617), .A3(new_n620), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n621), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n621), .A2(KEYINPUT54), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n791), .A2(KEYINPUT118), .A3(new_n626), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT118), .B1(new_n791), .B2(new_n626), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n790), .B(KEYINPUT55), .C1(new_n792), .C2(new_n793), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n796), .A2(new_n553), .A3(new_n628), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n534), .A2(new_n535), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n546), .A2(new_n547), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n543), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n548), .A2(new_n544), .A3(new_n549), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n629), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n604), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(new_n628), .A3(new_n797), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n604), .A2(new_n802), .A3(new_n801), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n579), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n630), .A2(new_n680), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n494), .A2(new_n428), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n463), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n374), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(KEYINPUT120), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(KEYINPUT120), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n788), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n657), .B1(new_n808), .B2(new_n809), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n683), .A2(new_n374), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n326), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n680), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n629), .A2(new_n278), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT121), .Z(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n819), .B2(new_n820), .ZN(new_n829));
  OAI21_X1  g628(.A(G120gat), .B1(new_n824), .B2(new_n748), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1341gat));
  NAND3_X1  g630(.A1(new_n818), .A2(new_n578), .A3(new_n266), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n824), .A2(new_n579), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n266), .B2(new_n833), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n604), .A2(new_n267), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n817), .A2(KEYINPUT56), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n824), .B2(new_n663), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT56), .B1(new_n817), .B2(new_n835), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(G1343gat));
  AOI21_X1  g638(.A(new_n428), .B1(new_n808), .B2(new_n809), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(KEYINPUT57), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n808), .A2(new_n809), .B1(new_n489), .B2(new_n488), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n841), .A2(new_n842), .B1(KEYINPUT57), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT122), .B1(new_n840), .B2(KEYINPUT57), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n498), .A2(new_n823), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n680), .A2(new_n389), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n498), .A2(new_n782), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n463), .A2(new_n810), .A3(new_n375), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(G141gat), .B1(new_n853), .B2(new_n553), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(KEYINPUT123), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n847), .B1(new_n844), .B2(new_n845), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n854), .B1(new_n859), .B2(new_n849), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT58), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(G1344gat));
  NAND3_X1  g662(.A1(new_n853), .A2(new_n391), .A3(new_n629), .ZN(new_n864));
  AOI211_X1 g663(.A(KEYINPUT59), .B(new_n391), .C1(new_n859), .C2(new_n629), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n840), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n843), .A2(new_n867), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n868), .A2(new_n629), .A3(new_n848), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n870), .B2(G148gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n864), .B1(new_n865), .B2(new_n871), .ZN(G1345gat));
  AOI21_X1  g671(.A(new_n376), .B1(new_n859), .B2(new_n578), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n853), .A2(new_n376), .A3(new_n578), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  AOI21_X1  g674(.A(G162gat), .B1(new_n853), .B2(new_n604), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n663), .A2(new_n377), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n859), .B2(new_n877), .ZN(G1347gat));
  AOI21_X1  g677(.A(new_n463), .B1(new_n808), .B2(new_n809), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(new_n374), .A3(new_n812), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n880), .A2(new_n553), .A3(new_n253), .A4(new_n254), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n375), .A2(new_n463), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n822), .A2(new_n738), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n680), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT124), .Z(G1348gat));
  NAND3_X1  g685(.A1(new_n880), .A2(new_n235), .A3(new_n629), .ZN(new_n887));
  OAI21_X1  g686(.A(G176gat), .B1(new_n883), .B2(new_n748), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n578), .A3(new_n216), .ZN(new_n890));
  OAI21_X1  g689(.A(G183gat), .B1(new_n883), .B2(new_n579), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g692(.A1(new_n880), .A2(new_n217), .A3(new_n604), .ZN(new_n894));
  OAI21_X1  g693(.A(G190gat), .B1(new_n883), .B2(new_n663), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1351gat));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n374), .A3(new_n852), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(G197gat), .B1(new_n900), .B2(new_n553), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n868), .A2(new_n869), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n498), .A2(new_n882), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n553), .A2(G197gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n901), .B1(new_n907), .B2(new_n908), .ZN(G1352gat));
  XNOR2_X1  g708(.A(KEYINPUT126), .B(G204gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n906), .B2(new_n748), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n899), .A2(new_n748), .A3(new_n910), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT62), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1353gat));
  NOR3_X1   g713(.A1(new_n899), .A2(G211gat), .A3(new_n579), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n868), .A2(new_n578), .A3(new_n869), .A4(new_n905), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT63), .B1(new_n916), .B2(G211gat), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n916), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1354gat));
  AOI21_X1  g721(.A(G218gat), .B1(new_n900), .B2(new_n604), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n604), .A2(G218gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n907), .B2(new_n924), .ZN(G1355gat));
endmodule


