//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1336, new_n1337, new_n1338, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n212), .B1(new_n216), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT7), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT7), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n258), .A3(new_n207), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(G68), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G58), .A2(G68), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(new_n201), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n262), .A2(G20), .B1(G159), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT16), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n214), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n261), .A2(new_n201), .ZN(new_n271));
  INV_X1    g0071(.A(G159), .ZN(new_n272));
  INV_X1    g0072(.A(new_n263), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n207), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n207), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n220), .B1(new_n277), .B2(KEYINPUT7), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n257), .A2(new_n213), .A3(new_n258), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n270), .B1(new_n280), .B2(KEYINPUT16), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n206), .A2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT8), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G58), .ZN(new_n288));
  INV_X1    g0088(.A(G58), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(KEYINPUT8), .ZN(new_n290));
  OAI211_X1 g0090(.A(KEYINPUT76), .B(new_n286), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n283), .A2(new_n214), .A3(new_n268), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n287), .A2(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT76), .B1(new_n296), .B2(new_n286), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n285), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT77), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT76), .ZN(new_n301));
  INV_X1    g0101(.A(new_n286), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n282), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(new_n292), .A3(new_n291), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n267), .A2(new_n281), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G1698), .ZN(new_n307));
  OAI211_X1 g0107(.A(G223), .B(new_n307), .C1(new_n255), .C2(new_n256), .ZN(new_n308));
  OAI211_X1 g0108(.A(G226), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G41), .ZN(new_n314));
  INV_X1    g0114(.A(G45), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n214), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G41), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n206), .A2(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G274), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n317), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n319), .A2(G232), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n313), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n313), .A2(KEYINPUT78), .A3(new_n324), .ZN(new_n328));
  AOI21_X1  g0128(.A(G200), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT79), .B(G190), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n306), .B(KEYINPUT17), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n313), .A2(KEYINPUT78), .A3(new_n324), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT78), .B1(new_n313), .B2(new_n324), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n331), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT17), .B1(new_n339), .B2(new_n306), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n213), .A2(G33), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n349), .A2(new_n213), .B1(new_n282), .B2(new_n273), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n269), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n292), .A2(G77), .A3(new_n286), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT72), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n284), .A2(new_n349), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n321), .A2(new_n323), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n317), .A2(new_n318), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n322), .ZN(new_n359));
  INV_X1    g0159(.A(G244), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(G1698), .B1(new_n275), .B2(new_n276), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G232), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n257), .A2(G107), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n361), .B1(new_n366), .B2(new_n312), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n367), .A2(G169), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n356), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n351), .A2(KEYINPUT73), .A3(new_n354), .A4(new_n355), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n312), .ZN(new_n373));
  INV_X1    g0173(.A(new_n361), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(G190), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n334), .B2(new_n367), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n356), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n371), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n325), .A2(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n327), .A2(new_n328), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n255), .A2(new_n256), .A3(G20), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n385), .B2(new_n258), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n257), .A2(new_n213), .A3(new_n258), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT16), .B(new_n264), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n269), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT16), .B1(new_n260), .B2(new_n264), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n304), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT77), .B1(new_n304), .B2(new_n285), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n389), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n380), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n383), .B1(new_n335), .B2(new_n336), .ZN(new_n395));
  INV_X1    g0195(.A(new_n381), .ZN(new_n396));
  AND4_X1   g0196(.A1(new_n380), .A2(new_n393), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n341), .A2(new_n379), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n286), .A2(G50), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n292), .A2(new_n401), .B1(new_n202), .B2(new_n284), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n347), .A2(KEYINPUT70), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT70), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n213), .A2(new_n404), .A3(G33), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n405), .A3(new_n296), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n263), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT9), .B(new_n402), .C1(new_n408), .C2(new_n270), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT9), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n270), .B1(new_n406), .B2(new_n407), .ZN(new_n411));
  INV_X1    g0211(.A(new_n402), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT10), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n253), .A2(G222), .A3(new_n307), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n253), .A2(G223), .A3(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n257), .A2(G77), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT69), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT69), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n416), .A2(new_n417), .A3(new_n421), .A4(new_n418), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n312), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G226), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n359), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n312), .A2(new_n320), .A3(new_n322), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT68), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT68), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n357), .B(new_n428), .C1(new_n359), .C2(new_n424), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n423), .A2(new_n430), .A3(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n423), .A2(new_n430), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n414), .A2(new_n415), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n433), .A2(new_n431), .A3(new_n409), .A4(new_n413), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT10), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n432), .A2(G179), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n411), .A2(new_n412), .ZN(new_n439));
  AOI21_X1  g0239(.A(G169), .B1(new_n423), .B2(new_n430), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT11), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n403), .A2(G77), .A3(new_n405), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n444), .B1(new_n447), .B2(new_n270), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n292), .A2(G68), .A3(new_n286), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT12), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n284), .B2(new_n220), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n270), .B1(new_n445), .B2(new_n446), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(KEYINPUT11), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT13), .ZN(new_n458));
  OAI211_X1 g0258(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT74), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT74), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n253), .A2(new_n461), .A3(G232), .A4(G1698), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n362), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n312), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n357), .B1(new_n359), .B2(new_n221), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n458), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n358), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n470), .A2(KEYINPUT13), .A3(new_n467), .ZN(new_n471));
  OAI211_X1 g0271(.A(G169), .B(new_n457), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n466), .A2(new_n458), .A3(new_n468), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT13), .B1(new_n470), .B2(new_n467), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(G179), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n474), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n457), .B1(new_n477), .B2(G169), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n456), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G190), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n469), .A2(new_n471), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n334), .B1(new_n473), .B2(new_n474), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n481), .A2(new_n482), .A3(new_n456), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n399), .A2(new_n443), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G250), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  OAI211_X1 g0288(.A(G244), .B(new_n307), .C1(new_n255), .C2(new_n256), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT4), .B1(new_n362), .B2(G244), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n312), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n206), .A2(G45), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n312), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(G257), .B1(new_n321), .B2(new_n498), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n383), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n258), .B1(new_n257), .B2(new_n213), .ZN(new_n503));
  NOR4_X1   g0303(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT7), .A4(G20), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n507));
  XNOR2_X1  g0307(.A(G97), .B(G107), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n510), .A2(new_n213), .B1(new_n349), .B2(new_n273), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n269), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n283), .A2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n206), .A2(G33), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n283), .A2(new_n514), .A3(new_n214), .A4(new_n268), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n493), .A2(new_n500), .A3(new_n368), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n502), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n501), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(new_n517), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n254), .A2(G107), .A3(new_n259), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n273), .A2(new_n349), .ZN(new_n524));
  AND2_X1   g0324(.A1(G97), .A2(G107), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G97), .A2(G107), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n509), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n524), .B1(new_n529), .B2(new_n252), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n522), .B1(new_n531), .B2(new_n269), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n493), .A2(new_n500), .A3(G190), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n521), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n520), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n253), .A2(KEYINPUT81), .A3(G244), .A4(G1698), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n253), .A2(G238), .A3(new_n307), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n312), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n223), .B1(new_n206), .B2(G45), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT80), .B1(new_n358), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n358), .A2(new_n544), .A3(KEYINPUT80), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n315), .A2(G1), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n546), .A2(new_n547), .B1(new_n321), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n543), .A2(G179), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n383), .B1(new_n543), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT82), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n543), .A2(new_n549), .A3(G179), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT82), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n321), .A2(new_n548), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n358), .A2(new_n544), .A3(KEYINPUT80), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(new_n545), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n312), .B2(new_n542), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n553), .B(new_n554), .C1(new_n558), .C2(new_n383), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n249), .A2(new_n251), .A3(G33), .A4(G97), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n213), .A2(new_n253), .A3(G68), .ZN(new_n563));
  NAND3_X1  g0363(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n249), .A2(new_n251), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n526), .A2(new_n222), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n269), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n346), .A2(new_n284), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n344), .A2(new_n345), .A3(new_n516), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT83), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT83), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n569), .A2(new_n574), .A3(new_n570), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n552), .A2(new_n559), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n516), .A2(G87), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n569), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(G190), .B2(new_n558), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n543), .A2(new_n549), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n535), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n249), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT22), .B1(new_n585), .B2(new_n222), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n213), .A2(new_n253), .A3(new_n587), .A4(G87), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND2_X1  g0390(.A1(KEYINPUT23), .A2(G107), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(G20), .ZN(new_n593));
  NOR2_X1   g0393(.A1(KEYINPUT23), .A2(G107), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n252), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n589), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n590), .B1(new_n589), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n269), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT25), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n283), .B2(G107), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n283), .A2(new_n599), .A3(G107), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n601), .A2(new_n602), .B1(new_n505), .B2(new_n515), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n498), .A2(new_n321), .ZN(new_n607));
  INV_X1    g0407(.A(new_n497), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n548), .B1(new_n608), .B2(new_n495), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(G264), .A3(new_n358), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G250), .A2(G1698), .ZN(new_n611));
  INV_X1    g0411(.A(G257), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(G1698), .ZN(new_n613));
  INV_X1    g0413(.A(G294), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT86), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT86), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G294), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n613), .A2(new_n253), .B1(new_n618), .B2(G33), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n607), .B(new_n610), .C1(new_n619), .C2(new_n358), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n612), .A2(G1698), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(G250), .B2(G1698), .ZN(new_n623));
  XNOR2_X1  g0423(.A(KEYINPUT86), .B(G294), .ZN(new_n624));
  INV_X1    g0424(.A(G33), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n623), .A2(new_n257), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n312), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n607), .A4(new_n610), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(G169), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n620), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G179), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n605), .A2(new_n606), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n606), .B1(new_n605), .B2(new_n633), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n620), .A2(new_n334), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n621), .A2(new_n629), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n480), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n605), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n641));
  OAI211_X1 g0441(.A(G257), .B(new_n307), .C1(new_n255), .C2(new_n256), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n312), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n609), .A2(G270), .A3(new_n358), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n607), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(G169), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n515), .A2(G116), .ZN(new_n649));
  INV_X1    g0449(.A(G116), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n283), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n625), .A2(G97), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n249), .A2(new_n251), .A3(new_n653), .A4(new_n488), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n268), .A2(new_n214), .B1(G20), .B2(new_n650), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n654), .A2(KEYINPUT20), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT20), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT84), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n652), .B(KEYINPUT84), .C1(new_n656), .C2(new_n657), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n648), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  INV_X1    g0465(.A(new_n647), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n644), .A2(new_n312), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n368), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n662), .A2(new_n664), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n648), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n664), .B1(new_n665), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n645), .A2(new_n647), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(G200), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n660), .A4(new_n661), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n670), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AND4_X1   g0479(.A1(new_n486), .A2(new_n584), .A3(new_n640), .A4(new_n679), .ZN(G372));
  NAND2_X1  g0480(.A1(new_n484), .A2(new_n371), .ZN(new_n681));
  AOI211_X1 g0481(.A(new_n340), .B(new_n333), .C1(new_n681), .C2(new_n479), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT90), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n394), .B2(new_n397), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT18), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n384), .A2(new_n380), .A3(new_n393), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT90), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n437), .B1(new_n682), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(new_n442), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n589), .A2(new_n595), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT24), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n589), .A2(new_n590), .A3(new_n595), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n603), .B1(new_n696), .B2(new_n269), .ZN(new_n697));
  AOI21_X1  g0497(.A(G190), .B1(new_n621), .B2(new_n629), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n636), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n553), .B1(new_n558), .B2(new_n383), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n700), .A2(new_n576), .B1(new_n580), .B2(new_n582), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n701), .A3(new_n535), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n665), .A2(new_n671), .A3(new_n664), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n665), .A2(new_n669), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n598), .A2(new_n604), .B1(new_n630), .B2(new_n632), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n706), .A3(new_n672), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n692), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n520), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n577), .A2(new_n709), .A3(new_n583), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT26), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n576), .A2(new_n700), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT26), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n709), .A3(new_n583), .A4(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(new_n712), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n520), .A2(new_n534), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n639), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n605), .A2(new_n633), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n670), .A2(new_n718), .A3(new_n673), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(new_n719), .A3(KEYINPUT89), .A4(new_n701), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n708), .A2(new_n711), .A3(new_n715), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n486), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n691), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT91), .ZN(G369));
  NAND3_X1  g0524(.A1(new_n213), .A2(new_n206), .A3(G13), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G213), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G343), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n665), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n679), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n705), .A2(new_n672), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(new_n731), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  INV_X1    g0535(.A(new_n633), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT88), .B1(new_n736), .B2(new_n697), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n706), .A2(new_n606), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n699), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n730), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n697), .A2(new_n740), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n739), .A2(new_n741), .B1(new_n718), .B2(new_n740), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n733), .A2(new_n730), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n640), .A2(new_n745), .B1(new_n706), .B2(new_n740), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(G399));
  INV_X1    g0547(.A(new_n210), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G41), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n206), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n526), .A2(new_n222), .A3(new_n650), .ZN(new_n752));
  INV_X1    g0552(.A(new_n749), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n751), .A2(new_n752), .B1(new_n218), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT28), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n712), .A2(new_n583), .ZN(new_n756));
  OAI21_X1  g0556(.A(KEYINPUT26), .B1(new_n756), .B2(new_n520), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n577), .A2(new_n713), .A3(new_n709), .A4(new_n583), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n757), .A2(new_n758), .A3(new_n712), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n634), .A2(new_n635), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n733), .ZN(new_n761));
  INV_X1    g0561(.A(new_n702), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n759), .A2(KEYINPUT93), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT93), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n757), .A2(new_n758), .A3(new_n764), .A4(new_n712), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n730), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT29), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n721), .A2(new_n740), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(KEYINPUT29), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n640), .A2(new_n584), .A3(new_n679), .A4(new_n740), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT92), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT30), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n558), .A2(new_n674), .A3(G179), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n493), .A2(new_n500), .A3(new_n610), .A4(new_n627), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n776), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n778), .A2(new_n669), .A3(KEYINPUT30), .A4(new_n558), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n631), .A2(G179), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n780), .A2(new_n501), .A3(new_n581), .A4(new_n668), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n782), .A2(KEYINPUT31), .A3(new_n730), .ZN(new_n783));
  AOI21_X1  g0583(.A(KEYINPUT31), .B1(new_n782), .B2(new_n730), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n773), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(new_n730), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT31), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n782), .A2(KEYINPUT31), .A3(new_n730), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n788), .A2(KEYINPUT92), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n772), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G330), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n771), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n755), .B1(new_n794), .B2(G1), .ZN(G364));
  AND2_X1   g0595(.A1(new_n213), .A2(G13), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G45), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n750), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n748), .A2(new_n257), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n650), .B2(new_n748), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n244), .A2(new_n315), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n748), .A2(new_n253), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G45), .B2(new_n218), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n800), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n214), .B1(G20), .B2(new_n383), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n798), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n807), .B(KEYINPUT100), .Z(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n213), .A2(new_n368), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT94), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(new_n480), .A3(new_n334), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n480), .A3(G200), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  OAI22_X1  g0617(.A1(new_n812), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n207), .A2(new_n480), .A3(new_n334), .A4(G179), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n253), .B1(new_n819), .B2(G303), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G179), .A2(G200), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n252), .B1(new_n480), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n213), .A2(KEYINPUT97), .A3(G190), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT97), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n252), .B2(new_n480), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n828), .A2(G179), .A3(new_n334), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n820), .B1(new_n624), .B2(new_n824), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n828), .A2(new_n822), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n818), .B(new_n832), .C1(G329), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G322), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n814), .A2(new_n334), .A3(new_n330), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT95), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G326), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n814), .A2(G200), .A3(new_n330), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT98), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n834), .B1(new_n835), .B2(new_n840), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT99), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n833), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n272), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT32), .ZN(new_n849));
  INV_X1    g0649(.A(new_n815), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n848), .A2(new_n849), .B1(new_n850), .B2(G77), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n851), .B1(new_n202), .B2(new_n842), .C1(new_n220), .C2(new_n816), .ZN(new_n852));
  INV_X1    g0652(.A(G97), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n824), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n819), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n222), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n854), .A2(new_n856), .A3(new_n257), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n857), .B1(new_n505), .B2(new_n830), .C1(new_n848), .C2(new_n849), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n840), .B(KEYINPUT96), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n289), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n844), .A2(new_n845), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n846), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n808), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n810), .B1(new_n734), .B2(new_n811), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n798), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n735), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(G330), .B2(new_n734), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G396));
  NAND2_X1  g0670(.A1(new_n371), .A2(new_n740), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n378), .A2(new_n372), .B1(new_n356), .B2(new_n730), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n371), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n769), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n873), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n721), .A2(new_n740), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n798), .B1(new_n879), .B2(new_n792), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n792), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(KEYINPUT104), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n881), .A2(KEYINPUT104), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n808), .A2(new_n805), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n798), .B1(new_n349), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n877), .B2(new_n806), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n829), .A2(G68), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n833), .A2(G132), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n253), .B1(new_n855), .B2(new_n202), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(G58), .B2(new_n823), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n842), .ZN(new_n893));
  AOI22_X1  g0693(.A1(G137), .A2(new_n893), .B1(new_n850), .B2(G159), .ZN(new_n894));
  INV_X1    g0694(.A(G150), .ZN(new_n895));
  INV_X1    g0695(.A(G143), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n894), .B1(new_n895), .B2(new_n816), .C1(new_n860), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT102), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT34), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n892), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n253), .B(new_n854), .C1(G107), .C2(new_n819), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n829), .A2(G87), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n902), .B(new_n903), .C1(new_n812), .C2(new_n847), .ZN(new_n904));
  AOI22_X1  g0704(.A1(G303), .A2(new_n893), .B1(new_n850), .B2(G116), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n831), .B2(new_n816), .ZN(new_n906));
  INV_X1    g0706(.A(new_n840), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n904), .B(new_n906), .C1(G294), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT101), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n887), .B1(new_n910), .B2(new_n808), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n884), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(G384));
  OR2_X1    g0713(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n914), .A2(new_n915), .A3(G116), .A4(new_n215), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT36), .Z(new_n917));
  OR3_X1    g0717(.A1(new_n218), .A2(new_n349), .A3(new_n261), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n202), .A2(G68), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n206), .B(G13), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n486), .B1(new_n768), .B2(new_n770), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n691), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n685), .A2(KEYINPUT106), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT37), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n306), .B1(new_n329), .B2(new_n331), .ZN(new_n928));
  INV_X1    g0728(.A(new_n728), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n393), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n928), .B(new_n930), .C1(new_n685), .C2(KEYINPUT106), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n298), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n280), .A2(KEYINPUT16), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n933), .B1(new_n389), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n395), .A3(new_n396), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT105), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n928), .A2(new_n936), .A3(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n929), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n932), .B1(new_n942), .B2(KEYINPUT37), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT38), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n341), .B2(new_n398), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n684), .A2(new_n341), .A3(new_n688), .ZN(new_n947));
  INV_X1    g0747(.A(new_n930), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n927), .A2(new_n931), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n928), .A2(new_n685), .A3(new_n930), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT37), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT38), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n924), .B1(new_n946), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(G169), .B1(new_n469), .B2(new_n471), .ZN(new_n956));
  INV_X1    g0756(.A(new_n457), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n475), .A3(new_n472), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(new_n456), .A3(new_n740), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n940), .A2(new_n941), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT105), .B1(new_n928), .B2(new_n936), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT37), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n950), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n341), .A2(new_n398), .ZN(new_n967));
  INV_X1    g0767(.A(new_n941), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(KEYINPUT38), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(KEYINPUT39), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n955), .A2(new_n961), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n456), .A2(new_n730), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n479), .A2(new_n484), .A3(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n456), .B(new_n730), .C1(new_n959), .C2(new_n483), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n878), .B2(new_n871), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n962), .A2(new_n970), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n689), .A2(new_n728), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n972), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n923), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G330), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n947), .A2(new_n948), .B1(new_n950), .B2(new_n952), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n970), .B1(new_n985), .B2(KEYINPUT38), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n783), .A2(new_n784), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n772), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n873), .B1(new_n974), .B2(new_n975), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT40), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n988), .A2(new_n993), .A3(new_n989), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n992), .A2(KEYINPUT40), .B1(new_n979), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n486), .A2(new_n988), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n984), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n996), .B2(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n983), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n206), .B2(new_n796), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n983), .A2(new_n998), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n921), .B1(new_n1000), .B2(new_n1001), .ZN(G367));
  NAND2_X1  g0802(.A1(new_n640), .A2(new_n745), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n535), .B1(new_n532), .B2(new_n740), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n520), .B2(new_n740), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT42), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n520), .B1(new_n760), .B2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n740), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(KEYINPUT42), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT108), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n730), .A2(new_n579), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n756), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n576), .A2(new_n1014), .A3(new_n700), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(new_n1018), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1019), .B1(new_n1022), .B2(new_n1013), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n743), .A2(new_n1006), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n749), .B(KEYINPUT41), .Z(new_n1026));
  NOR2_X1   g0826(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n746), .A2(new_n1006), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT45), .Z(new_n1029));
  NOR2_X1   g0829(.A1(new_n746), .A2(new_n1006), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT44), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1027), .B(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n742), .A2(new_n745), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT110), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1004), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1003), .A2(KEYINPUT110), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n1036), .A2(new_n735), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n735), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n794), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1026), .B1(new_n1042), .B2(new_n794), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n797), .A2(G1), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1025), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n202), .A2(new_n815), .B1(new_n816), .B2(new_n272), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n824), .A2(new_n220), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n257), .B(new_n1048), .C1(G58), .C2(new_n819), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n829), .A2(G77), .ZN(new_n1050));
  INV_X1    g0850(.A(G137), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1050), .C1(new_n1051), .C2(new_n847), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n843), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1047), .B(new_n1052), .C1(new_n1053), .C2(G143), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n895), .B2(new_n840), .ZN(new_n1055));
  INV_X1    g0855(.A(G303), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n860), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT46), .B1(new_n819), .B2(G116), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n819), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n257), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(G107), .C2(new_n823), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n829), .A2(G97), .ZN(new_n1062));
  INV_X1    g0862(.A(G317), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1062), .C1(new_n1063), .C2(new_n847), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n831), .A2(new_n815), .B1(new_n816), .B2(new_n624), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n812), .B2(new_n843), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1055), .B1(new_n1057), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT47), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n864), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n234), .A2(new_n802), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n809), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n346), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n748), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n798), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1071), .B(new_n1076), .C1(new_n811), .C2(new_n1020), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1046), .A2(new_n1077), .ZN(G387));
  NAND2_X1  g0878(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1056), .A2(new_n815), .B1(new_n816), .B2(new_n812), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1053), .B2(G322), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n860), .B2(new_n1063), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT48), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(KEYINPUT48), .B(new_n1082), .C1(new_n860), .C2(new_n1063), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n823), .A2(G283), .B1(new_n819), .B2(new_n618), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1080), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(KEYINPUT49), .A3(new_n1089), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n257), .B1(new_n847), .B2(new_n841), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G116), .B2(new_n829), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n346), .A2(new_n824), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n907), .B2(G50), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT113), .Z(new_n1100));
  AOI21_X1  g0900(.A(new_n257), .B1(new_n819), .B2(G77), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1062), .B(new_n1101), .C1(new_n895), .C2(new_n847), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT112), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n850), .A2(G68), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n816), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1105), .A2(new_n296), .B1(new_n893), .B2(G159), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n864), .B1(new_n1097), .B2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n799), .A2(new_n752), .B1(new_n505), .B2(new_n748), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n239), .A2(new_n315), .ZN(new_n1110));
  AOI211_X1 g0910(.A(G45), .B(new_n752), .C1(G68), .C2(G77), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT50), .B1(new_n296), .B2(new_n202), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n296), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n802), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1109), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n798), .B1(new_n1116), .B2(new_n809), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n742), .B2(new_n811), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1041), .A2(new_n749), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n794), .A2(new_n1040), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1079), .B1(new_n1108), .B2(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(G393));
  XNOR2_X1  g0921(.A(new_n1032), .B(new_n743), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1041), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1042), .A2(new_n749), .A3(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n840), .A2(new_n272), .B1(new_n895), .B2(new_n842), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT51), .Z(new_n1126));
  AOI21_X1  g0926(.A(new_n257), .B1(new_n819), .B2(G68), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n903), .B(new_n1127), .C1(new_n896), .C2(new_n847), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT115), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n850), .A2(new_n296), .B1(G77), .B2(new_n823), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n202), .B2(new_n816), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1126), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n840), .A2(new_n812), .B1(new_n1063), .B2(new_n842), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT52), .Z(new_n1134));
  OAI21_X1  g0934(.A(new_n257), .B1(new_n855), .B2(new_n831), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G116), .B2(new_n823), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n847), .B2(new_n835), .C1(new_n830), .C2(new_n505), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n614), .A2(new_n815), .B1(new_n816), .B2(new_n1056), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n808), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1005), .B(new_n807), .C1(new_n520), .C2(new_n740), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n802), .A2(new_n247), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1073), .B1(G97), .B2(new_n748), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n798), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1122), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n1045), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1124), .A2(new_n1147), .ZN(G390));
  INV_X1    g0948(.A(KEYINPUT118), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n535), .A2(new_n577), .A3(new_n583), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n739), .A2(new_n1150), .A3(new_n678), .A4(new_n730), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n788), .A2(new_n789), .ZN(new_n1152));
  OAI21_X1  g0952(.A(G330), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n875), .B1(new_n1153), .B2(KEYINPUT117), .ZN(new_n1154));
  AOI211_X1 g0954(.A(KEYINPUT117), .B(new_n984), .C1(new_n772), .C2(new_n987), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n976), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n759), .A2(KEYINPUT93), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n761), .A2(new_n762), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n765), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n872), .A2(new_n371), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n740), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n791), .A2(G330), .A3(new_n877), .A4(new_n976), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1163), .A3(new_n871), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1149), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n873), .B(KEYINPUT103), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n984), .B1(new_n772), .B2(new_n987), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT117), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n977), .B1(new_n1169), .B2(new_n1155), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n766), .A2(new_n1161), .B1(new_n371), .B2(new_n740), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1170), .A2(KEYINPUT118), .A3(new_n1171), .A4(new_n1163), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n977), .B1(new_n792), .B2(new_n873), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1167), .A2(new_n989), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n878), .A2(new_n871), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1165), .A2(new_n1172), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1167), .A2(new_n486), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT116), .Z(new_n1180));
  AND3_X1   g0980(.A1(new_n1180), .A2(new_n691), .A3(new_n922), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT119), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1174), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1176), .A2(new_n976), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1185), .A2(new_n960), .B1(new_n955), .B2(new_n971), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n960), .B1(new_n946), .B2(new_n954), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1162), .A2(new_n871), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n976), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1184), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n971), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n949), .A2(new_n953), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n944), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT39), .B1(new_n1193), .B2(new_n970), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n1191), .A2(new_n1194), .B1(new_n978), .B2(new_n961), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1171), .A2(new_n977), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1163), .C1(new_n1196), .C2(new_n1187), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n753), .B1(new_n1183), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1182), .A2(KEYINPUT119), .A3(new_n1198), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n805), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n819), .A2(G150), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT53), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n257), .B(new_n1205), .C1(G159), .C2(new_n823), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n833), .A2(G125), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n202), .C2(new_n830), .ZN(new_n1208));
  XOR2_X1   g1008(.A(KEYINPUT54), .B(G143), .Z(new_n1209));
  AOI22_X1  g1009(.A1(G128), .A2(new_n893), .B1(new_n850), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1051), .B2(new_n816), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(G132), .C2(new_n907), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n253), .B(new_n856), .C1(G77), .C2(new_n823), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n888), .C1(new_n614), .C2(new_n847), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G107), .A2(new_n1105), .B1(new_n850), .B2(G97), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n831), .B2(new_n842), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(G116), .C2(new_n907), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n864), .B1(new_n1218), .B2(KEYINPUT120), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(KEYINPUT120), .B2(new_n1218), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n798), .B1(new_n282), .B2(new_n885), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1203), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1045), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1198), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT121), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1224), .A2(KEYINPUT121), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1202), .A2(new_n1225), .A3(new_n1226), .ZN(G378));
  NOR2_X1   g1027(.A1(new_n439), .A2(new_n728), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n443), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n441), .B1(new_n434), .B2(new_n436), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1228), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1233), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n441), .B(new_n1228), .C1(new_n434), .C2(new_n436), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1234), .A2(new_n1238), .A3(KEYINPUT122), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT122), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n993), .B1(new_n986), .B2(new_n991), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n988), .A2(new_n989), .A3(new_n993), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n970), .B2(new_n962), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1241), .B(G330), .C1(new_n1242), .C2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n979), .A2(new_n994), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n990), .B1(new_n1193), .B2(new_n970), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n993), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1247), .B1(new_n1250), .B2(G330), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n982), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1247), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n995), .B2(new_n984), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n982), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1245), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1256), .A3(KEYINPUT123), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1255), .A3(new_n1258), .A4(new_n1245), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1045), .A3(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1241), .A2(new_n806), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n830), .A2(new_n289), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n847), .A2(new_n831), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n314), .B(new_n257), .C1(new_n855), .C2(new_n349), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1048), .A4(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n853), .A2(new_n816), .B1(new_n815), .B2(new_n346), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G116), .B2(new_n893), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1265), .B(new_n1267), .C1(new_n505), .C2(new_n840), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT58), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n257), .A2(new_n314), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G50), .B1(new_n625), .B2(new_n314), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1268), .A2(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n893), .A2(G125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n850), .A2(G137), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1105), .A2(G132), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n823), .A2(G150), .B1(new_n819), .B2(new_n1209), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n907), .B2(G128), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT59), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n625), .B(new_n314), .C1(new_n830), .C2(new_n272), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G124), .B2(new_n833), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT59), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1278), .B2(new_n1283), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1272), .B1(new_n1269), .B2(new_n1268), .C1(new_n1280), .C2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n808), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n798), .B1(new_n202), .B2(new_n885), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1261), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1260), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1178), .A2(new_n1197), .A3(new_n1190), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1181), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1294), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT57), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n753), .B1(new_n1297), .B2(new_n1294), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1295), .A2(KEYINPUT57), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1292), .B1(new_n1300), .B2(new_n1301), .ZN(G375));
  NOR3_X1   g1102(.A1(new_n808), .A2(G68), .A3(new_n805), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n253), .B(new_n1098), .C1(G97), .C2(new_n819), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1050), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(G303), .B2(new_n833), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n505), .A2(new_n815), .B1(new_n842), .B2(new_n614), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(G116), .B2(new_n1105), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1306), .B(new_n1308), .C1(new_n831), .C2(new_n840), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n860), .A2(new_n1051), .ZN(new_n1310));
  OAI221_X1 g1110(.A(new_n253), .B1(new_n855), .B2(new_n272), .C1(new_n824), .C2(new_n202), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1311), .B(new_n1262), .C1(G128), .C2(new_n833), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1105), .A2(new_n1209), .B1(new_n893), .B2(G132), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1312), .B(new_n1313), .C1(new_n895), .C2(new_n815), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1309), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n798), .B(new_n1303), .C1(new_n1315), .C2(new_n808), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n977), .A2(new_n805), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1178), .B2(new_n1045), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(KEYINPUT125), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1170), .A2(new_n1163), .A3(new_n1171), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1322), .A2(new_n1149), .B1(new_n1176), .B2(new_n1175), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1180), .A2(new_n922), .A3(new_n691), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1172), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1026), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1182), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1321), .A2(new_n1327), .ZN(G381));
  OR2_X1    g1128(.A1(G393), .A2(G396), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1124), .A2(new_n912), .A3(new_n1147), .ZN(new_n1330));
  NOR4_X1   g1130(.A1(G387), .A2(G381), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(G375), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1224), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  XOR2_X1   g1134(.A(new_n1334), .B(KEYINPUT126), .Z(G407));
  INV_X1    g1135(.A(G213), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1333), .A2(new_n729), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1332), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G407), .A2(new_n1338), .ZN(G409));
  XNOR2_X1  g1139(.A(G393), .B(new_n869), .ZN(new_n1340));
  OR2_X1    g1140(.A1(new_n1340), .A2(G390), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(G390), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(G387), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1343), .B(new_n1344), .ZN(new_n1345));
  OAI211_X1 g1145(.A(G378), .B(new_n1292), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1295), .A2(new_n1326), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1289), .B1(new_n1348), .B2(new_n1045), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1333), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1346), .A2(new_n1351), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1336), .A2(G343), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1323), .A2(KEYINPUT60), .A3(new_n1172), .A4(new_n1324), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n749), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1182), .A2(KEYINPUT60), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1357), .B1(new_n1325), .B2(new_n1358), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1320), .A2(KEYINPUT125), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT125), .ZN(new_n1361));
  AOI211_X1 g1161(.A(new_n1361), .B(new_n1319), .C1(new_n1178), .C2(new_n1045), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1360), .A2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n912), .B1(new_n1359), .B2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1358), .A2(new_n1325), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1365), .A2(new_n749), .A3(new_n1356), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1366), .A2(new_n1321), .A3(G384), .ZN(new_n1367));
  OR2_X1    g1167(.A1(new_n1354), .A2(KEYINPUT127), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1364), .A2(new_n1367), .A3(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1353), .A2(G2897), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1364), .A2(new_n1367), .A3(new_n1370), .A4(new_n1368), .ZN(new_n1373));
  AND2_X1   g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(KEYINPUT61), .B1(new_n1355), .B2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT63), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1364), .A2(new_n1367), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1376), .B1(new_n1355), .B2(new_n1377), .ZN(new_n1378));
  AOI21_X1  g1178(.A(new_n1353), .B1(new_n1346), .B2(new_n1351), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1377), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1379), .A2(KEYINPUT63), .A3(new_n1380), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1345), .A2(new_n1375), .A3(new_n1378), .A4(new_n1381), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT62), .ZN(new_n1383));
  AND3_X1   g1183(.A1(new_n1379), .A2(new_n1383), .A3(new_n1380), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT61), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1385), .B1(new_n1379), .B2(new_n1386), .ZN(new_n1387));
  AOI21_X1  g1187(.A(new_n1383), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1388));
  NOR3_X1   g1188(.A1(new_n1384), .A2(new_n1387), .A3(new_n1388), .ZN(new_n1389));
  OAI21_X1  g1189(.A(new_n1382), .B1(new_n1389), .B2(new_n1345), .ZN(G405));
  NAND2_X1  g1190(.A1(G375), .A2(new_n1333), .ZN(new_n1391));
  NAND3_X1  g1191(.A1(new_n1391), .A2(new_n1377), .A3(new_n1346), .ZN(new_n1392));
  INV_X1    g1192(.A(new_n1392), .ZN(new_n1393));
  AOI21_X1  g1193(.A(new_n1377), .B1(new_n1391), .B2(new_n1346), .ZN(new_n1394));
  NOR2_X1   g1194(.A1(new_n1393), .A2(new_n1394), .ZN(new_n1395));
  XNOR2_X1  g1195(.A(new_n1395), .B(new_n1345), .ZN(G402));
endmodule


