//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n214), .B1(new_n215), .B2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G13), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n217), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(G250), .B1(G257), .B2(G264), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n213), .B1(new_n222), .B2(KEYINPUT0), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n203), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G107), .A2(G264), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n215), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n223), .B(new_n232), .C1(KEYINPUT0), .C2(new_n222), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AOI21_X1  g0049(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT67), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(G222), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n250), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n265), .B(KEYINPUT66), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n250), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n269), .B2(G226), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G190), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n210), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n204), .A2(KEYINPUT68), .A3(G20), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G150), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT8), .B(G58), .Z(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n211), .A2(G33), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n275), .B(new_n277), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT68), .B1(new_n204), .B2(G20), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n274), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n217), .A2(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n201), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n274), .B1(new_n264), .B2(G20), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n201), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT9), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT70), .B1(new_n271), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n263), .A2(new_n270), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(G200), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n291), .A2(new_n293), .A3(new_n294), .A4(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n293), .A2(new_n297), .A3(new_n272), .A4(new_n290), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n295), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n289), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n284), .A2(G20), .A3(new_n203), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(KEYINPUT12), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(KEYINPUT12), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(KEYINPUT71), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(KEYINPUT71), .B2(new_n309), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT11), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n261), .B2(new_n280), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n274), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n311), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n312), .ZN(new_n317));
  INV_X1    g0117(.A(new_n287), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n203), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n267), .B1(new_n269), .B2(G238), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(new_n237), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n255), .A2(G226), .A3(new_n259), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n250), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n323), .B(new_n324), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n329), .B2(new_n330), .ZN(new_n334));
  INV_X1    g0134(.A(new_n267), .ZN(new_n335));
  INV_X1    g0135(.A(G41), .ZN(new_n336));
  INV_X1    g0136(.A(G45), .ZN(new_n337));
  AOI21_X1  g0137(.A(G1), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n332), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G238), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT13), .B1(new_n334), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n322), .B1(new_n333), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n333), .A2(G179), .A3(new_n344), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n345), .B2(new_n346), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n321), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n333), .A2(new_n344), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n292), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n333), .A2(new_n354), .A3(new_n344), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n321), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n285), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n278), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n318), .B2(new_n278), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n327), .A2(new_n259), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n255), .A2(G223), .A3(new_n259), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n332), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n335), .B1(new_n341), .B2(new_n237), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n292), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n267), .B1(new_n269), .B2(G232), .ZN(new_n369));
  INV_X1    g0169(.A(G226), .ZN(new_n370));
  INV_X1    g0170(.A(G87), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n256), .A2(new_n370), .B1(new_n252), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n365), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n250), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n354), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n255), .B2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G68), .ZN(new_n381));
  XNOR2_X1  g0181(.A(G58), .B(G68), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT16), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n386), .A3(new_n383), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n274), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n362), .B(new_n376), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n366), .A2(new_n367), .A3(G179), .ZN(new_n393));
  AOI21_X1  g0193(.A(G169), .B1(new_n369), .B2(new_n374), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n389), .B1(new_n385), .B2(new_n387), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n361), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT18), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n395), .B(new_n399), .C1(new_n396), .C2(new_n361), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n396), .A2(new_n361), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n376), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n392), .A2(new_n398), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n224), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n257), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n328), .A2(new_n259), .ZN(new_n407));
  INV_X1    g0207(.A(G107), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n255), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n250), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n267), .B1(new_n269), .B2(G244), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n292), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n354), .A3(new_n411), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT69), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n276), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n279), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT15), .B(G87), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n280), .B1(new_n211), .B2(new_n261), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n274), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n285), .A2(G77), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(G77), .B2(new_n287), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n412), .A2(G169), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n410), .A2(G179), .A3(new_n411), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n404), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n306), .A2(new_n358), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G250), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n253), .B2(new_n254), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n259), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n255), .A2(G257), .A3(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G294), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n250), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT5), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT75), .B1(new_n441), .B2(G41), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n336), .A3(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(G41), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n337), .A2(G1), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n442), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n332), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G264), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n264), .A2(G45), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n441), .B2(G41), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(G274), .A3(new_n444), .A4(new_n442), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n440), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G169), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n440), .A2(new_n450), .A3(G179), .A4(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n284), .A2(G20), .A3(new_n408), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT25), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n264), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n389), .A2(new_n285), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(G107), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n255), .A2(new_n211), .A3(G87), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT22), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n255), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT23), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n408), .A3(G20), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(KEYINPUT80), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT24), .B1(new_n468), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(KEYINPUT24), .A3(new_n466), .A4(new_n467), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n274), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n463), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n457), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n454), .A2(new_n292), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n454), .A2(G190), .ZN(new_n486));
  OAI221_X1 g0286(.A(new_n463), .B1(new_n478), .B2(new_n480), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n457), .A2(new_n481), .A3(KEYINPUT81), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g0290(.A(G1698), .B1(new_n435), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n490), .A2(G1698), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n255), .A2(G244), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G244), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n490), .B1(new_n327), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n491), .A2(new_n492), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n250), .ZN(new_n498));
  INV_X1    g0298(.A(G257), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n453), .B1(new_n448), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n354), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n497), .B2(new_n250), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G200), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n359), .A2(G97), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n461), .B2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT73), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT7), .B1(new_n327), .B2(new_n211), .ZN(new_n509));
  NOR4_X1   g0309(.A1(new_n325), .A2(new_n326), .A3(new_n377), .A4(G20), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n508), .B(G107), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n276), .A2(G77), .ZN(new_n512));
  OR2_X1    g0312(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n408), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  XOR2_X1   g0316(.A(KEYINPUT72), .B(KEYINPUT6), .Z(new_n517));
  XNOR2_X1  g0317(.A(G97), .B(G107), .ZN(new_n518));
  OAI211_X1 g0318(.A(G20), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n511), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n508), .B1(new_n380), .B2(G107), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT74), .B(new_n274), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n509), .B2(new_n510), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT73), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n519), .A2(new_n512), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n511), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT74), .B1(new_n527), .B2(new_n274), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n504), .B(new_n507), .C1(new_n523), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n255), .A2(new_n211), .A3(G68), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n211), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n371), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(G107), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n532), .B1(new_n531), .B2(G20), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n530), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n274), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n359), .A2(new_n420), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n539), .B(new_n540), .C1(new_n420), .C2(new_n461), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT76), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n266), .B1(new_n542), .B2(new_n434), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n446), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n451), .A2(new_n542), .A3(G250), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n250), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n255), .A2(G238), .A3(new_n259), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n255), .A2(G244), .A3(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n546), .B1(new_n550), .B2(new_n250), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G179), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n322), .B2(new_n551), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n250), .ZN(new_n554));
  INV_X1    g0354(.A(new_n546), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n354), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G200), .B2(new_n551), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n462), .A2(G87), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n539), .A2(new_n558), .A3(new_n540), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n541), .A2(new_n553), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n527), .A2(new_n274), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT74), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n506), .B1(new_n563), .B2(new_n522), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n498), .A2(new_n501), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G169), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n503), .A2(G179), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n529), .B(new_n560), .C1(new_n564), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n447), .A2(new_n332), .A3(G270), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n571), .A2(new_n453), .ZN(new_n572));
  OAI211_X1 g0372(.A(G264), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(new_n259), .C1(new_n325), .C2(new_n326), .ZN(new_n574));
  INV_X1    g0374(.A(G303), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(new_n255), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n250), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G20), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n274), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n492), .B(new_n211), .C1(G33), .C2(new_n534), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(KEYINPUT77), .A3(KEYINPUT20), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n274), .A3(new_n580), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n274), .A4(new_n580), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n583), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n285), .A2(G116), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n462), .B2(G116), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n578), .A2(G179), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n322), .B1(new_n572), .B2(new_n577), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(KEYINPUT21), .A3(new_n593), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n595), .A2(KEYINPUT78), .A3(new_n593), .A4(KEYINPUT21), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n578), .A2(new_n354), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(G200), .B2(new_n578), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n590), .A3(new_n592), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT79), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n595), .A2(new_n605), .A3(new_n593), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n595), .B2(new_n593), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n600), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n489), .A2(new_n570), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n433), .A2(new_n610), .ZN(G372));
  NAND2_X1  g0411(.A1(new_n553), .A2(new_n541), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n487), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n570), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n457), .A2(new_n481), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n457), .B2(new_n481), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n600), .B(new_n608), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n613), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n507), .B1(new_n523), .B2(new_n528), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n560), .A3(new_n568), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(KEYINPUT83), .A3(new_n623), .ZN(new_n627));
  XOR2_X1   g0427(.A(KEYINPUT84), .B(KEYINPUT26), .Z(new_n628));
  NAND4_X1  g0428(.A1(new_n621), .A2(new_n560), .A3(new_n568), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n433), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n305), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n398), .A2(new_n400), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n351), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n357), .B2(new_n430), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n392), .A2(new_n402), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n633), .B1(new_n639), .B2(new_n301), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT85), .ZN(G369));
  NAND2_X1  g0442(.A1(new_n600), .A2(new_n608), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n264), .A2(G13), .ZN(new_n644));
  OR3_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .A3(G20), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT27), .B1(new_n644), .B2(G20), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G343), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT86), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n593), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n609), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G330), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n484), .A2(new_n488), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n481), .A2(new_n649), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT87), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n657), .A3(new_n487), .ZN(new_n658));
  INV_X1    g0458(.A(new_n649), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n482), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n617), .A2(new_n618), .A3(new_n649), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n643), .A2(new_n659), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n658), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(G399));
  NOR2_X1   g0467(.A1(new_n220), .A2(G41), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n535), .A2(G107), .A3(G116), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n668), .A2(new_n264), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n209), .B2(new_n668), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT28), .Z(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n565), .A2(new_n454), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n578), .A2(G179), .A3(new_n551), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n551), .A2(new_n450), .A3(new_n440), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(G179), .A3(new_n578), .A4(new_n503), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n678), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n649), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT31), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(KEYINPUT88), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT31), .B(new_n649), .C1(new_n681), .C2(new_n682), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT88), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n683), .B2(new_n684), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n610), .A2(new_n659), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n674), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n621), .A2(new_n568), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n487), .A3(new_n560), .A4(new_n529), .ZN(new_n696));
  INV_X1    g0496(.A(new_n643), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n655), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n613), .B1(new_n622), .B2(new_n628), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(KEYINPUT26), .B2(new_n622), .ZN(new_n700));
  OAI211_X1 g0500(.A(KEYINPUT29), .B(new_n659), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n649), .B1(new_n620), .B2(new_n630), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(KEYINPUT29), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n673), .B1(new_n704), .B2(G1), .ZN(G364));
  NOR2_X1   g0505(.A1(new_n303), .A2(new_n292), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n211), .A2(G190), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(KEYINPUT33), .A2(G317), .ZN(new_n710));
  AND2_X1   g0510(.A1(KEYINPUT33), .A2(G317), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G283), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n292), .A2(G179), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n211), .A2(new_n354), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n714), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(G303), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT91), .B1(G179), .B2(G200), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(KEYINPUT91), .A2(G179), .A3(G200), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n211), .B1(new_n725), .B2(G190), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G294), .ZN(new_n728));
  INV_X1    g0528(.A(new_n707), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G329), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n717), .A2(new_n706), .ZN(new_n732));
  INV_X1    g0532(.A(G326), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n303), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n707), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G311), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n327), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n717), .A2(new_n735), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n734), .B(new_n738), .C1(G322), .C2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n720), .A2(new_n728), .A3(new_n731), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n726), .A2(new_n534), .ZN(new_n743));
  INV_X1    g0543(.A(new_n732), .ZN(new_n744));
  INV_X1    g0544(.A(new_n715), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n744), .A2(G50), .B1(new_n745), .B2(G107), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n202), .B2(new_n739), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n255), .B1(new_n708), .B2(new_n203), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n718), .A2(new_n371), .B1(new_n736), .B2(new_n261), .ZN(new_n749));
  OR4_X1    g0549(.A1(new_n743), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n730), .A2(G159), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT32), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n742), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n210), .B1(G20), .B2(new_n322), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n217), .A2(G20), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n668), .A2(new_n264), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n220), .A2(new_n327), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n761), .A2(G355), .B1(new_n579), .B2(new_n220), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n209), .A2(G45), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n245), .B2(G45), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n220), .A2(new_n255), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n762), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n754), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT90), .Z(new_n772));
  AOI21_X1  g0572(.A(new_n760), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n755), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT92), .Z(new_n775));
  NAND2_X1  g0575(.A1(new_n651), .A2(new_n652), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n770), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n777), .A2(G330), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT89), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n759), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(new_n781), .B2(new_n653), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n779), .B1(new_n783), .B2(new_n784), .ZN(G396));
  INV_X1    g0585(.A(new_n754), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n769), .ZN(new_n787));
  INV_X1    g0587(.A(G150), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n708), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G137), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n732), .A2(new_n790), .B1(new_n736), .B2(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n789), .B(new_n792), .C1(G143), .C2(new_n740), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G58), .B2(new_n727), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n327), .B1(new_n719), .B2(G50), .ZN(new_n796));
  INV_X1    g0596(.A(new_n730), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n203), .B2(new_n715), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(KEYINPUT34), .B2(new_n793), .ZN(new_n800));
  INV_X1    g0600(.A(new_n743), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n255), .B1(new_n740), .B2(G294), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n745), .A2(G87), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n575), .C2(new_n732), .ZN(new_n804));
  INV_X1    g0604(.A(new_n736), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G107), .A2(new_n719), .B1(new_n805), .B2(G116), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n713), .B2(new_n708), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(G311), .C2(new_n730), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n795), .A2(new_n800), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n759), .B1(G77), .B2(new_n787), .C1(new_n809), .C2(new_n786), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n426), .B(new_n649), .C1(new_n428), .C2(new_n429), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n649), .A2(new_n425), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n427), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(new_n813), .B2(new_n431), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n810), .B1(new_n815), .B2(new_n768), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n702), .B(new_n815), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(new_n693), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n759), .B1(new_n817), .B2(new_n693), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G384));
  NOR2_X1   g0621(.A1(new_n517), .A2(new_n518), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n517), .B2(new_n514), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT35), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(KEYINPUT35), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n824), .A2(G116), .A3(new_n212), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n827));
  XNOR2_X1  g0627(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n209), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n201), .A2(G68), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n264), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n433), .B(new_n701), .C1(KEYINPUT29), .C2(new_n702), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n640), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT99), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n635), .A2(new_n647), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n351), .B(new_n357), .C1(new_n320), .C2(new_n659), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT94), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n351), .B2(new_n659), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n352), .A2(G169), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT14), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(new_n347), .A3(new_n349), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n842), .A2(KEYINPUT94), .A3(new_n321), .A4(new_n649), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n837), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n627), .A2(new_n629), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT83), .B1(new_n622), .B2(new_n623), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n619), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n612), .B1(new_n848), .B2(new_n696), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n659), .B(new_n814), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n811), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT95), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n384), .A2(new_n853), .A3(new_n386), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n381), .B(new_n383), .C1(KEYINPUT95), .C2(KEYINPUT16), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n274), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n362), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n647), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n403), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n647), .B1(new_n396), .B2(new_n361), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n390), .A2(new_n397), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n857), .A2(new_n395), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n864), .A2(new_n858), .A3(new_n390), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n865), .B2(new_n861), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n860), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n860), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n836), .B1(new_n852), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT96), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT39), .B1(new_n867), .B2(new_n868), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n860), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n392), .A2(KEYINPUT98), .A3(new_n402), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT98), .B1(new_n392), .B2(new_n402), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n635), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n862), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n390), .A2(new_n397), .A3(new_n862), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n877), .A2(new_n878), .B1(new_n863), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n874), .B1(new_n881), .B2(KEYINPUT38), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n873), .B1(new_n882), .B2(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n636), .A2(new_n659), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT97), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n871), .A2(new_n872), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n871), .A2(new_n872), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n835), .B(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n685), .A2(new_n687), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n610), .B2(new_n659), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n891), .A2(new_n844), .A3(new_n815), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n882), .A3(KEYINPUT40), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n692), .A2(new_n685), .A3(new_n687), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n837), .A2(new_n839), .A3(new_n843), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n814), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n894), .B1(new_n897), .B2(new_n869), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n433), .A2(new_n895), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(G330), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n264), .B2(new_n756), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n889), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n832), .B1(new_n904), .B2(new_n905), .ZN(G367));
  OAI22_X1  g0706(.A1(new_n718), .A2(new_n202), .B1(new_n736), .B2(new_n201), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(G159), .B2(new_n709), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n327), .B1(new_n744), .B2(G143), .ZN(new_n909));
  AOI22_X1  g0709(.A1(G150), .A2(new_n740), .B1(new_n745), .B2(G77), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n911), .B1(new_n203), .B2(new_n726), .C1(new_n790), .C2(new_n797), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n726), .A2(new_n408), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n718), .A2(KEYINPUT46), .A3(new_n579), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT46), .B1(new_n718), .B2(new_n579), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(new_n730), .B2(G317), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n255), .B1(new_n805), .B2(G283), .ZN(new_n917));
  AOI22_X1  g0717(.A1(G311), .A2(new_n744), .B1(new_n740), .B2(G303), .ZN(new_n918));
  AOI22_X1  g0718(.A1(G294), .A2(new_n709), .B1(new_n745), .B2(G97), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n912), .B1(new_n913), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n786), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n771), .B1(new_n219), .B2(new_n420), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n241), .B2(new_n765), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n760), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n659), .A2(new_n559), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n560), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n612), .B2(new_n928), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n924), .B(new_n927), .C1(new_n930), .C2(new_n778), .ZN(new_n931));
  INV_X1    g0731(.A(new_n930), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n695), .B(new_n529), .C1(new_n564), .C2(new_n659), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n621), .A2(new_n568), .A3(new_n649), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(KEYINPUT100), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(KEYINPUT100), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT101), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n937), .B(KEYINPUT100), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(KEYINPUT101), .A3(new_n936), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n658), .A2(new_n664), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT42), .ZN(new_n948));
  INV_X1    g0748(.A(new_n655), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n649), .B1(new_n950), .B2(new_n695), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n934), .B(new_n935), .C1(new_n948), .C2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT42), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n947), .B(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n951), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(new_n933), .A4(new_n932), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n945), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n661), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n957), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n758), .A2(new_n264), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n658), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n482), .A2(new_n659), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n653), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n661), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n946), .B1(new_n968), .B2(new_n664), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n969), .A2(new_n703), .A3(new_n694), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n945), .A2(new_n666), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n945), .A2(KEYINPUT45), .A3(new_n666), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n942), .A2(new_n665), .A3(new_n944), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n977), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n942), .A2(new_n944), .A3(new_n665), .A4(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n975), .A2(new_n981), .A3(new_n661), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n970), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n661), .B1(new_n975), .B2(new_n981), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n704), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n668), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n963), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n931), .B1(new_n961), .B2(new_n988), .ZN(G387));
  AOI21_X1  g0789(.A(new_n766), .B1(new_n238), .B2(G45), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n670), .B2(new_n761), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n278), .A2(new_n201), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT50), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n337), .B1(new_n203), .B2(new_n261), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n993), .A2(new_n670), .A3(new_n994), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n991), .A2(new_n995), .B1(G107), .B2(new_n219), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n996), .A2(new_n772), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n718), .A2(new_n261), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n255), .B1(new_n715), .B2(new_n534), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G150), .C2(new_n730), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT104), .Z(new_n1001));
  OR2_X1    g0801(.A1(new_n726), .A2(new_n420), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G50), .A2(new_n740), .B1(new_n709), .B2(new_n278), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n744), .A2(G159), .B1(new_n805), .B2(G68), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n719), .A2(G294), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n744), .A2(G322), .B1(new_n805), .B2(G303), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(new_n737), .B2(new_n708), .C1(new_n1008), .C2(new_n739), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT48), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1006), .B1(new_n713), .B2(new_n726), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT105), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n327), .B1(new_n579), .B2(new_n715), .C1(new_n797), .C2(new_n733), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1005), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n760), .B(new_n997), .C1(new_n1018), .C2(new_n754), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n966), .A2(new_n770), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1019), .A2(new_n1020), .B1(new_n969), .B2(new_n963), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n970), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n668), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n704), .A2(new_n969), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G393));
  OAI21_X1  g0825(.A(new_n982), .B1(new_n984), .B2(KEYINPUT107), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n972), .B(new_n665), .C1(new_n942), .C2(new_n944), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT45), .B1(new_n945), .B2(new_n666), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n980), .B(new_n978), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n661), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT107), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT108), .B1(new_n1026), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n984), .A2(KEYINPUT107), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT108), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n982), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n963), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G303), .A2(new_n709), .B1(new_n805), .B2(G294), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n726), .B2(new_n579), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT111), .Z(new_n1043));
  OAI22_X1  g0843(.A1(new_n732), .A2(new_n1008), .B1(new_n739), .B2(new_n737), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n327), .B1(new_n715), .B2(new_n408), .C1(new_n713), .C2(new_n718), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G322), .B2(new_n730), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT112), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G68), .A2(new_n719), .B1(new_n805), .B2(new_n278), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n201), .B2(new_n708), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n727), .A2(G77), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1052), .A2(new_n1053), .A3(new_n255), .A4(new_n803), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT51), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n732), .A2(new_n788), .B1(new_n739), .B2(new_n791), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1055), .A2(new_n1056), .B1(new_n730), .B2(G143), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT110), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1048), .A2(KEYINPUT112), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1049), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n754), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n771), .B1(new_n534), .B2(new_n219), .C1(new_n766), .C2(new_n248), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1064), .A2(KEYINPUT109), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(KEYINPUT109), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1065), .A2(new_n1066), .A3(new_n760), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1063), .B(new_n1067), .C1(new_n945), .C2(new_n778), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n668), .B1(new_n983), .B2(new_n984), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1022), .B1(new_n1026), .B2(new_n1033), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1040), .A2(new_n1073), .ZN(G390));
  INV_X1    g0874(.A(new_n883), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT113), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n850), .A2(new_n851), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n896), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n885), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n852), .A2(KEYINPUT113), .A3(new_n885), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n813), .A2(new_n431), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n659), .B(new_n1083), .C1(new_n698), .C2(new_n700), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n851), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n882), .B(new_n1079), .C1(new_n1085), .C2(new_n844), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n693), .A2(new_n814), .A3(new_n896), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1082), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n814), .A2(G330), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n891), .A2(new_n844), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT113), .B1(new_n852), .B2(new_n885), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n811), .B1(new_n702), .B2(new_n814), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1076), .B(new_n1079), .C1(new_n1092), .C2(new_n844), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n883), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1086), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n433), .A2(G330), .A3(new_n895), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n833), .A2(new_n640), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n896), .B1(new_n693), .B2(new_n814), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1077), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n844), .B1(new_n891), .B2(new_n1089), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1087), .A2(new_n1085), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1098), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1088), .A2(new_n1096), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT114), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1088), .A2(new_n1096), .A3(new_n1106), .A4(new_n1103), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n668), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1088), .A2(new_n1096), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1103), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1110), .A2(new_n962), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n759), .B1(new_n278), .B2(new_n787), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n708), .A2(new_n408), .B1(new_n715), .B2(new_n203), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n255), .B(new_n1116), .C1(G87), .C2(new_n719), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n730), .A2(G294), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n732), .A2(new_n713), .B1(new_n739), .B2(new_n579), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G97), .B2(new_n805), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n1053), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n718), .A2(new_n788), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n805), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1123), .B(new_n1126), .C1(new_n1127), .C2(new_n797), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n732), .A2(new_n1129), .B1(new_n715), .B2(new_n201), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G137), .B2(new_n709), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n327), .B1(new_n740), .B2(G132), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n791), .C2(new_n726), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1121), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1115), .B1(new_n1134), .B2(new_n754), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n883), .B2(new_n769), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT116), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1114), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1113), .A2(new_n1138), .ZN(G378));
  OAI21_X1  g0939(.A(new_n759), .B1(G50), .B2(new_n787), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G116), .A2(new_n744), .B1(new_n740), .B2(G107), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n534), .B2(new_n708), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n327), .A2(new_n336), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n202), .A2(new_n715), .B1(new_n736), .B2(new_n420), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1142), .A2(new_n998), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n203), .B2(new_n726), .C1(new_n713), .C2(new_n797), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT58), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G50), .B1(new_n252), .B2(new_n336), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1146), .A2(new_n1147), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n708), .A2(new_n798), .B1(new_n736), .B2(new_n790), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n732), .A2(new_n1127), .B1(new_n739), .B2(new_n1129), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n719), .C2(new_n1125), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n788), .B2(new_n726), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n252), .B(new_n336), .C1(new_n715), .C2(new_n791), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G124), .B2(new_n730), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1149), .B1(new_n1147), .B2(new_n1146), .C1(new_n1155), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1140), .B1(new_n1160), .B2(new_n754), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n306), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n301), .A2(new_n305), .A3(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n289), .A2(new_n647), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT55), .Z(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1164), .A2(new_n1168), .A3(new_n1165), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1161), .B1(new_n1172), .B2(new_n769), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT119), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n893), .A2(new_n898), .A3(G330), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1172), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(new_n898), .A3(G330), .A4(new_n893), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1177), .A2(new_n886), .A3(new_n1179), .A4(new_n887), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1177), .A2(new_n1179), .B1(new_n886), .B2(new_n887), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT120), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n888), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT120), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(new_n1180), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1175), .B1(new_n1188), .B2(new_n962), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1098), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1108), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT57), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1109), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1098), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n1188), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1189), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n963), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n844), .A2(new_n768), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT121), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n759), .B1(G68), .B2(new_n787), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT122), .Z(new_n1206));
  AOI22_X1  g1006(.A1(new_n744), .A2(G294), .B1(new_n805), .B2(G107), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n534), .B2(new_n718), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n255), .B1(new_n745), .B2(G77), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n579), .B2(new_n708), .C1(new_n713), .C2(new_n739), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G303), .C2(new_n730), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n739), .A2(new_n790), .B1(new_n736), .B2(new_n788), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G132), .B2(new_n744), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1125), .A2(new_n709), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n327), .B1(new_n745), .B2(G58), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G50), .B2(new_n727), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n730), .A2(G128), .B1(G159), .B2(new_n719), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT123), .Z(new_n1219));
  AOI22_X1  g1019(.A1(new_n1211), .A2(new_n1002), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1204), .B(new_n1206), .C1(new_n786), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1202), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1201), .A2(new_n1190), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1111), .A2(new_n987), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1199), .A2(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G384), .A2(G381), .A3(G387), .A4(new_n1230), .ZN(new_n1231));
  OR3_X1    g1031(.A1(new_n1229), .A2(new_n1231), .A3(G390), .ZN(G407));
  INV_X1    g1032(.A(G343), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G213), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT125), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(new_n1229), .C2(new_n1236), .ZN(G409));
  NAND3_X1  g1037(.A1(G387), .A2(new_n1040), .A3(new_n1073), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n931), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n985), .A2(new_n987), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n962), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n957), .B(new_n959), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1239), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(G390), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1238), .A2(new_n1244), .ZN(new_n1245));
  XOR2_X1   g1045(.A(G393), .B(G396), .Z(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1243), .B2(G390), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n970), .B1(new_n1250), .B2(new_n1036), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1068), .B1(new_n1251), .B2(new_n1070), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n962), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT126), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1040), .A2(new_n1073), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1243), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1248), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(KEYINPUT127), .B(new_n1243), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1247), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1225), .A2(new_n1263), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1201), .A2(new_n1190), .A3(KEYINPUT60), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n668), .B(new_n1111), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1224), .A2(G384), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G384), .B1(new_n1224), .B2(new_n1266), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G2897), .B(new_n1235), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1268), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1224), .A2(G384), .A3(new_n1266), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1235), .A2(G2897), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1187), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1186), .B1(new_n1185), .B2(new_n1180), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1191), .A2(new_n987), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1174), .B1(new_n1192), .B2(new_n963), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G378), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1199), .B2(G378), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1274), .B1(new_n1281), .B2(new_n1235), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1174), .B1(new_n1277), .B2(new_n963), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1277), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n668), .B1(new_n1197), .B2(new_n1193), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1284), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1197), .A2(new_n1188), .A3(new_n986), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1279), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1228), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1236), .A4(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1282), .A2(new_n1283), .A3(new_n1295), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1235), .B(new_n1293), .C1(new_n1287), .C2(new_n1290), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(new_n1292), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1262), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1261), .A2(new_n1283), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(KEYINPUT63), .B2(new_n1297), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1235), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1294), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1301), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1299), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(new_n1262), .A2(new_n1294), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1199), .B(G378), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1261), .A2(new_n1293), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(G402));
endmodule


