//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n461), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n461), .A2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n461), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n478), .B1(G136), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n462), .B2(new_n463), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n463), .C2(new_n462), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(G50), .A3(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT70), .B1(new_n504), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT5), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n505), .A2(new_n508), .B1(new_n504), .B2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n499), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  OAI221_X1 g086(.A(new_n502), .B1(new_n503), .B2(new_n510), .C1(new_n496), .C2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  XOR2_X1   g088(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n516), .B(KEYINPUT73), .C1(new_n517), .C2(new_n510), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  INV_X1    g097(.A(new_n498), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n497), .A2(KEYINPUT71), .A3(new_n498), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G543), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(G51), .B1(new_n509), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n520), .A2(new_n521), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n496), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n510), .A2(new_n535), .B1(new_n527), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G171));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n510), .A2(new_n542), .B1(new_n527), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI221_X1 g121(.A(KEYINPUT76), .B1(new_n527), .B2(new_n543), .C1(new_n510), .C2(new_n542), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n505), .A2(new_n508), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n504), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n496), .B1(new_n553), .B2(KEYINPUT75), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n546), .A2(new_n547), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT78), .Z(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n527), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n507), .B1(new_n499), .B2(new_n522), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .A3(G53), .A4(new_n526), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  AND2_X1   g145(.A1(KEYINPUT79), .A2(G65), .ZN(new_n571));
  NOR2_X1   g146(.A1(KEYINPUT79), .A2(G65), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n570), .B1(new_n551), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n499), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n551), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n575), .A2(G651), .B1(new_n577), .B2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n569), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  NAND2_X1  g155(.A1(new_n531), .A2(KEYINPUT80), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n520), .A2(new_n582), .A3(new_n521), .A4(new_n530), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G286));
  NAND2_X1  g160(.A1(new_n577), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n528), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G288));
  AOI22_X1  g168(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n496), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n509), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n576), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n496), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n510), .A2(new_n602), .B1(new_n527), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n601), .A2(new_n604), .ZN(G290));
  NAND3_X1  g180(.A1(new_n577), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n510), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n551), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(G651), .B1(new_n528), .B2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g192(.A(new_n616), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n566), .A2(new_n568), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n509), .A2(G91), .A3(new_n499), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n509), .A2(new_n573), .B1(G78), .B2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n496), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n619), .B1(new_n624), .B2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  MUX2_X1   g201(.A(new_n619), .B(new_n625), .S(new_n626), .Z(G297));
  MUX2_X1   g202(.A(new_n619), .B(new_n625), .S(new_n626), .Z(G280));
  AND2_X1   g203(.A1(new_n610), .A2(new_n614), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n634), .B(new_n635), .C1(G868), .C2(new_n556), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n472), .A2(new_n468), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n480), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n474), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n461), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n643), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT85), .Z(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT86), .Z(G401));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT17), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n669), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n671), .A3(new_n669), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n671), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n670), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n688), .A2(new_n689), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(new_n692), .A3(new_n690), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n697), .C1(new_n692), .C2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G33), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT25), .Z(new_n708));
  INV_X1    g283(.A(G139), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n479), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n714));
  OAI22_X1  g289(.A1(new_n712), .A2(new_n713), .B1(new_n461), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT96), .Z(new_n716));
  OAI21_X1  g291(.A(new_n706), .B1(new_n716), .B2(new_n705), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G2072), .Z(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G5), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G171), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  NOR2_X1   g297(.A1(G29), .A2(G35), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G162), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT29), .Z(new_n725));
  OAI221_X1 g300(.A(new_n718), .B1(G1961), .B2(new_n721), .C1(new_n722), .C2(new_n725), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(new_n722), .B1(G1961), .B2(new_n721), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT31), .B(G11), .Z(new_n728));
  NOR2_X1   g303(.A1(new_n648), .A2(new_n705), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT97), .B(G28), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n730), .B2(KEYINPUT30), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n728), .B(new_n729), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G27), .A2(G29), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G164), .B2(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G2078), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n705), .B1(new_n737), .B2(G34), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n737), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G160), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n733), .A2(new_n736), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n705), .A2(G32), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  INV_X1    g321(.A(G129), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n473), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n468), .A2(G105), .ZN(new_n749));
  INV_X1    g324(.A(G141), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n479), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n744), .B1(new_n753), .B2(new_n705), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G2078), .B2(new_n735), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n629), .A2(G16), .ZN(new_n759));
  OR2_X1    g334(.A1(G4), .A2(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n743), .B(new_n757), .C1(new_n758), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n705), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  OR2_X1    g339(.A1(G104), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT93), .Z(new_n767));
  INV_X1    g342(.A(G128), .ZN(new_n768));
  INV_X1    g343(.A(G140), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n768), .A2(new_n473), .B1(new_n479), .B2(new_n769), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n767), .A2(KEYINPUT94), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT94), .B1(new_n767), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n764), .B1(new_n773), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n761), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(G1348), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n719), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n719), .ZN(new_n780));
  INV_X1    g355(.A(G1966), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n727), .A2(new_n762), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n556), .B2(G16), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n719), .A2(G20), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT23), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G299), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n726), .A2(new_n783), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n719), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n719), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1971), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n719), .A2(G6), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n598), .B2(new_n719), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT90), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n719), .A2(G23), .ZN(new_n802));
  INV_X1    g377(.A(new_n589), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n719), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT33), .B(G1976), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT91), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n795), .A2(new_n800), .A3(new_n801), .A4(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(G16), .Z(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(G1986), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n480), .A2(G131), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n474), .A2(G119), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n461), .A2(G107), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G25), .B(new_n817), .S(G29), .Z(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n812), .A2(KEYINPUT92), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G1986), .B2(new_n811), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n809), .A2(new_n810), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n792), .A2(new_n825), .A3(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  AOI22_X1  g404(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n496), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT98), .B(G93), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n510), .A2(new_n832), .B1(new_n527), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n629), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  INV_X1    g416(.A(new_n835), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n556), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n836), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n838), .B1(new_n846), .B2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n773), .B(G164), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n716), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n753), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n753), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n480), .A2(G142), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT100), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n474), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n461), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n817), .B(new_n639), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n851), .A2(new_n852), .A3(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n648), .B(G160), .Z(new_n862));
  XNOR2_X1  g437(.A(G162), .B(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n851), .A2(new_n852), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n860), .B(KEYINPUT101), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n861), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n863), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n851), .A2(new_n852), .A3(new_n865), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n851), .B2(new_n852), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(new_n843), .B(new_n632), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n629), .A2(new_n624), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n615), .A2(G299), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(KEYINPUT41), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n881), .A3(new_n876), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(KEYINPUT102), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n878), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n879), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n589), .B(KEYINPUT103), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G303), .ZN(new_n891));
  XNOR2_X1  g466(.A(G290), .B(new_n598), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n891), .B(new_n892), .Z(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n888), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n889), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n889), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(G868), .B2(new_n835), .ZN(G295));
  OAI21_X1  g473(.A(new_n897), .B1(G868), .B2(new_n835), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n584), .A2(G171), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n556), .B(new_n835), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n539), .A2(new_n531), .A3(new_n540), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n581), .A2(new_n583), .B1(new_n539), .B2(new_n540), .ZN(new_n906));
  INV_X1    g481(.A(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n843), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n878), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n891), .B(new_n892), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n905), .A2(new_n908), .A3(new_n883), .A4(new_n885), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n880), .A2(new_n914), .A3(new_n882), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n878), .A2(KEYINPUT104), .A3(new_n881), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n905), .A2(new_n908), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n871), .B(new_n913), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  AND4_X1   g495(.A1(new_n905), .A2(new_n908), .A3(new_n915), .A4(new_n916), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n877), .B1(new_n905), .B2(new_n908), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n893), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(KEYINPUT105), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n901), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n913), .A2(new_n871), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n918), .A2(new_n919), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(KEYINPUT106), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n900), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n912), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n893), .B1(new_n931), .B2(new_n922), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT43), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n920), .A2(new_n924), .A3(KEYINPUT43), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n900), .B1(new_n926), .B2(new_n932), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(G164), .B2(G1384), .ZN(new_n941));
  INV_X1    g516(.A(G40), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n466), .A2(new_n470), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n491), .A2(new_n493), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n483), .A2(new_n486), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n941), .A2(new_n943), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n951), .A3(new_n947), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n943), .A3(new_n952), .ZN(new_n953));
  OAI22_X1  g528(.A1(new_n949), .A2(G1971), .B1(G2090), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G8), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n502), .B1(new_n503), .B2(new_n510), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n511), .A2(new_n496), .ZN(new_n957));
  OAI21_X1  g532(.A(G8), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n955), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(G8), .A3(new_n954), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n944), .B2(new_n945), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n943), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(G8), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n803), .A2(G1976), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n967), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1976), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n590), .A2(new_n974), .A3(new_n591), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n589), .A2(new_n974), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n976), .A2(new_n970), .A3(KEYINPUT52), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G1981), .B1(new_n595), .B2(new_n597), .ZN(new_n979));
  INV_X1    g554(.A(G1981), .ZN(new_n980));
  OAI221_X1 g555(.A(new_n980), .B1(new_n596), .B2(new_n576), .C1(new_n496), .C2(new_n594), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT49), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n970), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n981), .A3(KEYINPUT49), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n978), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n943), .B1(new_n968), .B2(new_n951), .ZN(new_n991));
  NOR3_X1   g566(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n941), .A2(new_n943), .A3(new_n948), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n993), .A2(new_n741), .B1(new_n994), .B2(new_n781), .ZN(new_n995));
  NOR3_X1   g570(.A1(G286), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n966), .A2(new_n989), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(KEYINPUT112), .A2(KEYINPUT63), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(KEYINPUT112), .A2(KEYINPUT63), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n966), .A2(new_n989), .A3(new_n996), .A4(new_n998), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n988), .A2(new_n974), .A3(new_n592), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n981), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n970), .B(KEYINPUT111), .Z(new_n1005));
  INV_X1    g580(.A(new_n965), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1004), .A2(new_n1005), .B1(new_n989), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1001), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1956), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n991), .B2(new_n992), .ZN(new_n1011));
  OR2_X1    g586(.A1(KEYINPUT113), .A2(KEYINPUT57), .ZN(new_n1012));
  NAND2_X1  g587(.A1(KEYINPUT113), .A2(KEYINPUT57), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n569), .A2(new_n578), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT113), .B(KEYINPUT57), .C1(new_n620), .C2(new_n623), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n941), .A2(new_n948), .A3(new_n943), .A4(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(KEYINPUT114), .A3(new_n1011), .A4(new_n1017), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1011), .A2(new_n1017), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n758), .B1(new_n991), .B2(new_n992), .ZN(new_n1025));
  INV_X1    g600(.A(new_n969), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n775), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n629), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1020), .A2(new_n1022), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(KEYINPUT60), .A3(new_n1027), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n615), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n615), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1028), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(KEYINPUT60), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1024), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT61), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1024), .A2(KEYINPUT61), .A3(new_n1018), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  INV_X1    g623(.A(new_n556), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT58), .B(G1341), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(new_n969), .B2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g628(.A(KEYINPUT115), .B(new_n1051), .C1(new_n968), .C2(new_n943), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1996), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n941), .A2(new_n948), .A3(new_n1056), .A4(new_n943), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1049), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT117), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT59), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n493), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n492), .B1(new_n472), .B2(new_n489), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n947), .B1(new_n1065), .B2(new_n487), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G160), .A2(G40), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1052), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT115), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n969), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1057), .A3(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1071), .A2(new_n1061), .A3(new_n556), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1060), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n556), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1059), .B1(new_n1074), .B2(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(KEYINPUT117), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1048), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1047), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1048), .A3(new_n1077), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1030), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n963), .A2(new_n978), .A3(new_n988), .A4(new_n965), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n990), .B1(new_n995), .B2(G168), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(G168), .B2(new_n995), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1082), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  INV_X1    g665(.A(G1961), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n953), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(G2078), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n994), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1090), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1092), .B(KEYINPUT120), .C1(new_n994), .C2(new_n1096), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n994), .B2(G2078), .ZN(new_n1102));
  AOI21_X1  g677(.A(G301), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1096), .B1(new_n1067), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n943), .A2(KEYINPUT122), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n941), .A3(new_n948), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1092), .A3(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(G171), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1089), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1100), .A2(G301), .A3(new_n1102), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1089), .B1(new_n1108), .B2(G171), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1088), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT123), .B(new_n1009), .C1(new_n1081), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n629), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1031), .A2(new_n1032), .A3(new_n615), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1038), .B1(new_n1120), .B2(new_n1033), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1023), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1046), .B1(new_n1122), .B2(KEYINPUT61), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1061), .B1(new_n1071), .B2(new_n556), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n1126));
  NOR4_X1   g701(.A1(new_n1072), .A2(new_n1125), .A3(new_n1126), .A4(new_n1059), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1071), .A2(new_n1059), .A3(new_n556), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1126), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1131), .A3(new_n1080), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1030), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1114), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1116), .B1(new_n1134), .B2(new_n1008), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT62), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n966), .A2(new_n1103), .A3(new_n989), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT124), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n1144));
  NOR4_X1   g719(.A1(new_n1137), .A2(new_n1140), .A3(new_n1144), .A4(new_n1141), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1115), .A2(new_n1135), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n773), .B(new_n775), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1056), .B2(new_n753), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n941), .A2(new_n1067), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1056), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT108), .Z(new_n1152));
  AOI22_X1  g727(.A1(new_n1149), .A2(new_n1150), .B1(new_n753), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n819), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n817), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n817), .A2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1150), .ZN(new_n1159));
  AND2_X1   g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT107), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT107), .B1(G290), .B2(G1986), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT109), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1147), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1152), .A2(KEYINPUT46), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1159), .B1(new_n1148), .B2(new_n753), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(KEYINPUT46), .B2(new_n1152), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT47), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(G2067), .B2(new_n773), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1150), .ZN(new_n1178));
  NOR2_X1   g753(.A1(G290), .A2(G1986), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1150), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT126), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT48), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1158), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT127), .B1(new_n1175), .B2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1186), .A2(new_n1187), .A3(new_n1183), .A4(new_n1178), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1167), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g765(.A1(G229), .A2(new_n459), .A3(new_n667), .A4(G227), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n872), .B(new_n1192), .C1(new_n937), .C2(new_n936), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


