

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731;

  INV_X1 U364 ( .A(G953), .ZN(n716) );
  XOR2_X1 U365 ( .A(n497), .B(n548), .Z(n343) );
  NOR2_X2 U366 ( .A1(n531), .A2(n656), .ZN(n661) );
  INV_X2 U367 ( .A(n545), .ZN(n653) );
  XNOR2_X2 U368 ( .A(n521), .B(KEYINPUT33), .ZN(n672) );
  NOR2_X2 U369 ( .A1(n530), .A2(n563), .ZN(n521) );
  XNOR2_X2 U370 ( .A(n498), .B(KEYINPUT19), .ZN(n571) );
  NOR2_X2 U371 ( .A1(n653), .A2(n512), .ZN(n636) );
  XNOR2_X2 U372 ( .A(n713), .B(G101), .ZN(n350) );
  XNOR2_X2 U373 ( .A(n483), .B(n421), .ZN(n713) );
  AND2_X1 U374 ( .A1(n346), .A2(n371), .ZN(n370) );
  XNOR2_X1 U375 ( .A(G104), .B(G110), .ZN(n424) );
  XNOR2_X1 U376 ( .A(G113), .B(KEYINPUT3), .ZN(n357) );
  XNOR2_X1 U377 ( .A(n368), .B(n367), .ZN(n700) );
  NAND2_X1 U378 ( .A1(n370), .A2(n369), .ZN(n368) );
  AND2_X1 U379 ( .A1(n380), .A2(n378), .ZN(n377) );
  NOR2_X1 U380 ( .A1(n516), .A2(n502), .ZN(n503) );
  XNOR2_X1 U381 ( .A(n438), .B(n429), .ZN(n624) );
  XNOR2_X1 U382 ( .A(n350), .B(n710), .ZN(n438) );
  XNOR2_X1 U383 ( .A(n357), .B(G119), .ZN(n447) );
  XNOR2_X1 U384 ( .A(n424), .B(G107), .ZN(n445) );
  XNOR2_X1 U385 ( .A(KEYINPUT4), .B(G146), .ZN(n420) );
  INV_X1 U386 ( .A(n360), .ZN(n359) );
  INV_X1 U387 ( .A(KEYINPUT85), .ZN(n355) );
  XNOR2_X1 U388 ( .A(n431), .B(n430), .ZN(n505) );
  XNOR2_X1 U389 ( .A(n725), .B(n513), .ZN(n349) );
  XNOR2_X1 U390 ( .A(n388), .B(n387), .ZN(n478) );
  INV_X1 U391 ( .A(KEYINPUT8), .ZN(n387) );
  NAND2_X1 U392 ( .A1(n716), .A2(G234), .ZN(n388) );
  XNOR2_X1 U393 ( .A(G113), .B(G143), .ZN(n461) );
  XOR2_X1 U394 ( .A(G122), .B(G104), .Z(n462) );
  XNOR2_X1 U395 ( .A(n451), .B(n450), .ZN(n453) );
  INV_X1 U396 ( .A(KEYINPUT18), .ZN(n450) );
  NOR2_X1 U397 ( .A1(n457), .A2(n363), .ZN(n361) );
  NAND2_X1 U398 ( .A1(n457), .A2(n363), .ZN(n362) );
  OR2_X1 U399 ( .A1(n608), .A2(n365), .ZN(n364) );
  XNOR2_X1 U400 ( .A(n501), .B(n500), .ZN(n516) );
  XNOR2_X1 U401 ( .A(n438), .B(n437), .ZN(n599) );
  XNOR2_X1 U402 ( .A(G110), .B(G128), .ZN(n397) );
  XNOR2_X1 U403 ( .A(n400), .B(n399), .ZN(n401) );
  INV_X1 U404 ( .A(KEYINPUT96), .ZN(n399) );
  XNOR2_X1 U405 ( .A(n549), .B(KEYINPUT39), .ZN(n590) );
  NAND2_X1 U406 ( .A1(n459), .A2(n343), .ZN(n549) );
  XNOR2_X1 U407 ( .A(n351), .B(KEYINPUT83), .ZN(n579) );
  XNOR2_X1 U408 ( .A(n575), .B(n355), .ZN(n354) );
  AND2_X1 U409 ( .A1(n353), .A2(n578), .ZN(n352) );
  INV_X1 U410 ( .A(n598), .ZN(n363) );
  XOR2_X1 U411 ( .A(G116), .B(G122), .Z(n477) );
  XNOR2_X1 U412 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n523) );
  AND2_X1 U413 ( .A1(n372), .A2(n522), .ZN(n383) );
  NOR2_X1 U414 ( .A1(n518), .A2(n517), .ZN(n520) );
  NAND2_X1 U415 ( .A1(n344), .A2(n358), .ZN(n498) );
  NOR2_X1 U416 ( .A1(n359), .A2(n366), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n505), .B(KEYINPUT1), .ZN(n518) );
  INV_X1 U418 ( .A(KEYINPUT45), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n472), .B(n471), .ZN(n616) );
  XNOR2_X1 U420 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U421 ( .A(G125), .B(KEYINPUT17), .ZN(n452) );
  NOR2_X1 U422 ( .A1(n566), .A2(n656), .ZN(n556) );
  INV_X1 U423 ( .A(n382), .ZN(n375) );
  NAND2_X1 U424 ( .A1(n383), .A2(n381), .ZN(n376) );
  OR2_X1 U425 ( .A1(n384), .A2(n381), .ZN(n380) );
  NOR2_X1 U426 ( .A1(n443), .A2(n444), .ZN(n459) );
  OR2_X1 U427 ( .A1(n599), .A2(G902), .ZN(n439) );
  BUF_X1 U428 ( .A(n518), .Z(n651) );
  XNOR2_X1 U429 ( .A(n503), .B(n504), .ZN(n356) );
  XNOR2_X1 U430 ( .A(n402), .B(n401), .ZN(n407) );
  XNOR2_X1 U431 ( .A(KEYINPUT40), .B(n550), .ZN(n730) );
  NOR2_X2 U432 ( .A1(n529), .A2(n528), .ZN(n642) );
  INV_X1 U433 ( .A(n664), .ZN(n366) );
  AND2_X1 U434 ( .A1(n364), .A2(n362), .ZN(n344) );
  AND2_X1 U435 ( .A1(n547), .A2(n629), .ZN(n345) );
  AND2_X1 U436 ( .A1(n525), .A2(n345), .ZN(n346) );
  NAND2_X1 U437 ( .A1(n347), .A2(n526), .ZN(n369) );
  NAND2_X1 U438 ( .A1(n348), .A2(KEYINPUT66), .ZN(n347) );
  NAND2_X1 U439 ( .A1(n349), .A2(n524), .ZN(n348) );
  XNOR2_X1 U440 ( .A(n455), .B(n350), .ZN(n608) );
  NAND2_X1 U441 ( .A1(n354), .A2(n352), .ZN(n351) );
  XNOR2_X1 U442 ( .A(n577), .B(KEYINPUT84), .ZN(n353) );
  NAND2_X1 U443 ( .A1(n490), .A2(n522), .ZN(n575) );
  NOR2_X1 U444 ( .A1(n558), .A2(n557), .ZN(n572) );
  NAND2_X1 U445 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U446 ( .A1(n356), .A2(n507), .ZN(n508) );
  NAND2_X1 U447 ( .A1(n356), .A2(n510), .ZN(n511) );
  AND2_X1 U448 ( .A1(n356), .A2(n563), .ZN(n543) );
  NAND2_X1 U449 ( .A1(n344), .A2(n360), .ZN(n497) );
  NAND2_X1 U450 ( .A1(n608), .A2(n361), .ZN(n360) );
  INV_X1 U451 ( .A(n457), .ZN(n365) );
  NAND2_X1 U452 ( .A1(n515), .A2(n514), .ZN(n371) );
  NAND2_X1 U453 ( .A1(n382), .A2(n383), .ZN(n379) );
  NAND2_X1 U454 ( .A1(n539), .A2(KEYINPUT34), .ZN(n372) );
  NAND2_X1 U455 ( .A1(n672), .A2(KEYINPUT34), .ZN(n382) );
  NAND2_X2 U456 ( .A1(n377), .A2(n373), .ZN(n725) );
  NAND2_X1 U457 ( .A1(n384), .A2(n374), .ZN(n373) );
  NOR2_X1 U458 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U459 ( .A1(n379), .A2(n523), .ZN(n378) );
  INV_X1 U460 ( .A(n523), .ZN(n381) );
  NAND2_X1 U461 ( .A1(n386), .A2(n385), .ZN(n384) );
  NOR2_X1 U462 ( .A1(n539), .A2(KEYINPUT34), .ZN(n385) );
  INV_X1 U463 ( .A(n672), .ZN(n386) );
  AND2_X1 U464 ( .A1(n391), .A2(n579), .ZN(n580) );
  XNOR2_X1 U465 ( .A(n445), .B(n425), .ZN(n426) );
  XNOR2_X1 U466 ( .A(n509), .B(KEYINPUT67), .ZN(n727) );
  XNOR2_X2 U467 ( .A(n419), .B(n418), .ZN(n483) );
  XNOR2_X2 U468 ( .A(G143), .B(G128), .ZN(n419) );
  BUF_X1 U469 ( .A(n688), .Z(n692) );
  XNOR2_X2 U470 ( .A(KEYINPUT65), .B(KEYINPUT81), .ZN(n418) );
  XOR2_X1 U471 ( .A(n404), .B(n403), .Z(n389) );
  XOR2_X1 U472 ( .A(n469), .B(n468), .Z(n390) );
  AND2_X1 U473 ( .A1(n728), .A2(n574), .ZN(n391) );
  XOR2_X1 U474 ( .A(n562), .B(KEYINPUT46), .Z(n392) );
  XNOR2_X1 U475 ( .A(G140), .B(KEYINPUT80), .ZN(n425) );
  INV_X1 U476 ( .A(KEYINPUT76), .ZN(n519) );
  XNOR2_X1 U477 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U478 ( .A(KEYINPUT70), .B(KEYINPUT0), .ZN(n500) );
  XNOR2_X1 U479 ( .A(n449), .B(n448), .ZN(n703) );
  XNOR2_X1 U480 ( .A(n470), .B(n390), .ZN(n472) );
  NOR2_X1 U481 ( .A1(n497), .A2(n583), .ZN(n568) );
  BUF_X1 U482 ( .A(n505), .Z(n558) );
  XNOR2_X1 U483 ( .A(n405), .B(n389), .ZN(n406) );
  XNOR2_X1 U484 ( .A(n407), .B(n406), .ZN(n408) );
  AND2_X1 U485 ( .A1(n602), .A2(G953), .ZN(n696) );
  XOR2_X1 U486 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n395) );
  XNOR2_X1 U487 ( .A(G902), .B(KEYINPUT15), .ZN(n598) );
  NAND2_X1 U488 ( .A1(G234), .A2(n598), .ZN(n393) );
  XNOR2_X1 U489 ( .A(KEYINPUT20), .B(n393), .ZN(n411) );
  NAND2_X1 U490 ( .A1(n411), .A2(G217), .ZN(n394) );
  XNOR2_X1 U491 ( .A(n395), .B(n394), .ZN(n410) );
  XOR2_X1 U492 ( .A(G140), .B(G125), .Z(n396) );
  XNOR2_X1 U493 ( .A(KEYINPUT10), .B(n396), .ZN(n711) );
  XNOR2_X1 U494 ( .A(G146), .B(n711), .ZN(n471) );
  XOR2_X1 U495 ( .A(KEYINPUT97), .B(KEYINPUT86), .Z(n398) );
  XNOR2_X1 U496 ( .A(n398), .B(n397), .ZN(n402) );
  XNOR2_X1 U497 ( .A(G119), .B(G137), .ZN(n400) );
  NAND2_X1 U498 ( .A1(G221), .A2(n478), .ZN(n405) );
  XOR2_X1 U499 ( .A(KEYINPUT24), .B(KEYINPUT79), .Z(n404) );
  XNOR2_X1 U500 ( .A(KEYINPUT23), .B(KEYINPUT95), .ZN(n403) );
  XNOR2_X1 U501 ( .A(n471), .B(n408), .ZN(n693) );
  NOR2_X1 U502 ( .A1(G902), .A2(n693), .ZN(n409) );
  XNOR2_X1 U503 ( .A(n410), .B(n409), .ZN(n545) );
  XOR2_X1 U504 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n413) );
  NAND2_X1 U505 ( .A1(n411), .A2(G221), .ZN(n412) );
  XNOR2_X1 U506 ( .A(n413), .B(n412), .ZN(n654) );
  NAND2_X1 U507 ( .A1(n653), .A2(n654), .ZN(n517) );
  NAND2_X1 U508 ( .A1(G234), .A2(G237), .ZN(n414) );
  XNOR2_X1 U509 ( .A(n414), .B(KEYINPUT14), .ZN(n415) );
  NAND2_X1 U510 ( .A1(G952), .A2(n415), .ZN(n679) );
  NOR2_X1 U511 ( .A1(n679), .A2(G953), .ZN(n495) );
  NAND2_X1 U512 ( .A1(G902), .A2(n415), .ZN(n493) );
  OR2_X1 U513 ( .A1(n716), .A2(n493), .ZN(n416) );
  NOR2_X1 U514 ( .A1(n416), .A2(G900), .ZN(n417) );
  NOR2_X1 U515 ( .A1(n495), .A2(n417), .ZN(n554) );
  NOR2_X1 U516 ( .A1(n517), .A2(n554), .ZN(n432) );
  XNOR2_X1 U517 ( .A(n420), .B(KEYINPUT64), .ZN(n421) );
  XNOR2_X1 U518 ( .A(G137), .B(G134), .ZN(n423) );
  INV_X1 U519 ( .A(G131), .ZN(n422) );
  XNOR2_X1 U520 ( .A(n423), .B(n422), .ZN(n710) );
  XOR2_X1 U521 ( .A(KEYINPUT94), .B(n426), .Z(n428) );
  NAND2_X1 U522 ( .A1(G227), .A2(n716), .ZN(n427) );
  XNOR2_X1 U523 ( .A(n428), .B(n427), .ZN(n429) );
  INV_X1 U524 ( .A(G902), .ZN(n486) );
  NAND2_X1 U525 ( .A1(n624), .A2(n486), .ZN(n431) );
  INV_X1 U526 ( .A(G469), .ZN(n430) );
  INV_X1 U527 ( .A(n558), .ZN(n536) );
  NAND2_X1 U528 ( .A1(n432), .A2(n536), .ZN(n444) );
  NOR2_X1 U529 ( .A1(G953), .A2(G237), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n467), .A2(G210), .ZN(n433) );
  XNOR2_X1 U531 ( .A(n433), .B(G116), .ZN(n435) );
  XNOR2_X1 U532 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n434) );
  XNOR2_X1 U533 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U534 ( .A(n447), .B(n436), .ZN(n437) );
  XNOR2_X2 U535 ( .A(n439), .B(G472), .ZN(n535) );
  NOR2_X1 U536 ( .A1(G902), .A2(G237), .ZN(n440) );
  XNOR2_X1 U537 ( .A(KEYINPUT77), .B(n440), .ZN(n456) );
  NAND2_X1 U538 ( .A1(n456), .A2(G214), .ZN(n664) );
  NAND2_X1 U539 ( .A1(n535), .A2(n664), .ZN(n442) );
  XNOR2_X1 U540 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n441) );
  XNOR2_X1 U541 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n445), .B(n477), .ZN(n449) );
  XNOR2_X1 U543 ( .A(KEYINPUT16), .B(KEYINPUT75), .ZN(n446) );
  NAND2_X1 U544 ( .A1(G224), .A2(n716), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n703), .B(n454), .ZN(n455) );
  NAND2_X1 U546 ( .A1(n456), .A2(G210), .ZN(n457) );
  INV_X1 U547 ( .A(n497), .ZN(n458) );
  NAND2_X1 U548 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U549 ( .A(n460), .B(KEYINPUT111), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT13), .B(G475), .ZN(n474) );
  XNOR2_X1 U551 ( .A(n462), .B(n461), .ZN(n466) );
  XOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n464) );
  XNOR2_X1 U553 ( .A(KEYINPUT12), .B(KEYINPUT102), .ZN(n463) );
  XNOR2_X1 U554 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U555 ( .A(n466), .B(n465), .ZN(n470) );
  XOR2_X1 U556 ( .A(G131), .B(KEYINPUT101), .Z(n469) );
  NAND2_X1 U557 ( .A1(G214), .A2(n467), .ZN(n468) );
  NOR2_X1 U558 ( .A1(G902), .A2(n616), .ZN(n473) );
  XNOR2_X1 U559 ( .A(n474), .B(n473), .ZN(n527) );
  XOR2_X1 U560 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n476) );
  XNOR2_X1 U561 ( .A(G107), .B(KEYINPUT7), .ZN(n475) );
  XNOR2_X1 U562 ( .A(n476), .B(n475), .ZN(n482) );
  XOR2_X1 U563 ( .A(n477), .B(G134), .Z(n480) );
  NAND2_X1 U564 ( .A1(G217), .A2(n478), .ZN(n479) );
  XNOR2_X1 U565 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U566 ( .A(n482), .B(n481), .ZN(n485) );
  INV_X1 U567 ( .A(n483), .ZN(n484) );
  XNOR2_X1 U568 ( .A(n485), .B(n484), .ZN(n690) );
  NAND2_X1 U569 ( .A1(n690), .A2(n486), .ZN(n487) );
  XNOR2_X1 U570 ( .A(n487), .B(G478), .ZN(n529) );
  AND2_X1 U571 ( .A1(n527), .A2(n529), .ZN(n489) );
  INV_X1 U572 ( .A(KEYINPUT107), .ZN(n488) );
  XNOR2_X1 U573 ( .A(n489), .B(n488), .ZN(n522) );
  XNOR2_X1 U574 ( .A(n575), .B(G143), .ZN(G45) );
  XOR2_X1 U575 ( .A(KEYINPUT22), .B(KEYINPUT73), .Z(n491) );
  XNOR2_X1 U576 ( .A(KEYINPUT74), .B(n491), .ZN(n504) );
  XNOR2_X1 U577 ( .A(G898), .B(KEYINPUT91), .ZN(n699) );
  NAND2_X1 U578 ( .A1(n699), .A2(G953), .ZN(n492) );
  XNOR2_X1 U579 ( .A(n492), .B(KEYINPUT92), .ZN(n704) );
  NOR2_X1 U580 ( .A1(n704), .A2(n493), .ZN(n494) );
  NOR2_X1 U581 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U582 ( .A(KEYINPUT93), .B(n496), .ZN(n499) );
  NAND2_X1 U583 ( .A1(n499), .A2(n571), .ZN(n501) );
  NOR2_X1 U584 ( .A1(n529), .A2(n527), .ZN(n551) );
  NAND2_X1 U585 ( .A1(n551), .A2(n654), .ZN(n502) );
  XNOR2_X1 U586 ( .A(n535), .B(KEYINPUT6), .ZN(n563) );
  NOR2_X1 U587 ( .A1(n651), .A2(n653), .ZN(n506) );
  AND2_X1 U588 ( .A1(n563), .A2(n506), .ZN(n507) );
  XNOR2_X1 U589 ( .A(n508), .B(KEYINPUT32), .ZN(n509) );
  INV_X1 U590 ( .A(n651), .ZN(n585) );
  NOR2_X1 U591 ( .A1(n585), .A2(n535), .ZN(n510) );
  XNOR2_X1 U592 ( .A(KEYINPUT68), .B(n511), .ZN(n512) );
  NOR2_X2 U593 ( .A1(n727), .A2(n636), .ZN(n526) );
  INV_X1 U594 ( .A(KEYINPUT71), .ZN(n513) );
  NAND2_X1 U595 ( .A1(n526), .A2(n513), .ZN(n515) );
  AND2_X1 U596 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n514) );
  INV_X1 U597 ( .A(KEYINPUT44), .ZN(n524) );
  INV_X1 U598 ( .A(n516), .ZN(n532) );
  INV_X1 U599 ( .A(n532), .ZN(n539) );
  XNOR2_X1 U600 ( .A(n520), .B(n519), .ZN(n530) );
  OR2_X1 U601 ( .A1(n524), .A2(n725), .ZN(n525) );
  XOR2_X1 U602 ( .A(n527), .B(KEYINPUT104), .Z(n528) );
  AND2_X1 U603 ( .A1(n529), .A2(n528), .ZN(n645) );
  XNOR2_X1 U604 ( .A(n645), .B(KEYINPUT106), .ZN(n589) );
  NOR2_X1 U605 ( .A1(n589), .A2(n642), .ZN(n669) );
  BUF_X1 U606 ( .A(n530), .Z(n531) );
  INV_X1 U607 ( .A(n535), .ZN(n656) );
  NAND2_X1 U608 ( .A1(n532), .A2(n661), .ZN(n534) );
  XNOR2_X1 U609 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n533) );
  XNOR2_X1 U610 ( .A(n534), .B(n533), .ZN(n646) );
  NOR2_X1 U611 ( .A1(n517), .A2(n535), .ZN(n537) );
  NAND2_X1 U612 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U613 ( .A1(n539), .A2(n538), .ZN(n632) );
  NOR2_X1 U614 ( .A1(n646), .A2(n632), .ZN(n540) );
  NOR2_X1 U615 ( .A1(n669), .A2(n540), .ZN(n542) );
  NOR2_X1 U616 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n541) );
  NOR2_X1 U617 ( .A1(n542), .A2(n541), .ZN(n547) );
  XNOR2_X1 U618 ( .A(KEYINPUT89), .B(n543), .ZN(n544) );
  NOR2_X1 U619 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U620 ( .A1(n651), .A2(n546), .ZN(n629) );
  INV_X1 U621 ( .A(n700), .ZN(n595) );
  INV_X1 U622 ( .A(KEYINPUT38), .ZN(n548) );
  NAND2_X1 U623 ( .A1(n642), .A2(n590), .ZN(n550) );
  NAND2_X1 U624 ( .A1(n343), .A2(n664), .ZN(n668) );
  INV_X1 U625 ( .A(n551), .ZN(n667) );
  NOR2_X1 U626 ( .A1(n668), .A2(n667), .ZN(n553) );
  XNOR2_X1 U627 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n552) );
  XNOR2_X1 U628 ( .A(n553), .B(n552), .ZN(n680) );
  NOR2_X1 U629 ( .A1(n653), .A2(n554), .ZN(n555) );
  NAND2_X1 U630 ( .A1(n654), .A2(n555), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT28), .B(n556), .Z(n557) );
  INV_X1 U632 ( .A(n572), .ZN(n559) );
  NOR2_X1 U633 ( .A1(n680), .A2(n559), .ZN(n561) );
  XNOR2_X1 U634 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n560) );
  XNOR2_X1 U635 ( .A(n561), .B(n560), .ZN(n731) );
  NAND2_X1 U636 ( .A1(n730), .A2(n731), .ZN(n562) );
  INV_X1 U637 ( .A(n563), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n564), .A2(n642), .ZN(n565) );
  NOR2_X1 U639 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U640 ( .A1(n567), .A2(n664), .ZN(n583) );
  XNOR2_X1 U641 ( .A(KEYINPUT36), .B(n568), .ZN(n569) );
  NAND2_X1 U642 ( .A1(n569), .A2(n585), .ZN(n570) );
  XNOR2_X1 U643 ( .A(n570), .B(KEYINPUT114), .ZN(n728) );
  INV_X1 U644 ( .A(n576), .ZN(n640) );
  NOR2_X1 U645 ( .A1(n669), .A2(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n640), .A2(n573), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n669), .A2(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n576), .A2(KEYINPUT47), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n392), .A2(n580), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT72), .B(KEYINPUT48), .Z(n581) );
  XNOR2_X1 U651 ( .A(n582), .B(n581), .ZN(n593) );
  XNOR2_X1 U652 ( .A(KEYINPUT108), .B(n583), .ZN(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U654 ( .A(KEYINPUT43), .B(n586), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT109), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n588), .A2(n497), .ZN(n649) );
  INV_X1 U657 ( .A(n649), .ZN(n591) );
  AND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n648) );
  NOR2_X1 U659 ( .A1(n591), .A2(n648), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n715) );
  INV_X1 U661 ( .A(n715), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n597) );
  INV_X1 U663 ( .A(KEYINPUT2), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n597), .B(n596), .ZN(n650) );
  NOR2_X2 U665 ( .A1(n650), .A2(n598), .ZN(n688) );
  NAND2_X1 U666 ( .A1(n688), .A2(G472), .ZN(n601) );
  XOR2_X1 U667 ( .A(KEYINPUT62), .B(n599), .Z(n600) );
  XNOR2_X1 U668 ( .A(n601), .B(n600), .ZN(n603) );
  INV_X1 U669 ( .A(G952), .ZN(n602) );
  INV_X1 U670 ( .A(n696), .ZN(n619) );
  NAND2_X1 U671 ( .A1(n603), .A2(n619), .ZN(n605) );
  XNOR2_X1 U672 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n605), .B(n604), .ZN(G57) );
  NAND2_X1 U674 ( .A1(n688), .A2(G210), .ZN(n610) );
  XNOR2_X1 U675 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n606) );
  XOR2_X1 U676 ( .A(n606), .B(KEYINPUT55), .Z(n607) );
  XNOR2_X1 U677 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n611), .A2(n619), .ZN(n614) );
  XNOR2_X1 U680 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(KEYINPUT88), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n614), .B(n613), .ZN(G51) );
  NAND2_X1 U683 ( .A1(n688), .A2(G475), .ZN(n618) );
  XNOR2_X1 U684 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U686 ( .A(n618), .B(n617), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n622) );
  XNOR2_X1 U688 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n621) );
  XNOR2_X1 U689 ( .A(n622), .B(n621), .ZN(G60) );
  NAND2_X1 U690 ( .A1(n692), .A2(G469), .ZN(n626) );
  XNOR2_X1 U691 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X1 U694 ( .A1(n627), .A2(n696), .ZN(G54) );
  XOR2_X1 U695 ( .A(G101), .B(KEYINPUT115), .Z(n628) );
  XNOR2_X1 U696 ( .A(n629), .B(n628), .ZN(G3) );
  NAND2_X1 U697 ( .A1(n632), .A2(n642), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n630), .B(KEYINPUT116), .ZN(n631) );
  XNOR2_X1 U699 ( .A(G104), .B(n631), .ZN(G6) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n634) );
  NAND2_X1 U701 ( .A1(n632), .A2(n645), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U703 ( .A(G107), .B(n635), .ZN(G9) );
  XNOR2_X1 U704 ( .A(G110), .B(n636), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n637), .B(KEYINPUT117), .ZN(G12) );
  XOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .Z(n639) );
  NAND2_X1 U707 ( .A1(n640), .A2(n645), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n639), .B(n638), .ZN(G30) );
  NAND2_X1 U709 ( .A1(n640), .A2(n642), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n641), .B(G146), .ZN(G48) );
  NAND2_X1 U711 ( .A1(n646), .A2(n642), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(KEYINPUT118), .ZN(n644) );
  XNOR2_X1 U713 ( .A(G113), .B(n644), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(G116), .ZN(G18) );
  XOR2_X1 U716 ( .A(G134), .B(n648), .Z(G36) );
  XNOR2_X1 U717 ( .A(G140), .B(n649), .ZN(G42) );
  INV_X1 U718 ( .A(n650), .ZN(n686) );
  NAND2_X1 U719 ( .A1(n651), .A2(n517), .ZN(n652) );
  XOR2_X1 U720 ( .A(KEYINPUT50), .B(n652), .Z(n659) );
  NOR2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n655), .B(KEYINPUT49), .ZN(n657) );
  NAND2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U726 ( .A(KEYINPUT51), .B(n662), .Z(n663) );
  NOR2_X1 U727 ( .A1(n680), .A2(n663), .ZN(n676) );
  NOR2_X1 U728 ( .A1(n343), .A2(n664), .ZN(n665) );
  XOR2_X1 U729 ( .A(KEYINPUT119), .B(n665), .Z(n666) );
  NOR2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U732 ( .A1(n671), .A2(n670), .ZN(n674) );
  BUF_X1 U733 ( .A(n672), .Z(n673) );
  NOR2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U736 ( .A(n677), .B(KEYINPUT52), .ZN(n678) );
  NOR2_X1 U737 ( .A1(n679), .A2(n678), .ZN(n682) );
  NOR2_X1 U738 ( .A1(n680), .A2(n673), .ZN(n681) );
  NOR2_X1 U739 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n683), .B(KEYINPUT120), .ZN(n684) );
  NAND2_X1 U741 ( .A1(n684), .A2(n716), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U743 ( .A(n687), .B(KEYINPUT53), .ZN(G75) );
  AND2_X1 U744 ( .A1(n688), .A2(G478), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U746 ( .A1(n696), .A2(n691), .ZN(G63) );
  NAND2_X1 U747 ( .A1(n692), .A2(G217), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U749 ( .A1(n696), .A2(n695), .ZN(G66) );
  NAND2_X1 U750 ( .A1(G953), .A2(G224), .ZN(n697) );
  XOR2_X1 U751 ( .A(KEYINPUT61), .B(n697), .Z(n698) );
  NOR2_X1 U752 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U753 ( .A1(G953), .A2(n700), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(n709) );
  XOR2_X1 U755 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n707) );
  XOR2_X1 U756 ( .A(G101), .B(n703), .Z(n705) );
  NAND2_X1 U757 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n709), .B(n708), .ZN(G69) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U761 ( .A(n713), .B(n712), .Z(n718) );
  XOR2_X1 U762 ( .A(n718), .B(KEYINPUT125), .Z(n714) );
  XNOR2_X1 U763 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U764 ( .A1(n717), .A2(n716), .ZN(n724) );
  XNOR2_X1 U765 ( .A(n718), .B(G227), .ZN(n719) );
  XNOR2_X1 U766 ( .A(n719), .B(KEYINPUT126), .ZN(n720) );
  NAND2_X1 U767 ( .A1(n720), .A2(G900), .ZN(n721) );
  XOR2_X1 U768 ( .A(KEYINPUT127), .B(n721), .Z(n722) );
  NAND2_X1 U769 ( .A1(G953), .A2(n722), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n724), .A2(n723), .ZN(G72) );
  BUF_X1 U771 ( .A(n725), .Z(n726) );
  XNOR2_X1 U772 ( .A(n726), .B(G122), .ZN(G24) );
  XOR2_X1 U773 ( .A(G119), .B(n727), .Z(G21) );
  XOR2_X1 U774 ( .A(n728), .B(G125), .Z(n729) );
  XNOR2_X1 U775 ( .A(KEYINPUT37), .B(n729), .ZN(G27) );
  XNOR2_X1 U776 ( .A(G131), .B(n730), .ZN(G33) );
  XNOR2_X1 U777 ( .A(G137), .B(n731), .ZN(G39) );
endmodule

