//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n442, new_n443, new_n444, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G237));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n442));
  OR2_X1    g017(.A1(new_n442), .A2(G108), .ZN(new_n443));
  NAND2_X1  g018(.A1(new_n442), .A2(G108), .ZN(new_n444));
  NAND2_X1  g019(.A1(new_n443), .A2(new_n444), .ZN(G238));
  NAND4_X1  g020(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g028(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n440), .A2(G120), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n443), .A2(new_n444), .A3(G69), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(new_n458), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  OAI21_X1  g036(.A(G567), .B1(new_n456), .B2(new_n457), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G2106), .B1(KEYINPUT67), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G137), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n473), .B2(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n481), .B2(new_n472), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n485), .A3(G125), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n479), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  INV_X1    g063(.A(new_n472), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n478), .B1(new_n482), .B2(new_n490), .ZN(G160));
  NAND2_X1  g066(.A1(new_n483), .A2(new_n485), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n473), .A2(KEYINPUT70), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G136), .A4(new_n468), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n494), .A2(new_n495), .A3(new_n489), .A4(G124), .ZN(new_n500));
  OAI221_X1 g075(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n472), .C2(G112), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(G162));
  NAND3_X1  g078(.A1(new_n472), .A2(new_n473), .A3(G138), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  XOR2_X1   g082(.A(KEYINPUT72), .B(G114), .Z(new_n508));
  OAI211_X1 g083(.A(G2104), .B(new_n507), .C1(new_n508), .C2(new_n468), .ZN(new_n509));
  INV_X1    g084(.A(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n469), .B2(new_n471), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(KEYINPUT4), .B1(G126), .B2(G2105), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n506), .B(new_n509), .C1(new_n512), .C2(new_n492), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT74), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n517), .A2(new_n519), .B1(new_n516), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(G62), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT75), .Z(new_n529));
  NAND3_X1  g104(.A1(new_n524), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT6), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n525), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(G543), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(G88), .B1(new_n540), .B2(G50), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n530), .A2(KEYINPUT76), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n533), .A2(new_n541), .A3(new_n542), .ZN(G303));
  INV_X1    g118(.A(G303), .ZN(G166));
  NAND2_X1  g119(.A1(new_n540), .A2(G51), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n525), .A2(G89), .A3(new_n538), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  AOI22_X1  g129(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n534), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n525), .A2(new_n538), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n538), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT78), .B(G52), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n556), .A2(new_n561), .ZN(G171));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n557), .A2(new_n563), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n525), .A2(G56), .ZN(new_n566));
  NAND2_X1  g141(.A1(G68), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n534), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n538), .A2(G53), .A3(G543), .A4(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n535), .A2(new_n537), .A3(G53), .A4(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n580), .A2(new_n576), .A3(KEYINPUT9), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n579), .B1(new_n578), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G65), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n522), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(new_n539), .B2(G91), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G299));
  OR2_X1    g164(.A1(new_n556), .A2(new_n561), .ZN(G301));
  OAI21_X1  g165(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(KEYINPUT81), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n539), .A2(G87), .B1(new_n540), .B2(G49), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(KEYINPUT81), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND4_X1  g170(.A1(new_n535), .A2(new_n537), .A3(G48), .A4(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n525), .A2(G86), .A3(new_n538), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n599), .C1(new_n534), .C2(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n534), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n557), .A2(new_n604), .B1(new_n559), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT83), .B1(new_n557), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n525), .A2(new_n612), .A3(G92), .A4(new_n538), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n522), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(G54), .B2(new_n540), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n611), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n616), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(new_n583), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n578), .A2(new_n581), .A3(new_n579), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n587), .A2(G651), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n539), .A2(G91), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(G868), .B2(new_n633), .ZN(G297));
  OAI21_X1  g209(.A(new_n626), .B1(G868), .B2(new_n633), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n623), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n623), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g216(.A1(new_n494), .A2(new_n495), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n642), .A2(KEYINPUT85), .A3(G135), .A4(new_n468), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(G123), .A3(new_n489), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n472), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n494), .A2(new_n495), .A3(G135), .A4(new_n468), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n643), .A2(new_n644), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  INV_X1    g229(.A(G2100), .ZN(new_n655));
  AOI22_X1  g230(.A1(new_n653), .A2(new_n654), .B1(KEYINPUT84), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n473), .A2(new_n476), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT12), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(KEYINPUT84), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT13), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n656), .B(new_n661), .C1(new_n654), .C2(new_n653), .ZN(G156));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2427), .B(G2430), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT14), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n667), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2451), .B(G2454), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT16), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2443), .B(G2446), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1341), .B(G1348), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n672), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n683), .A3(G14), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT88), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n679), .A2(new_n683), .A3(new_n686), .A4(G14), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G401));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT89), .ZN(new_n691));
  XOR2_X1   g266(.A(G2084), .B(G2090), .Z(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2072), .B(G2078), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(KEYINPUT17), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n695), .A2(KEYINPUT17), .ZN(new_n698));
  AOI211_X1 g273(.A(new_n693), .B(new_n697), .C1(new_n698), .C2(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n695), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT18), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G2096), .B(G2100), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G227));
  XOR2_X1   g279(.A(G1956), .B(G2474), .Z(new_n705));
  XOR2_X1   g280(.A(G1961), .B(G1966), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1971), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT19), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(new_n706), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n708), .A2(new_n710), .A3(new_n712), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n715), .B(new_n716), .C1(new_n714), .C2(new_n713), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(G1991), .B(G1996), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1981), .ZN(new_n721));
  INV_X1    g296(.A(G1986), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n719), .B(new_n723), .ZN(G229));
  OAI21_X1  g299(.A(KEYINPUT91), .B1(G29), .B2(G33), .ZN(new_n725));
  OR3_X1    g300(.A1(KEYINPUT91), .A2(G29), .A3(G33), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n494), .A2(new_n495), .A3(G139), .A4(new_n468), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(new_n472), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n725), .B(new_n726), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G2072), .Z(new_n737));
  INV_X1    g312(.A(G1348), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n623), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G4), .B2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(G29), .A2(G32), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n642), .A2(G129), .A3(new_n489), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n476), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  NAND4_X1  g321(.A1(new_n494), .A2(new_n495), .A3(G141), .A4(new_n468), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n743), .A2(new_n744), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n742), .B1(new_n748), .B2(new_n735), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT24), .A2(G34), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n752), .A2(new_n735), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G160), .B2(new_n735), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(G2084), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G28), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n758), .A2(new_n759), .A3(new_n735), .ZN(new_n760));
  NOR2_X1   g335(.A1(G5), .A2(G16), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G171), .B2(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G1961), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n751), .A2(new_n756), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G16), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n765), .A2(KEYINPUT23), .A3(G20), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT23), .ZN(new_n767));
  INV_X1    g342(.A(G20), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G16), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n769), .C1(new_n633), .C2(new_n765), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n764), .B(new_n771), .C1(G2084), .C2(new_n755), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  NAND2_X1  g348(.A1(G164), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G27), .B2(G29), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n741), .B(new_n772), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(new_n773), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G21), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G168), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT94), .B(G1966), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n740), .A2(new_n738), .B1(new_n782), .B2(G11), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n782), .B2(G11), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n765), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n569), .B2(new_n765), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1341), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n749), .A2(new_n750), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT93), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n762), .A2(G1961), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT28), .ZN(new_n791));
  INV_X1    g366(.A(G26), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G29), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(G29), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n494), .A2(new_n495), .A3(new_n489), .A4(G128), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n494), .A2(new_n495), .A3(G140), .A4(new_n468), .ZN(new_n796));
  OAI221_X1 g371(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n472), .C2(G116), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n798), .B2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(new_n791), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n790), .B(new_n801), .C1(G29), .C2(new_n653), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n784), .A2(new_n787), .A3(new_n789), .A4(new_n802), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n776), .A2(new_n777), .A3(new_n781), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n735), .A2(G35), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n735), .ZN(new_n806));
  MUX2_X1   g381(.A(new_n805), .B(new_n806), .S(KEYINPUT95), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT97), .B(G2090), .Z(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n807), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n765), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n765), .ZN(new_n813));
  INV_X1    g388(.A(G1971), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n765), .A2(G6), .ZN(new_n816));
  INV_X1    g391(.A(G305), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n765), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT90), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n765), .A2(G23), .ZN(new_n823));
  INV_X1    g398(.A(G288), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n765), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1976), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT34), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G1976), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n827), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n831), .A2(new_n832), .A3(new_n815), .A4(new_n821), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n765), .A2(G24), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n607), .B2(new_n765), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n722), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n494), .A2(new_n495), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(new_n472), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G119), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(G2105), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G131), .ZN(new_n841));
  OAI221_X1 g416(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n472), .C2(G107), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  MUX2_X1   g418(.A(G25), .B(new_n843), .S(G29), .Z(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT35), .B(G1991), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n844), .B(new_n845), .Z(new_n846));
  NAND4_X1  g421(.A1(new_n829), .A2(new_n833), .A3(new_n836), .A4(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT36), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(KEYINPUT36), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n804), .B(new_n811), .C1(new_n848), .C2(new_n849), .ZN(G150));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  NAND2_X1  g426(.A1(G150), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n847), .B(KEYINPUT36), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n853), .A2(KEYINPUT98), .A3(new_n804), .A4(new_n811), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G311));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n557), .A2(new_n856), .B1(new_n559), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n525), .A2(G67), .ZN(new_n859));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n534), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(G860), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT37), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n623), .A2(G559), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  INV_X1    g440(.A(new_n565), .ZN(new_n866));
  INV_X1    g441(.A(new_n568), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n866), .B(new_n867), .C1(new_n861), .C2(new_n858), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n539), .A2(G93), .B1(new_n540), .B2(G55), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n859), .A2(new_n860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G651), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n869), .B(new_n871), .C1(new_n568), .C2(new_n565), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT39), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n865), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n863), .B1(new_n875), .B2(G860), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT99), .Z(G145));
  XOR2_X1   g452(.A(new_n843), .B(new_n658), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n652), .A2(G160), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n838), .A2(G123), .B1(new_n645), .B2(new_n647), .ZN(new_n881));
  INV_X1    g456(.A(new_n478), .ZN(new_n882));
  AOI211_X1 g457(.A(KEYINPUT69), .B(new_n472), .C1(new_n486), .C2(new_n479), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n881), .A2(new_n885), .A3(new_n651), .A4(new_n643), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n886), .A3(G162), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G162), .B1(new_n880), .B2(new_n886), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND4_X1   g465(.A1(new_n743), .A2(new_n744), .A3(new_n746), .A4(new_n747), .ZN(new_n891));
  NAND2_X1  g466(.A1(G164), .A2(new_n798), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n513), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(G164), .A2(new_n798), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n513), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n748), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n734), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n898), .A2(new_n733), .A3(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n890), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n838), .A2(G130), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT100), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n840), .A2(G142), .ZN(new_n904));
  OAI221_X1 g479(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n472), .C2(G118), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(KEYINPUT100), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n880), .A2(new_n886), .ZN(new_n911));
  INV_X1    g486(.A(G162), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n887), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n898), .A2(new_n895), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n733), .B(KEYINPUT92), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n898), .A2(new_n733), .A3(new_n895), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n901), .A2(new_n910), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n910), .B1(new_n901), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n879), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n890), .A2(new_n899), .A3(new_n900), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n914), .B1(new_n918), .B2(new_n917), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n901), .A2(new_n910), .A3(new_n919), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n878), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT103), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n922), .A2(new_n927), .A3(new_n931), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g509(.A(new_n638), .B(new_n873), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n622), .A2(new_n633), .ZN(new_n936));
  NAND4_X1  g511(.A1(G299), .A2(new_n620), .A3(new_n621), .A4(new_n616), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT41), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n942), .B2(new_n935), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n530), .A2(KEYINPUT76), .A3(G651), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT76), .B1(new_n530), .B2(G651), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n817), .B1(new_n947), .B2(new_n541), .ZN(new_n948));
  AND4_X1   g523(.A1(new_n541), .A2(new_n533), .A3(new_n542), .A4(new_n817), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n541), .A3(new_n817), .ZN(new_n951));
  NAND2_X1  g526(.A1(G303), .A2(G305), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT105), .ZN(new_n953));
  NAND2_X1  g528(.A1(G290), .A2(KEYINPUT104), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n607), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n824), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(G288), .A3(new_n956), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n950), .A2(new_n953), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n948), .A2(new_n949), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n962), .A2(KEYINPUT105), .A3(new_n959), .A4(new_n958), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n943), .B(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n966));
  AND2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(G868), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n858), .A2(new_n861), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n969), .B1(G868), .B2(new_n970), .ZN(G295));
  OAI21_X1  g546(.A(new_n969), .B1(G868), .B2(new_n970), .ZN(G331));
  OAI21_X1  g547(.A(KEYINPUT107), .B1(new_n556), .B2(new_n561), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n873), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n976));
  AOI21_X1  g551(.A(G286), .B1(new_n976), .B2(G171), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n868), .A2(new_n872), .A3(new_n973), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n549), .B(new_n552), .C1(G301), .C2(KEYINPUT107), .ZN(new_n980));
  INV_X1    g555(.A(new_n978), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n973), .B1(new_n868), .B2(new_n872), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n979), .B(new_n983), .C1(new_n939), .C2(new_n938), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n981), .A2(new_n982), .A3(new_n980), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n977), .B1(new_n975), .B2(new_n978), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n941), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(KEYINPUT108), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n964), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n928), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n964), .B2(new_n992), .ZN(new_n993));
  NOR4_X1   g568(.A1(new_n991), .A2(new_n993), .A3(KEYINPUT109), .A4(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n964), .A2(new_n992), .ZN(new_n995));
  INV_X1    g570(.A(new_n988), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n928), .A4(new_n990), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n964), .A2(new_n988), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n961), .A2(new_n963), .A3(new_n984), .A4(new_n987), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n928), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1003), .B2(KEYINPUT43), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n994), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n991), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n998), .B1(new_n1008), .B2(new_n997), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1009), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(G397));
  OAI211_X1 g590(.A(G40), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT111), .B1(G160), .B2(G40), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n513), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G2067), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n798), .B(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n748), .B(G1996), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT112), .Z(new_n1032));
  NOR2_X1   g607(.A1(new_n843), .A2(new_n845), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n893), .A2(new_n1027), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1026), .A2(new_n1037), .A3(G1996), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1025), .B1(new_n748), .B2(new_n1029), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1026), .B2(G1996), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n1041), .B(KEYINPUT47), .Z(new_n1042));
  AND2_X1   g617(.A1(new_n843), .A2(new_n845), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1025), .B1(new_n1033), .B2(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1032), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G290), .A2(G1986), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1025), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT126), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT48), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1036), .B(new_n1042), .C1(new_n1045), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G160), .A2(KEYINPUT111), .A3(G40), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1022), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  AND3_X1   g634(.A1(G305), .A2(new_n1059), .A3(G1981), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(G305), .B2(G1981), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1056), .B(new_n1058), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1056), .B1(G305), .B2(G1981), .ZN(new_n1064));
  NAND3_X1  g639(.A1(G305), .A2(new_n1059), .A3(G1981), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1055), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n830), .A3(new_n824), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1058), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1055), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n824), .A2(G1976), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n830), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1055), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n513), .A2(new_n1021), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1076), .A2(G8), .A3(new_n1071), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1067), .B(new_n1073), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT116), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1055), .A2(new_n1071), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1067), .A4(new_n1073), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G303), .A2(G8), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1086), .B(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1024), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT113), .B1(new_n1020), .B2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT45), .B1(new_n513), .B2(new_n1021), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1074), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1971), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1022), .B(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1074), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(G2090), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1089), .B(G8), .C1(new_n1098), .C2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1070), .B1(new_n1085), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  OAI21_X1  g680(.A(G8), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1086), .B(new_n1087), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1079), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1075), .A2(new_n1099), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1022), .A2(KEYINPUT50), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT117), .B(G2084), .Z(new_n1113));
  AND4_X1   g688(.A1(new_n1074), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n780), .B1(new_n1095), .B2(new_n1074), .ZN(new_n1115));
  OAI211_X1 g690(.A(G8), .B(G168), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1105), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1116), .A2(new_n1105), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1103), .A3(new_n1108), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1104), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n780), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1020), .B2(new_n1091), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1074), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(G168), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G168), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n1127));
  OAI211_X1 g702(.A(G8), .B(new_n1125), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1114), .A2(new_n1115), .A3(G286), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT51), .B1(new_n1129), .B2(new_n1054), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1092), .A2(new_n773), .A3(new_n1097), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1961), .B1(new_n1100), .B2(new_n1074), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n882), .B(G40), .C1(new_n472), .C2(new_n481), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1138), .A2(KEYINPUT122), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1133), .A2(G2078), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(KEYINPUT122), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1139), .A2(new_n1095), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1134), .A2(G301), .A3(new_n1136), .A4(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1095), .A2(new_n1074), .A3(new_n1140), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1135), .B(new_n1145), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1146), .B2(G301), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1131), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT56), .B(G2072), .Z(new_n1150));
  OR3_X1    g725(.A1(new_n1020), .A2(new_n1091), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n584), .B2(new_n588), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n578), .A2(new_n581), .ZN(new_n1154));
  AND4_X1   g729(.A1(new_n1152), .A2(new_n630), .A3(new_n631), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT119), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT57), .B1(new_n629), .B2(new_n632), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n588), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT118), .B(G1956), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(new_n1020), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1151), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1053), .A2(new_n1027), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(G1348), .B1(new_n1100), .B2(new_n1074), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n623), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1095), .A2(new_n1074), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1171), .A2(new_n1150), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1162), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1100), .B2(new_n1074), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1170), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1169), .B1(new_n1175), .B2(KEYINPUT120), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1161), .B1(new_n1151), .B2(new_n1164), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1165), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1168), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1181), .A2(new_n623), .A3(new_n1166), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n622), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1182), .A2(new_n1183), .A3(KEYINPUT60), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1171), .A2(G1996), .ZN(new_n1185));
  XNOR2_X1  g760(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(G1341), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1053), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n569), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(KEYINPUT59), .B(new_n569), .C1(new_n1185), .C2(new_n1188), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT60), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1181), .A2(new_n1193), .A3(new_n623), .A4(new_n1166), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1184), .A2(new_n1191), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1165), .B1(new_n1177), .B2(KEYINPUT61), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1151), .A2(new_n1197), .A3(new_n1161), .A4(new_n1164), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1180), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1134), .A2(G301), .A3(new_n1136), .A4(new_n1144), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(KEYINPUT54), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1135), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1203));
  AOI21_X1  g778(.A(G301), .B1(new_n1203), .B2(new_n1142), .ZN(new_n1204));
  OAI21_X1  g779(.A(KEYINPUT124), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1142), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(G171), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1207), .A2(new_n1208), .A3(KEYINPUT54), .A4(new_n1201), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1149), .A2(new_n1200), .A3(new_n1205), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1110), .A2(KEYINPUT123), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1108), .A2(new_n1103), .A3(new_n1212), .A4(new_n1109), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1121), .B1(new_n1210), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1128), .A2(new_n1130), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(G301), .B1(new_n1203), .B2(new_n1144), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(KEYINPUT125), .B1(new_n1214), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n1223));
  AOI211_X1 g798(.A(new_n1223), .B(new_n1220), .C1(new_n1211), .C2(new_n1213), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  OR2_X1    g800(.A1(new_n1131), .A2(new_n1217), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1216), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n607), .A2(new_n722), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1025), .B1(new_n1046), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1045), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1050), .B1(new_n1227), .B2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n688), .A2(G319), .ZN(new_n1234));
  INV_X1    g808(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n933), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n1004), .A2(new_n999), .ZN(new_n1237));
  NAND4_X1  g811(.A1(new_n1008), .A2(new_n1000), .A3(new_n998), .A4(new_n997), .ZN(new_n1238));
  NOR2_X1   g812(.A1(G229), .A2(G227), .ZN(new_n1239));
  NAND3_X1  g813(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g814(.A(new_n1233), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g815(.A(new_n1234), .B1(new_n930), .B2(new_n932), .ZN(new_n1242));
  NAND4_X1  g816(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n1239), .A4(new_n1242), .ZN(new_n1243));
  AND2_X1   g817(.A1(new_n1241), .A2(new_n1243), .ZN(G308));
  NAND2_X1  g818(.A1(new_n1241), .A2(new_n1243), .ZN(G225));
endmodule


