//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n547, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n581,
    new_n582, new_n583, new_n586, new_n588, new_n589, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n453), .A2(G2106), .B1(KEYINPUT66), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  XOR2_X1   g040(.A(new_n465), .B(KEYINPUT67), .Z(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  OAI221_X1 g049(.A(new_n466), .B1(new_n472), .B2(new_n473), .C1(new_n474), .C2(new_n464), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n472), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n471), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n464), .B2(G112), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n468), .A3(new_n470), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n487), .A2(new_n468), .A3(new_n470), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(KEYINPUT71), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n489), .A2(new_n495), .A3(KEYINPUT4), .A4(new_n491), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(new_n464), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G102), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(new_n464), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n471), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n494), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n507), .A2(KEYINPUT72), .A3(KEYINPUT5), .A4(G543), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(KEYINPUT73), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(new_n510), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(KEYINPUT74), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(G88), .B1(G50), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n520), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n522), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n520), .A2(G90), .B1(G52), .B2(new_n522), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n516), .B2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(new_n520), .A2(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n521), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n516), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT76), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  NAND3_X1  g126(.A1(new_n519), .A2(G53), .A3(G543), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n520), .A2(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n553), .B(new_n554), .C1(new_n516), .C2(new_n555), .ZN(G299));
  NAND2_X1  g131(.A1(new_n520), .A2(G87), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n522), .A2(G49), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(G288));
  NAND2_X1  g135(.A1(new_n522), .A2(G48), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n514), .A2(new_n519), .A3(G86), .ZN(new_n562));
  NAND2_X1  g137(.A1(G73), .A2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT77), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n514), .B2(G61), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n561), .B(new_n562), .C1(new_n565), .C2(new_n516), .ZN(G305));
  AOI22_X1  g141(.A1(new_n520), .A2(G85), .B1(G47), .B2(new_n522), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT79), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT78), .Z(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n516), .B2(new_n570), .ZN(G290));
  NAND2_X1  g146(.A1(G301), .A2(G868), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n520), .A2(G92), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT10), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n522), .A2(G54), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n516), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n572), .B1(new_n578), .B2(G868), .ZN(G284));
  OAI21_X1  g154(.A(new_n572), .B1(new_n578), .B2(G868), .ZN(G321));
  NAND2_X1  g155(.A1(G286), .A2(G868), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT80), .Z(new_n582));
  INV_X1    g157(.A(G299), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(G868), .B2(new_n583), .ZN(G297));
  OAI21_X1  g159(.A(new_n582), .B1(G868), .B2(new_n583), .ZN(G280));
  INV_X1    g160(.A(G559), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n578), .B1(new_n586), .B2(G860), .ZN(G148));
  NAND2_X1  g162(.A1(new_n578), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G868), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g165(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g166(.A(G135), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n472), .A2(KEYINPUT82), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n479), .A2(G123), .ZN(new_n594));
  OR2_X1    g169(.A1(G99), .A2(G2105), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n595), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n472), .B2(new_n592), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(G2096), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT12), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT13), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT81), .B(G2100), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n598), .A2(G2096), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g182(.A(KEYINPUT15), .B(G2430), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2435), .ZN(new_n609));
  XOR2_X1   g184(.A(G2427), .B(G2438), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT14), .ZN(new_n612));
  XNOR2_X1  g187(.A(G2443), .B(G2446), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2451), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2454), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n612), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(G1341), .B(G1348), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n618), .B(new_n619), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G14), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(G401));
  XOR2_X1   g197(.A(G2072), .B(G2078), .Z(new_n623));
  XOR2_X1   g198(.A(G2067), .B(G2678), .Z(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G2084), .B(G2090), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n623), .B1(new_n627), .B2(KEYINPUT18), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2096), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2100), .Z(new_n630));
  AND2_X1   g205(.A1(new_n627), .A2(KEYINPUT17), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n625), .A2(new_n626), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT18), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(G227));
  XOR2_X1   g209(.A(G1956), .B(G2474), .Z(new_n635));
  XOR2_X1   g210(.A(G1961), .B(G1966), .Z(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1971), .B(G1976), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT19), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(new_n636), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n640), .A3(new_n642), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n645), .B(new_n646), .C1(new_n644), .C2(new_n643), .ZN(new_n647));
  XOR2_X1   g222(.A(G1991), .B(G1996), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1981), .B(G1986), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n651), .B(new_n653), .Z(G229));
  INV_X1    g229(.A(KEYINPUT28), .ZN(new_n655));
  INV_X1    g230(.A(G26), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n655), .B1(new_n656), .B2(G29), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(G29), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n477), .A2(G140), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n479), .A2(G128), .ZN(new_n660));
  NOR2_X1   g235(.A1(G104), .A2(G2105), .ZN(new_n661));
  OAI21_X1  g236(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n659), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n658), .B1(new_n663), .B2(G29), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n657), .B1(new_n664), .B2(new_n655), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(G2067), .ZN(new_n666));
  INV_X1    g241(.A(G16), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n544), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n667), .B2(G19), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(G1341), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(G1341), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(G2067), .ZN(new_n673));
  AND4_X1   g248(.A1(new_n666), .A2(new_n671), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(KEYINPUT93), .B1(G5), .B2(G16), .ZN(new_n675));
  OR3_X1    g250(.A1(KEYINPUT93), .A2(G5), .A3(G16), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(G301), .C2(new_n667), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT94), .B(G1961), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  AOI22_X1  g254(.A1(G141), .A2(new_n477), .B1(new_n479), .B2(G129), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n681));
  NAND3_X1  g256(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT26), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G29), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G29), .B2(G32), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT27), .B(G1996), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n679), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(KEYINPUT90), .B1(G4), .B2(G16), .ZN(new_n691));
  OR3_X1    g266(.A1(KEYINPUT90), .A2(G4), .A3(G16), .ZN(new_n692));
  INV_X1    g267(.A(new_n578), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n667), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1348), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G21), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G168), .B2(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(G1966), .ZN(new_n698));
  INV_X1    g273(.A(new_n598), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G29), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT92), .B(G28), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT30), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  INV_X1    g278(.A(G34), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(KEYINPUT24), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(KEYINPUT24), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G160), .B2(new_n703), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n700), .B1(G29), .B2(new_n702), .C1(new_n708), .C2(G2084), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n698), .B(new_n709), .C1(G2084), .C2(new_n708), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n674), .A2(new_n690), .A3(new_n695), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n703), .A2(G35), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G162), .B2(new_n703), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT29), .Z(new_n714));
  INV_X1    g289(.A(G2090), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n688), .B2(new_n689), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n714), .A2(new_n715), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  INV_X1    g295(.A(G139), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n720), .B1(new_n472), .B2(new_n721), .C1(new_n722), .C2(new_n464), .ZN(new_n723));
  MUX2_X1   g298(.A(G33), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G2072), .Z(new_n725));
  INV_X1    g300(.A(G1966), .ZN(new_n726));
  INV_X1    g301(.A(new_n697), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n711), .A2(new_n717), .A3(new_n718), .A4(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n667), .A2(G24), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G290), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT87), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1986), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n667), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n667), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1971), .ZN(new_n736));
  NOR2_X1   g311(.A1(G6), .A2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G305), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT32), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1981), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G23), .ZN(new_n742));
  INV_X1    g317(.A(G288), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT33), .B(G1976), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n744), .B(new_n745), .Z(new_n746));
  NOR3_X1   g321(.A1(new_n736), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT34), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(new_n464), .B2(G107), .ZN(new_n750));
  INV_X1    g325(.A(G95), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n464), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT86), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n479), .A2(G119), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n477), .A2(G131), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G25), .B(new_n756), .S(G29), .Z(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT35), .B(G1991), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n757), .B(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n733), .A2(new_n749), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT88), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n748), .B2(new_n747), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT89), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n729), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(KEYINPUT89), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n766), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n703), .A2(G27), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n703), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n667), .A2(G20), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT95), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n583), .B2(new_n667), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT96), .B(G1956), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n769), .A2(new_n770), .A3(new_n774), .A4(new_n780), .ZN(G150));
  INV_X1    g356(.A(G150), .ZN(G311));
  AOI22_X1  g357(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n516), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n522), .A2(G55), .ZN(new_n786));
  INV_X1    g361(.A(new_n520), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT98), .B(G93), .Z(new_n788));
  OAI211_X1 g363(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G860), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT37), .Z(new_n791));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n792), .B2(new_n544), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n792), .B2(new_n544), .ZN(new_n794));
  INV_X1    g369(.A(new_n544), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n789), .A2(KEYINPUT99), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n578), .A2(G559), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT39), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n799), .B(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n791), .B1(new_n802), .B2(G860), .ZN(G145));
  XNOR2_X1  g378(.A(new_n484), .B(new_n475), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(new_n699), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(new_n601), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(new_n756), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n685), .B(new_n663), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(new_n505), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n723), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n723), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n477), .A2(G142), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n479), .A2(G130), .ZN(new_n814));
  NOR2_X1   g389(.A1(G106), .A2(G2105), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n812), .B(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n811), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n807), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G37), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g398(.A1(new_n789), .A2(G868), .ZN(new_n824));
  XNOR2_X1  g399(.A(G303), .B(new_n743), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G290), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G305), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT42), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(KEYINPUT102), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT102), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n797), .B(new_n588), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n578), .B(G299), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n834), .B(KEYINPUT41), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n831), .A2(new_n832), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n832), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n831), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n824), .B1(new_n841), .B2(G868), .ZN(G295));
  AOI21_X1  g417(.A(new_n824), .B1(new_n841), .B2(G868), .ZN(G331));
  XNOR2_X1  g418(.A(G301), .B(G286), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n797), .B(new_n844), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n834), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n797), .B(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n836), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n849), .A2(KEYINPUT104), .A3(new_n827), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT104), .B1(new_n849), .B2(new_n827), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n821), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n845), .A2(new_n834), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n846), .A2(KEYINPUT105), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(new_n827), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n852), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n849), .A2(new_n827), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n850), .A2(new_n821), .A3(new_n851), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT44), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(KEYINPUT43), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n852), .A2(new_n858), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n867), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g443(.A(KEYINPUT125), .ZN(new_n869));
  INV_X1    g444(.A(G40), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n475), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G1384), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT50), .B1(new_n505), .B2(new_n872), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n715), .B(new_n871), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n871), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT45), .B1(new_n505), .B2(new_n872), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT106), .B(G1384), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT108), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT108), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n505), .A2(new_n881), .A3(KEYINPUT45), .A4(new_n878), .ZN(new_n882));
  AOI211_X1 g457(.A(new_n876), .B(new_n877), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(KEYINPUT115), .B(new_n875), .C1(new_n883), .C2(G1971), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT115), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n877), .A2(new_n876), .ZN(new_n887));
  AOI21_X1  g462(.A(G1971), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n875), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(KEYINPUT110), .B(G8), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(G303), .A2(G8), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n871), .A2(new_n872), .A3(new_n505), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n743), .A2(G1976), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n891), .ZN(new_n899));
  NAND2_X1  g474(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n743), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n897), .A2(new_n898), .A3(new_n891), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n897), .A2(new_n891), .ZN(new_n906));
  NAND2_X1  g481(.A1(G305), .A2(KEYINPUT49), .ZN(new_n907));
  INV_X1    g482(.A(G1981), .ZN(new_n908));
  INV_X1    g483(.A(G61), .ZN(new_n909));
  OAI21_X1  g484(.A(G543), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n512), .B2(new_n510), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n911), .B2(new_n508), .ZN(new_n912));
  OAI21_X1  g487(.A(G651), .B1(new_n912), .B2(new_n564), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n908), .B1(new_n913), .B2(KEYINPUT112), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT49), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n913), .A2(new_n915), .A3(new_n561), .A4(new_n562), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n907), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n914), .B1(new_n907), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n906), .A2(new_n919), .A3(KEYINPUT113), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT113), .B1(new_n906), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n905), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(G8), .B1(new_n888), .B2(new_n889), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n895), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n896), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT119), .B(G2072), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT56), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n886), .A2(new_n887), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n932));
  INV_X1    g507(.A(G1956), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT57), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n583), .A2(KEYINPUT118), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT118), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT57), .B1(G299), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n931), .A2(new_n934), .A3(new_n940), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(KEYINPUT61), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT121), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n942), .A2(new_n946), .A3(KEYINPUT61), .A4(new_n943), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n886), .A2(new_n887), .ZN(new_n949));
  INV_X1    g524(.A(new_n897), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT58), .B(G1341), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n949), .A2(G1996), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n544), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT60), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n505), .A2(new_n872), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n872), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n876), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n960), .A2(G1348), .B1(G2067), .B2(new_n897), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n578), .ZN(new_n962));
  INV_X1    g537(.A(G1348), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n932), .A2(new_n963), .B1(new_n964), .B2(new_n950), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n693), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n955), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT120), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n942), .A2(new_n968), .A3(new_n943), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n940), .B1(new_n931), .B2(new_n934), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT61), .B1(new_n970), .B2(KEYINPUT120), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n967), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n955), .A3(new_n578), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n948), .A2(new_n954), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n962), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n970), .B1(new_n975), .B2(new_n943), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n872), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n505), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n872), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n887), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n773), .A2(KEYINPUT53), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n886), .A2(new_n773), .A3(new_n887), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1961), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n932), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n985), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G171), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n876), .B1(new_n880), .B2(new_n882), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n505), .B2(new_n878), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n984), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n986), .A2(new_n987), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT123), .B1(new_n960), .B2(G1961), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT123), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n932), .A2(new_n999), .A3(new_n989), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n992), .B(new_n993), .C1(G171), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT124), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n1002), .B2(G171), .ZN(new_n1005));
  AOI211_X1 g580(.A(KEYINPUT124), .B(G301), .C1(new_n997), .C2(new_n1001), .ZN(new_n1006));
  AND4_X1   g581(.A1(G301), .A2(new_n985), .A3(new_n988), .A4(new_n990), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1003), .B1(new_n1008), .B2(new_n993), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1966), .B1(new_n982), .B2(new_n887), .ZN(new_n1010));
  INV_X1    g585(.A(G2084), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(new_n871), .C1(new_n873), .C2(new_n874), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n891), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n1015));
  INV_X1    g590(.A(new_n891), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G168), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT122), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n983), .A2(new_n726), .B1(new_n1011), .B2(new_n960), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT51), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1014), .A2(KEYINPUT122), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1017), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AND4_X1   g605(.A1(new_n928), .A2(new_n977), .A3(new_n1009), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(G168), .A3(new_n891), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n896), .A2(new_n1033), .A3(new_n926), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT63), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(KEYINPUT117), .A3(new_n1035), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n923), .B2(new_n895), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1033), .A2(new_n926), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n922), .A2(new_n923), .A3(new_n895), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n920), .A2(new_n921), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G288), .A2(G1976), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1044), .A2(new_n1045), .B1(new_n908), .B2(new_n738), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1043), .B1(new_n1048), .B2(new_n906), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n869), .B1(new_n1031), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n977), .A2(new_n1009), .A3(new_n928), .A4(new_n1030), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(KEYINPUT125), .A3(new_n1049), .A4(new_n1042), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT62), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1027), .A2(new_n1054), .A3(new_n1029), .ZN(new_n1055));
  INV_X1    g630(.A(new_n992), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n927), .B1(new_n1030), .B2(KEYINPUT62), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT126), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT126), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1051), .A2(new_n1053), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n995), .A2(new_n871), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(G290), .A2(G1986), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT107), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G290), .A2(G1986), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1996), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n686), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n663), .B(new_n964), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n685), .A2(G1996), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n756), .B(new_n759), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1064), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1062), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n756), .A2(new_n758), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n663), .A2(G2067), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1063), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1064), .B1(new_n1073), .B2(new_n685), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1064), .A2(KEYINPUT46), .A3(new_n1070), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT46), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1063), .B2(G1996), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(new_n1088), .B(KEYINPUT47), .Z(new_n1089));
  NAND2_X1  g664(.A1(new_n1077), .A2(new_n1064), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1065), .A2(new_n1063), .ZN(new_n1091));
  XOR2_X1   g666(.A(new_n1091), .B(KEYINPUT48), .Z(new_n1092));
  AOI211_X1 g667(.A(new_n1083), .B(new_n1089), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1079), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT127), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT127), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1079), .A2(new_n1096), .A3(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g673(.A(G229), .ZN(new_n1100));
  NAND2_X1  g674(.A1(new_n822), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g675(.A1(G227), .A2(new_n462), .ZN(new_n1102));
  NAND2_X1  g676(.A1(new_n621), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g677(.A1(new_n867), .A2(new_n1101), .A3(new_n1103), .ZN(G308));
  MUX2_X1   g678(.A(new_n862), .B(new_n866), .S(new_n859), .Z(new_n1105));
  INV_X1    g679(.A(new_n1101), .ZN(new_n1106));
  NAND4_X1  g680(.A1(new_n1105), .A2(new_n621), .A3(new_n1106), .A4(new_n1102), .ZN(G225));
endmodule


