//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G137), .A4(new_n461), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT70), .ZN(G160));
  AND3_X1   g050(.A1(new_n467), .A2(new_n469), .A3(new_n461), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n467), .A2(new_n469), .A3(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT71), .A2(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n461), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(new_n494), .A3(G138), .A4(new_n461), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT72), .B1(new_n498), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT73), .B1(new_n501), .B2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n498), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n503), .A2(new_n507), .A3(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n497), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n503), .A2(new_n507), .A3(G88), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(G50), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n510), .A2(new_n514), .ZN(G166));
  AOI22_X1  g090(.A1(new_n499), .A2(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(new_n511), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n511), .A2(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(G51), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n519), .A3(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(G90), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n497), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n497), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n516), .A2(new_n511), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n511), .A2(G543), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT75), .B(G43), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n520), .A2(new_n548), .A3(G53), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n550), .B1(new_n549), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n503), .A2(new_n507), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(G91), .A2(new_n517), .B1(new_n560), .B2(G651), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n555), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n556), .B1(new_n555), .B2(new_n561), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  NAND2_X1  g141(.A1(new_n508), .A2(new_n509), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n512), .A2(new_n513), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT78), .B1(new_n510), .B2(new_n514), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n503), .A2(new_n507), .A3(G87), .A4(new_n511), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n503), .A2(new_n507), .A3(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n520), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n503), .A2(new_n507), .A3(G86), .A4(new_n511), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n516), .A2(KEYINPUT79), .A3(G86), .A4(new_n511), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n581), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(KEYINPUT80), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(G651), .A3(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n517), .A2(G85), .B1(G47), .B2(new_n520), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n558), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n536), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n602), .A2(new_n605), .B1(G54), .B2(new_n520), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n594), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n594), .B1(new_n607), .B2(G868), .ZN(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n607), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n476), .A2(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n476), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n478), .A2(G123), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n461), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n623), .A3(new_n629), .ZN(G156));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n631), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g222(.A(KEYINPUT82), .B(new_n645), .C1(new_n642), .C2(new_n643), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n644), .B2(new_n646), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(KEYINPUT83), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT83), .B1(new_n649), .B2(new_n651), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n669), .A2(new_n670), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n678), .A2(new_n674), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n671), .A3(new_n674), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n683), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n690), .ZN(new_n693));
  INV_X1    g268(.A(new_n686), .ZN(new_n694));
  INV_X1    g269(.A(new_n687), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n684), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n693), .B1(new_n696), .B2(new_n688), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n692), .A2(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G23), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n575), .A2(new_n576), .ZN(new_n701));
  INV_X1    g276(.A(G74), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n497), .B1(new_n558), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(KEYINPUT87), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n574), .A2(new_n705), .A3(new_n575), .A4(new_n576), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n700), .B1(new_n708), .B2(new_n699), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT88), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT33), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n699), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n699), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n712), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n476), .A2(G131), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n478), .A2(G119), .ZN(new_n727));
  OR2_X1    g302(.A1(G95), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n724), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n591), .A2(new_n592), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G16), .B2(G24), .ZN(new_n737));
  INV_X1    g312(.A(G1986), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(new_n737), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n722), .A2(new_n723), .A3(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT36), .Z(new_n742));
  AND2_X1   g317(.A1(new_n699), .A2(G21), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G286), .B2(G16), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G33), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n476), .A2(G139), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n750), .B(new_n751), .C1(new_n461), .C2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n748), .B1(new_n753), .B2(new_n724), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G2072), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT30), .B(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n756), .A2(new_n724), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n628), .B2(new_n724), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n724), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n476), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n478), .A2(G128), .ZN(new_n764));
  OR2_X1    g339(.A1(G104), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n724), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  OR4_X1    g344(.A1(new_n746), .A2(new_n755), .A3(new_n760), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G164), .A2(new_n724), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G27), .B2(new_n724), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n745), .A2(new_n744), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n724), .A2(G32), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n476), .A2(G141), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n478), .A2(G129), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n471), .A2(G105), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n779), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n779), .B2(new_n783), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n775), .B1(new_n788), .B2(new_n724), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT27), .B(G1996), .Z(new_n790));
  OAI221_X1 g365(.A(new_n774), .B1(new_n773), .B2(new_n772), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n724), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n724), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT29), .Z(new_n794));
  INV_X1    g369(.A(G2090), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n541), .A2(new_n699), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n699), .B2(G19), .ZN(new_n798));
  INV_X1    g373(.A(G1341), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n699), .A2(G5), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G171), .B2(new_n699), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(G1961), .ZN(new_n803));
  NAND2_X1  g378(.A1(G160), .A2(G29), .ZN(new_n804));
  INV_X1    g379(.A(G34), .ZN(new_n805));
  AOI21_X1  g380(.A(G29), .B1(new_n805), .B2(KEYINPUT24), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(KEYINPUT24), .B2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G2084), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n796), .A2(new_n800), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n798), .A2(new_n799), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n770), .A2(new_n791), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n802), .A2(KEYINPUT95), .A3(G1961), .ZN(new_n814));
  AOI21_X1  g389(.A(KEYINPUT95), .B1(new_n802), .B2(G1961), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n789), .B2(new_n790), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(G299), .A2(G16), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n699), .A2(G20), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT23), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G1956), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n794), .A2(new_n795), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n823), .A2(KEYINPUT96), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n699), .A2(G4), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n607), .B2(new_n699), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT91), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT90), .B(G1348), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT89), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n817), .A2(new_n827), .A3(new_n828), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n742), .A2(new_n835), .ZN(G311));
  OR2_X1    g411(.A1(new_n742), .A2(new_n835), .ZN(G150));
  NAND2_X1  g412(.A1(new_n520), .A2(G55), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n536), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n516), .A2(G67), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n497), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT98), .B1(new_n840), .B2(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n607), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n535), .A2(new_n540), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n846), .A2(new_n853), .A3(new_n847), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT97), .B1(new_n853), .B2(new_n844), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n541), .B(new_n856), .C1(new_n843), .C2(new_n840), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n858), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n861), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n866), .B2(KEYINPUT39), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n864), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n850), .B1(new_n868), .B2(new_n869), .ZN(G145));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n753), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n788), .A2(new_n767), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n493), .A2(new_n495), .ZN(new_n875));
  AND2_X1   g450(.A1(KEYINPUT71), .A2(G114), .ZN(new_n876));
  NOR2_X1   g451(.A1(KEYINPUT71), .A2(G114), .ZN(new_n877));
  OAI21_X1  g452(.A(G2105), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n490), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n478), .A2(G126), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT101), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n875), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n767), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n787), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n874), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n874), .B2(new_n888), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n873), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n753), .A2(new_n871), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n889), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n478), .A2(G130), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n461), .A2(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(G142), .B2(new_n476), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n619), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n731), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n892), .A2(new_n895), .A3(new_n903), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G160), .B(new_n628), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(G162), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(KEYINPUT103), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n892), .A2(new_n895), .A3(new_n912), .A4(new_n903), .ZN(new_n913));
  INV_X1    g488(.A(new_n909), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n911), .A2(new_n905), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g492(.A1(new_n848), .A2(G868), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n735), .A2(new_n708), .ZN(new_n919));
  NAND2_X1  g494(.A1(G290), .A2(new_n707), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(KEYINPUT105), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(G166), .A2(KEYINPUT104), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n510), .B2(new_n514), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(G305), .Z(new_n926));
  NOR2_X1   g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n921), .A2(new_n926), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n919), .A2(new_n920), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n927), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT42), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n601), .A2(new_n606), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n563), .A2(new_n935), .A3(new_n564), .ZN(new_n936));
  INV_X1    g511(.A(new_n554), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n551), .B(new_n548), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n550), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n941));
  INV_X1    g516(.A(G91), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n941), .A2(new_n497), .B1(new_n942), .B2(new_n536), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT77), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n944), .A2(new_n562), .B1(new_n601), .B2(new_n606), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n934), .B1(new_n936), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n935), .B1(new_n563), .B2(new_n564), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n607), .A2(new_n944), .A3(new_n562), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n614), .B(new_n858), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n936), .A2(new_n945), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n952), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n933), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n931), .A2(new_n921), .A3(new_n926), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n921), .A2(new_n926), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n954), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n961), .A3(KEYINPUT106), .ZN(new_n962));
  OR3_X1    g537(.A1(new_n933), .A2(KEYINPUT106), .A3(new_n955), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n918), .B1(new_n964), .B2(G868), .ZN(G295));
  AOI21_X1  g540(.A(new_n918), .B1(new_n964), .B2(G868), .ZN(G331));
  NAND2_X1  g541(.A1(G171), .A2(G168), .ZN(new_n967));
  OAI21_X1  g542(.A(G286), .B1(new_n530), .B2(new_n532), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n858), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n968), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(new_n854), .A3(new_n857), .A4(new_n855), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n950), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n970), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n858), .A2(new_n969), .A3(KEYINPUT107), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n932), .B(new_n974), .C1(new_n978), .C2(new_n953), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n953), .B1(new_n976), .B2(new_n977), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n946), .A2(new_n949), .B1(new_n970), .B2(new_n972), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n959), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G37), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n980), .A2(new_n981), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n986), .B2(new_n932), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n936), .A2(new_n945), .A3(new_n934), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT41), .B1(new_n947), .B2(new_n948), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n976), .B(new_n977), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n947), .A2(new_n948), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n970), .A3(new_n993), .A4(new_n972), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT108), .B1(new_n973), .B2(new_n953), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n959), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n987), .A2(new_n988), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n985), .A2(new_n998), .A3(KEYINPUT109), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n987), .A2(new_n1001), .A3(new_n997), .A4(new_n988), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n987), .A2(new_n997), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1004), .B2(KEYINPUT43), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT110), .B1(new_n984), .B2(KEYINPUT43), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n987), .A2(new_n1007), .A3(new_n988), .A4(new_n982), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1003), .A2(new_n1009), .ZN(G397));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n571), .A2(G8), .A3(new_n572), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n473), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n463), .A2(new_n464), .ZN(new_n1018));
  OAI211_X1 g593(.A(G40), .B(new_n1017), .C1(new_n1018), .C2(new_n461), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n881), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n1020), .A4(new_n884), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n718), .ZN(new_n1026));
  INV_X1    g601(.A(G40), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n465), .A2(new_n473), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n875), .B2(new_n880), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g606(.A(KEYINPUT50), .B(G1384), .C1(new_n875), .C2(new_n880), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1031), .A2(G2090), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1016), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n704), .A2(G1976), .A3(new_n706), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .A4(KEYINPUT52), .ZN(new_n1044));
  NOR2_X1   g619(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G288), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  INV_X1    g623(.A(G1981), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n581), .A2(new_n1049), .A3(new_n586), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n581), .B2(new_n582), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n520), .A2(G48), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n582), .B(new_n1053), .C1(new_n1054), .C2(new_n497), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G1981), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n581), .A2(new_n1049), .A3(new_n586), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT49), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(new_n1058), .A3(new_n1039), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1047), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1011), .B1(new_n1036), .B2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1040), .A2(new_n1042), .B1(G288), .B2(new_n1045), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1039), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(new_n1048), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1062), .A2(new_n1044), .B1(new_n1065), .B2(new_n1058), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1971), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n1067), .B2(new_n1033), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1070), .A3(KEYINPUT116), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT63), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n881), .A2(new_n1030), .A3(new_n1020), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n809), .A3(new_n1074), .A4(new_n1028), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1019), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n809), .A4(new_n1074), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1028), .B1(new_n1029), .B2(KEYINPUT45), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n745), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1076), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(G8), .A3(G168), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1072), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1061), .A2(new_n1071), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1016), .B(G8), .C1(new_n1067), .C2(new_n1033), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1066), .A2(new_n1070), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1087), .B1(new_n1089), .B2(new_n1084), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1057), .B(KEYINPUT113), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1059), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(new_n1063), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1060), .A2(new_n1088), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g673(.A(KEYINPUT114), .B1(new_n1060), .B2(new_n1088), .C1(new_n1063), .C2(new_n1095), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1091), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1089), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1066), .A2(new_n1070), .A3(KEYINPUT124), .A4(new_n1088), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  OR4_X1    g680(.A1(new_n1105), .A2(new_n1080), .A3(new_n1081), .A4(G2078), .ZN(new_n1106));
  INV_X1    g681(.A(G1961), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1105), .B1(new_n1025), .B2(G2078), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OR3_X1    g685(.A1(new_n530), .A2(KEYINPUT54), .A3(new_n532), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n530), .B2(new_n532), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1109), .A2(new_n1108), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1022), .B1(new_n886), .B2(G1384), .ZN(new_n1115));
  AND4_X1   g690(.A1(KEYINPUT53), .A2(new_n1024), .A3(new_n773), .A4(new_n1028), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1110), .A2(new_n1113), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1103), .A2(new_n1104), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1083), .A2(G8), .ZN(new_n1121));
  NOR2_X1   g696(.A1(G168), .A2(new_n1038), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(KEYINPUT51), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(G8), .C1(new_n1083), .C2(G286), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1083), .A2(KEYINPUT122), .A3(new_n1122), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT122), .B1(new_n1083), .B2(new_n1122), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1120), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1083), .A2(new_n1122), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1083), .A2(KEYINPUT122), .A3(new_n1122), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(KEYINPUT123), .A3(new_n1126), .A4(new_n1124), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1119), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1996), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1023), .A2(new_n1024), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1029), .A2(new_n1028), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT59), .B1(new_n1144), .B2(new_n541), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1146), .B(new_n853), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n561), .A2(new_n937), .A3(new_n939), .A4(KEYINPUT57), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n943), .B2(new_n938), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT56), .B(G2072), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1023), .A2(new_n1024), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n822), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1152), .B1(new_n1155), .B2(new_n1154), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1156), .B(new_n1157), .C1(new_n1158), .C2(KEYINPUT61), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1152), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT61), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1148), .A2(new_n1159), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n832), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1141), .A2(G2067), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT118), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT118), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  OAI211_X1 g744(.A(KEYINPUT121), .B(KEYINPUT60), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n607), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT118), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT118), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT121), .B1(new_n1176), .B2(KEYINPUT60), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT60), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n1180), .A3(new_n935), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1168), .A2(new_n1169), .A3(KEYINPUT60), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1165), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1176), .A2(new_n935), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1160), .A2(KEYINPUT119), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1152), .B1(new_n1160), .B2(KEYINPUT119), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1185), .A2(new_n1156), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1101), .B1(new_n1138), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1131), .A2(new_n1191), .A3(new_n1137), .ZN(new_n1192));
  AND4_X1   g767(.A1(G171), .A2(new_n1103), .A3(new_n1104), .A4(new_n1110), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1192), .B(new_n1193), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g771(.A(KEYINPUT125), .B(new_n1191), .C1(new_n1131), .C2(new_n1137), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1190), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1115), .A2(new_n1019), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1199), .A2(new_n738), .A3(new_n735), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1199), .A2(G1986), .A3(G290), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT111), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n767), .B(G2067), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n788), .A2(G1996), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n787), .A2(new_n1139), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  XOR2_X1   g782(.A(new_n730), .B(new_n733), .Z(new_n1208));
  OR2_X1    g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1203), .B1(new_n1199), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1198), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1199), .A2(new_n1139), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT46), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n788), .A2(new_n1204), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1212), .A2(new_n1213), .B1(new_n1199), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(new_n1213), .B2(new_n1212), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1216), .B(KEYINPUT47), .Z(new_n1217));
  NAND2_X1  g792(.A1(new_n731), .A2(new_n733), .ZN(new_n1218));
  OAI22_X1  g793(.A1(new_n1207), .A2(new_n1218), .B1(G2067), .B2(new_n887), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(new_n1199), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1200), .B(KEYINPUT48), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1209), .A2(new_n1199), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1221), .B1(new_n1222), .B2(KEYINPUT126), .ZN(new_n1223));
  AND2_X1   g798(.A1(new_n1222), .A2(KEYINPUT126), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1220), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1217), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1211), .A2(new_n1226), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g802(.A1(G227), .A2(new_n459), .ZN(new_n1229));
  XNOR2_X1  g803(.A(new_n1229), .B(KEYINPUT127), .ZN(new_n1230));
  AOI21_X1  g804(.A(new_n1230), .B1(new_n692), .B2(new_n697), .ZN(new_n1231));
  OAI21_X1  g805(.A(new_n1231), .B1(new_n653), .B2(new_n654), .ZN(new_n1232));
  AOI21_X1  g806(.A(new_n1232), .B1(new_n910), .B2(new_n915), .ZN(new_n1233));
  AND3_X1   g807(.A1(new_n1233), .A2(new_n999), .A3(new_n1002), .ZN(G308));
  NAND3_X1  g808(.A1(new_n1233), .A2(new_n999), .A3(new_n1002), .ZN(G225));
endmodule


