//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n452), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n463), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n486), .B1(new_n468), .B2(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n486), .B(new_n489), .C1(new_n469), .C2(new_n468), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n463), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n479), .A2(G126), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n491), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n491), .B2(new_n496), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT72), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT71), .A2(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(KEYINPUT6), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n505), .B2(new_n507), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n509), .A2(new_n514), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n508), .A2(G51), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n500), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n524), .A2(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n521), .A2(new_n522), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(G64), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(G52), .A2(new_n508), .B1(new_n513), .B2(G90), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n538), .B1(new_n535), .B2(new_n536), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT73), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n508), .A2(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n513), .A2(G81), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT75), .B1(new_n510), .B2(new_n511), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n527), .A2(new_n558), .A3(new_n528), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n556), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n513), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT74), .A2(G53), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n565), .B1(new_n508), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT71), .B1(KEYINPUT72), .B2(G651), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n507), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND4_X1   g145(.A1(new_n565), .A2(new_n570), .A3(G543), .A4(new_n566), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n563), .B(new_n564), .C1(new_n567), .C2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n570), .A2(G91), .A3(new_n529), .ZN(new_n575));
  NOR3_X1   g150(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT75), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n558), .B1(new_n527), .B2(new_n528), .ZN(new_n577));
  OAI21_X1  g152(.A(G65), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(new_n561), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n575), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n508), .A2(new_n565), .A3(new_n566), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n570), .A2(G543), .A3(new_n566), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n580), .A2(KEYINPUT76), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n574), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  NAND3_X1  g162(.A1(new_n570), .A2(G87), .A3(new_n529), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n570), .A2(G49), .A3(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n570), .A2(new_n529), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT77), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n513), .A2(new_n595), .A3(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n512), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n508), .A2(G48), .B1(new_n600), .B2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n538), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT79), .B(G85), .Z(new_n607));
  NAND2_X1  g182(.A1(new_n513), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n508), .ZN(new_n609));
  INV_X1    g184(.A(G47), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n608), .B(new_n613), .C1(new_n609), .C2(new_n610), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n606), .A2(new_n612), .A3(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n557), .A2(new_n559), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(new_n538), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n508), .A2(G54), .ZN(new_n620));
  AOI21_X1  g195(.A(KEYINPUT10), .B1(new_n513), .B2(G92), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n513), .A2(KEYINPUT10), .A3(G92), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n616), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NOR2_X1   g202(.A1(G286), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n586), .B2(new_n627), .ZN(G297));
  AOI21_X1  g204(.A(new_n628), .B1(new_n586), .B2(new_n627), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n624), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g211(.A(new_n472), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n464), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n477), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n479), .A2(G123), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n646), .A2(KEYINPUT81), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(KEYINPUT81), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(G111), .B2(new_n463), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n644), .B(new_n645), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n642), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT82), .ZN(G156));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(G1341), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G1348), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n669), .B1(new_n668), .B2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n658), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n675), .A2(new_n657), .A3(new_n671), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n674), .A2(new_n676), .A3(G14), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G401));
  XOR2_X1   g253(.A(G2067), .B(G2678), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n682), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n681), .B1(new_n687), .B2(KEYINPUT17), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n685), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G2096), .B(G2100), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1956), .B(G2474), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1961), .B(G1966), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n701), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(KEYINPUT20), .ZN(new_n707));
  OAI221_X1 g282(.A(new_n702), .B1(new_n699), .B2(new_n703), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1991), .B(G1996), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n710), .A2(new_n712), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n696), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n715), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n717), .A2(new_n695), .A3(new_n713), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n716), .A2(new_n718), .ZN(G229));
  INV_X1    g294(.A(KEYINPUT100), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G5), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G301), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(G16), .A2(G19), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n549), .B2(new_n721), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n725), .A2(G1961), .B1(new_n667), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2090), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n483), .A2(G29), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G35), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n730), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n729), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(new_n463), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n477), .A2(G139), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n740), .A2(new_n743), .A3(G29), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G33), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT91), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(G160), .A2(G29), .ZN(new_n751));
  AND2_X1   g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  NOR2_X1   g327(.A1(KEYINPUT24), .A2(G34), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n731), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n745), .A2(G2072), .A3(new_n747), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n751), .A2(G2084), .A3(new_n755), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n750), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n728), .A2(new_n738), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n721), .A2(G4), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n623), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT99), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n735), .A2(new_n729), .A3(new_n737), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n764), .A2(new_n669), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n764), .A2(new_n669), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n731), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n731), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(G2078), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n727), .A2(new_n667), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(G2078), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n731), .A2(G32), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT94), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT26), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n479), .A2(G129), .B1(G105), .B2(new_n637), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n477), .A2(G141), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n778), .B(new_n779), .C1(new_n786), .C2(new_n731), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n731), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT90), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n477), .A2(G140), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n479), .A2(G128), .ZN(new_n792));
  OR2_X1    g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G29), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n790), .A2(new_n796), .A3(G2067), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n778), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n731), .B1(new_n782), .B2(new_n785), .ZN(new_n803));
  INV_X1    g378(.A(new_n779), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n787), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n766), .A2(new_n765), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n762), .A2(new_n769), .A3(new_n776), .A4(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n650), .A2(new_n810), .A3(new_n731), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n650), .B2(new_n731), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT31), .B(G11), .Z(new_n813));
  INV_X1    g388(.A(G28), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(KEYINPUT30), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT97), .Z(new_n816));
  AOI21_X1  g391(.A(G29), .B1(new_n814), .B2(KEYINPUT30), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n811), .A2(new_n812), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n725), .B2(G1961), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n721), .A2(G21), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G286), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1966), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(KEYINPUT98), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n825));
  INV_X1    g400(.A(new_n819), .ZN(new_n826));
  INV_X1    g401(.A(G1961), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n724), .ZN(new_n828));
  INV_X1    g403(.A(G1966), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n822), .B(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n825), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n574), .A2(G16), .A3(new_n585), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n721), .A2(G20), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT23), .ZN(new_n835));
  AOI21_X1  g410(.A(G1956), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n833), .A2(G1956), .A3(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n720), .B1(new_n809), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n761), .A2(new_n738), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n727), .A2(new_n667), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n827), .B2(new_n724), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n842), .A2(new_n844), .A3(new_n807), .A4(new_n806), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(new_n775), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n824), .A2(new_n831), .B1(new_n838), .B2(new_n837), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT100), .A4(new_n769), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n721), .A2(G22), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G303), .B2(G16), .ZN(new_n851));
  INV_X1    g426(.A(G1971), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n721), .A2(G6), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G305), .B2(G16), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT32), .B(G1981), .Z(new_n856));
  AND2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G23), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(G16), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(G288), .B2(G16), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT87), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT33), .B(G1976), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT34), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT34), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n859), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT88), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n731), .A2(G25), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n477), .A2(G131), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n479), .A2(G119), .ZN(new_n876));
  OR2_X1    g451(.A1(G95), .A2(G2105), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n874), .B1(new_n880), .B2(new_n731), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G1991), .Z(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n881), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(G290), .A2(G16), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n721), .A2(G24), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G1986), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(G1986), .A3(new_n886), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n872), .A2(new_n873), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n873), .B1(new_n872), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n870), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT36), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(KEYINPUT89), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI221_X1 g472(.A(new_n870), .B1(KEYINPUT89), .B2(new_n895), .C1(new_n892), .C2(new_n893), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n849), .B1(new_n897), .B2(new_n898), .ZN(G311));
  NOR2_X1   g474(.A1(G311), .A2(KEYINPUT101), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n901));
  AOI211_X1 g476(.A(new_n901), .B(new_n849), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(G150));
  NAND2_X1  g478(.A1(new_n624), .A2(G559), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n508), .A2(G55), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n513), .A2(G93), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n906), .B(new_n907), .C1(new_n538), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n549), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n905), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n912));
  AOI21_X1  g487(.A(G860), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n912), .B2(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(G860), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT37), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(G145));
  NAND2_X1  g492(.A1(new_n479), .A2(G130), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n463), .A2(G118), .ZN(new_n919));
  OAI21_X1  g494(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(G142), .B2(new_n477), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(new_n639), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(new_n880), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n740), .A2(new_n744), .A3(new_n743), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT102), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(new_n786), .ZN(new_n927));
  INV_X1    g502(.A(new_n795), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n491), .A2(new_n496), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n929), .A2(new_n491), .A3(new_n496), .A4(new_n930), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n924), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(G160), .B(new_n650), .Z(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(new_n483), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT103), .A4(new_n924), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n933), .A2(new_n934), .ZN(new_n941));
  INV_X1    g516(.A(new_n924), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n937), .B1(new_n945), .B2(new_n935), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(G395));
  XOR2_X1   g525(.A(G290), .B(G305), .Z(new_n951));
  XNOR2_X1  g526(.A(G303), .B(G288), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT42), .Z(new_n954));
  XNOR2_X1  g529(.A(new_n633), .B(new_n910), .ZN(new_n955));
  NAND2_X1  g530(.A1(G299), .A2(new_n624), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n586), .A2(new_n623), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(KEYINPUT41), .A3(new_n957), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n955), .B2(new_n958), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n954), .A2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n909), .A2(new_n627), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  NAND2_X1  g544(.A1(new_n960), .A2(new_n961), .ZN(new_n970));
  XNOR2_X1  g545(.A(G301), .B(G286), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(new_n910), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n971), .A2(KEYINPUT105), .A3(new_n910), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT105), .B1(new_n971), .B2(new_n910), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n910), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n956), .B2(new_n957), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n970), .A2(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n953), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n974), .A2(new_n975), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n982), .A2(new_n978), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n960), .A2(new_n961), .B1(new_n973), .B2(new_n977), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n953), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n981), .A2(KEYINPUT43), .A3(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n979), .A2(new_n980), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT43), .B1(new_n987), .B2(new_n981), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT44), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n981), .A2(new_n990), .A3(new_n985), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n987), .B2(new_n981), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n993), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g569(.A(KEYINPUT106), .B(G1384), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n491), .B2(new_n496), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  INV_X1    g573(.A(G40), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n467), .A2(new_n999), .A3(new_n473), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT107), .Z(new_n1002));
  XNOR2_X1  g577(.A(new_n795), .B(new_n798), .ZN(new_n1003));
  INV_X1    g578(.A(G1996), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(new_n786), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1001), .A2(G1996), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1002), .A2(new_n1005), .B1(new_n786), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1002), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n879), .B(new_n882), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(G290), .A2(G1986), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1001), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT108), .Z(new_n1015));
  INV_X1    g590(.A(KEYINPUT61), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n1017), .B(KEYINPUT57), .C1(new_n572), .C2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n572), .B2(new_n1018), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n572), .B2(new_n1017), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1019), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n465), .A2(new_n466), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G2105), .ZN(new_n1026));
  INV_X1    g601(.A(new_n473), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(G40), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(KEYINPUT45), .B2(new_n996), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT56), .B(G2072), .ZN(new_n1030));
  INV_X1    g605(.A(new_n490), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n489), .B1(new_n464), .B2(new_n486), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n479), .A2(G126), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n493), .A2(new_n495), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT70), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n491), .A2(new_n492), .A3(new_n496), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1029), .B(new_n1030), .C1(new_n1039), .C2(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT121), .ZN(new_n1041));
  INV_X1    g616(.A(G1384), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n497), .B2(new_n498), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n998), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT118), .B(G1956), .ZN(new_n1048));
  NOR2_X1   g623(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1053));
  OAI21_X1  g628(.A(new_n1000), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1024), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n582), .B(new_n565), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n563), .A2(new_n564), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1018), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(KEYINPUT120), .A3(new_n1022), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n572), .A2(new_n1017), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT57), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1060), .B(new_n1055), .C1(new_n1062), .C2(new_n1020), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1016), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT119), .B1(new_n580), .B2(new_n584), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT57), .B(new_n1061), .C1(new_n1066), .C2(new_n1017), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1067), .A2(new_n1055), .A3(new_n1060), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1047), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n932), .A2(new_n1042), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1053), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1028), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1049), .B1(new_n497), .B2(new_n498), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1041), .A2(new_n1046), .B1(new_n1074), .B2(new_n1048), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1069), .B(KEYINPUT61), .C1(new_n1024), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1000), .A2(new_n1052), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G2067), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1000), .B(new_n1079), .C1(new_n1039), .C2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1081), .B2(new_n669), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n669), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1078), .ZN(new_n1085));
  AND4_X1   g660(.A1(KEYINPUT60), .A2(new_n1084), .A3(new_n623), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n623), .B1(new_n1082), .B2(KEYINPUT60), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1044), .A2(new_n1004), .A3(new_n1029), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1077), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n549), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1065), .A2(new_n1076), .A3(new_n1088), .A4(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1082), .A2(new_n623), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1069), .B1(new_n1056), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT122), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n1069), .C1(new_n1056), .C2(new_n1096), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1102));
  AND3_X1   g677(.A1(G303), .A2(G8), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(G303), .B2(G8), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT115), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1072), .A2(new_n1073), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1109), .A3(new_n729), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1029), .B1(new_n1039), .B2(KEYINPUT45), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n852), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1106), .B1(new_n1113), .B2(G8), .ZN(new_n1114));
  INV_X1    g689(.A(G8), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1116), .A2(new_n729), .A3(new_n1000), .A4(new_n1079), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n1115), .B(new_n1105), .C1(new_n1112), .C2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1115), .B1(new_n1000), .B2(new_n1052), .ZN(new_n1120));
  INV_X1    g695(.A(G1981), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n513), .A2(G86), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n601), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n595), .B1(new_n513), .B2(G86), .ZN(new_n1124));
  AND4_X1   g699(.A1(new_n595), .A2(new_n570), .A3(G86), .A4(new_n529), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n601), .B(new_n1121), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT113), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT113), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n597), .A2(new_n1128), .A3(new_n1121), .A4(new_n601), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1123), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1120), .B1(new_n1130), .B2(KEYINPUT49), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT49), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1132), .B(new_n1123), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT111), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n589), .A2(new_n590), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1138), .A2(KEYINPUT111), .A3(G1976), .A4(new_n588), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1120), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT52), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1120), .A2(new_n1137), .A3(new_n1142), .A4(new_n1139), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT112), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1141), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1134), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1043), .A2(KEYINPUT50), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1028), .A2(G2084), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT45), .B(new_n1042), .C1(new_n497), .C2(new_n498), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1028), .B1(new_n1070), .B2(new_n998), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1150), .A2(new_n1151), .B1(new_n1154), .B2(new_n829), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1115), .B1(new_n1155), .B2(G168), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n829), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1079), .B(new_n1151), .C1(new_n1039), .C2(new_n1080), .ZN(new_n1158));
  AOI21_X1  g733(.A(G168), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1149), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(G168), .A3(new_n1158), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(G8), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1163), .A2(KEYINPUT51), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1119), .B(new_n1148), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G2078), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1029), .B(new_n1166), .C1(new_n1039), .C2(KEYINPUT45), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT53), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1081), .A2(new_n827), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n997), .A2(new_n998), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n996), .A2(KEYINPUT45), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1166), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1173), .B(new_n467), .C1(new_n1174), .C2(new_n473), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1027), .A2(KEYINPUT123), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1169), .A2(new_n1170), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(G171), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1168), .A2(new_n1167), .B1(new_n1081), .B2(new_n827), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1152), .A2(new_n1153), .A3(KEYINPUT53), .A4(new_n1166), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1179), .B(KEYINPUT54), .C1(G171), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n1184));
  AOI21_X1  g759(.A(G301), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1185));
  AND4_X1   g760(.A1(G301), .A2(new_n1169), .A3(new_n1170), .A4(new_n1177), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1165), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1101), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1115), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1191), .A2(KEYINPUT116), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(KEYINPUT116), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1192), .A2(new_n1105), .A3(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1143), .B(new_n1144), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1195), .B(new_n1141), .C1(new_n1133), .C2(new_n1131), .ZN(new_n1196));
  NAND2_X1  g771(.A1(G168), .A2(G8), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1155), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT63), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1202), .A2(G8), .A3(new_n1106), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1155), .A2(KEYINPUT63), .A3(new_n1197), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1203), .B1(new_n1205), .B2(new_n1114), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1138), .A2(new_n1136), .A3(new_n588), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1207), .B1(new_n1134), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1120), .B(KEYINPUT114), .Z(new_n1210));
  AOI22_X1  g785(.A1(new_n1206), .A2(new_n1148), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT117), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1201), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1214));
  AOI21_X1  g789(.A(G2090), .B1(new_n1074), .B2(KEYINPUT115), .ZN(new_n1215));
  AOI22_X1  g790(.A1(new_n1215), .A2(new_n1109), .B1(new_n852), .B2(new_n1111), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1105), .B1(new_n1216), .B2(new_n1115), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1118), .B1(new_n1217), .B2(new_n1204), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1214), .B1(new_n1218), .B2(new_n1196), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT63), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1220), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1221));
  OAI21_X1  g796(.A(KEYINPUT117), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1190), .A2(new_n1213), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n1225));
  OAI21_X1  g800(.A(KEYINPUT51), .B1(new_n1163), .B2(new_n1159), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1156), .A2(new_n1149), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1148), .A2(new_n1217), .A3(new_n1185), .A4(new_n1203), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1226), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1224), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1115), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1203), .B1(new_n1233), .B2(new_n1106), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1182), .A2(G171), .ZN(new_n1235));
  NOR3_X1   g810(.A1(new_n1234), .A2(new_n1235), .A3(new_n1196), .ZN(new_n1236));
  OAI21_X1  g811(.A(KEYINPUT62), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1237));
  AND4_X1   g812(.A1(new_n1224), .A2(new_n1236), .A3(new_n1237), .A4(new_n1231), .ZN(new_n1238));
  NOR2_X1   g813(.A1(new_n1232), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g814(.A(new_n1015), .B1(new_n1223), .B2(new_n1239), .ZN(new_n1240));
  XOR2_X1   g815(.A(new_n1006), .B(KEYINPUT46), .Z(new_n1241));
  NAND2_X1  g816(.A1(new_n1003), .A2(new_n786), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g819(.A(new_n1244), .B(KEYINPUT47), .ZN(new_n1245));
  NOR2_X1   g820(.A1(new_n1011), .A2(new_n1001), .ZN(new_n1246));
  XNOR2_X1  g821(.A(new_n1246), .B(KEYINPUT48), .ZN(new_n1247));
  OAI21_X1  g822(.A(new_n1245), .B1(new_n1010), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g823(.A1(new_n879), .A2(new_n883), .ZN(new_n1249));
  XNOR2_X1  g824(.A(new_n1249), .B(KEYINPUT125), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1007), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n928), .A2(new_n798), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1008), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g828(.A(KEYINPUT126), .ZN(new_n1254));
  AND2_X1   g829(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g830(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1256));
  NOR3_X1   g831(.A1(new_n1248), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1240), .A2(new_n1257), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g833(.A1(G227), .A2(new_n461), .ZN(new_n1260));
  AOI21_X1  g834(.A(new_n1260), .B1(new_n716), .B2(new_n718), .ZN(new_n1261));
  AND3_X1   g835(.A1(new_n1261), .A2(new_n677), .A3(KEYINPUT127), .ZN(new_n1262));
  AOI21_X1  g836(.A(KEYINPUT127), .B1(new_n1261), .B2(new_n677), .ZN(new_n1263));
  OAI21_X1  g837(.A(new_n948), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g838(.A1(new_n1264), .A2(new_n993), .ZN(G308));
  OAI221_X1 g839(.A(new_n948), .B1(new_n1262), .B2(new_n1263), .C1(new_n991), .C2(new_n992), .ZN(G225));
endmodule


