//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n203), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  INV_X1    g0011(.A(KEYINPUT1), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n212), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n203), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n217), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AND3_X1   g0023(.A1(new_n213), .A2(new_n214), .A3(new_n223), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G58), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(KEYINPUT68), .ZN(new_n241));
  AND2_X1   g0041(.A1(KEYINPUT3), .A2(G33), .ZN(new_n242));
  NOR2_X1   g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n246), .A2(G223), .B1(G77), .B2(new_n244), .ZN(new_n247));
  INV_X1    g0047(.A(G222), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G1698), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n249), .B(new_n251), .C1(new_n242), .C2(new_n243), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n247), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n254), .A2(new_n260), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(G226), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G169), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n241), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G179), .ZN(new_n267));
  INV_X1    g0067(.A(new_n264), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(KEYINPUT68), .A3(new_n267), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n218), .B1(new_n203), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n219), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G58), .A2(G68), .ZN(new_n279));
  INV_X1    g0079(.A(G50), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n219), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n272), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G13), .A3(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT66), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT66), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n286), .A2(new_n283), .A3(G13), .A4(G20), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n272), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n219), .A2(G1), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n289), .A2(KEYINPUT67), .A3(new_n280), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT67), .B1(new_n289), .B2(new_n280), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n285), .A2(new_n287), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n282), .B(new_n292), .C1(G50), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n270), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n269), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n262), .A2(G244), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n246), .A2(G238), .B1(G107), .B2(new_n244), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n226), .B2(new_n252), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n261), .B(new_n297), .C1(new_n299), .C2(new_n254), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(new_n267), .ZN(new_n301));
  INV_X1    g0101(.A(new_n273), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n303));
  XOR2_X1   g0103(.A(KEYINPUT15), .B(G87), .Z(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n274), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G77), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n285), .A2(new_n287), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n306), .A2(new_n272), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n289), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n288), .A2(G77), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n300), .B2(G169), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n301), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n300), .B2(G190), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n300), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n264), .A2(KEYINPUT69), .A3(G200), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n264), .A2(G200), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n268), .A2(G190), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n294), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n294), .A2(new_n328), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT70), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n331), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n333), .A2(new_n322), .A3(new_n334), .A4(new_n325), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n323), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT10), .ZN(new_n338));
  AOI211_X1 g0138(.A(new_n296), .B(new_n319), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n273), .A2(new_n289), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n308), .A2(new_n273), .B1(new_n288), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n343));
  INV_X1    g0143(.A(G68), .ZN(new_n344));
  NAND2_X1  g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n271), .A2(KEYINPUT76), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT76), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n346), .B1(new_n350), .B2(KEYINPUT3), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n271), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(new_n219), .A3(new_n345), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n344), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G58), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n344), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n279), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n276), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n343), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT79), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n343), .C1(new_n357), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT76), .B(G33), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n219), .B(new_n353), .C1(new_n368), .C2(new_n352), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n355), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n355), .A2(G20), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n353), .B(new_n371), .C1(new_n368), .C2(new_n352), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT77), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n350), .A2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n353), .A4(new_n371), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G68), .ZN(new_n378));
  INV_X1    g0178(.A(new_n362), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n367), .A2(new_n380), .A3(new_n272), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n272), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n362), .B1(new_n377), .B2(G68), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(KEYINPUT16), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT80), .A3(new_n367), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n342), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n261), .B1(G232), .B2(new_n262), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT65), .B(G1698), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G223), .ZN(new_n391));
  INV_X1    g0191(.A(G226), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n245), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n353), .B1(new_n368), .B2(new_n352), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(G33), .B2(G87), .ZN(new_n395));
  INV_X1    g0195(.A(new_n254), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n389), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G169), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n267), .B2(new_n397), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n388), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n386), .A2(KEYINPUT80), .A3(new_n367), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT80), .B1(new_n386), .B2(new_n367), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n341), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n399), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n397), .A2(new_n317), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(G190), .B2(new_n397), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n341), .B(new_n408), .C1(new_n402), .C2(new_n403), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n388), .A2(KEYINPUT17), .A3(new_n408), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n401), .A2(new_n406), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n261), .B1(G238), .B2(new_n262), .ZN(new_n415));
  OAI211_X1 g0215(.A(G232), .B(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT71), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n353), .A2(new_n345), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT71), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(G232), .A4(G1698), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n390), .A3(G226), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n417), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT72), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(new_n254), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(new_n423), .B2(new_n254), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n415), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n415), .C1(new_n425), .C2(new_n426), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G200), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n308), .A2(new_n344), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT12), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n277), .A2(new_n280), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n274), .A2(new_n307), .B1(new_n219), .B2(G68), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n272), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT11), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n288), .A2(G68), .A3(new_n310), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT73), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n428), .A2(G190), .A3(new_n430), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n432), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT14), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n423), .A2(new_n254), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT72), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n423), .A2(new_n424), .A3(new_n254), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n429), .B1(new_n449), .B2(new_n415), .ZN(new_n450));
  INV_X1    g0250(.A(new_n430), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n445), .B(G169), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(G169), .B1(new_n450), .B2(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT14), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n431), .A2(KEYINPUT74), .A3(new_n445), .A4(G169), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n428), .A2(G179), .A3(new_n430), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n454), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n441), .B(KEYINPUT75), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n444), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n339), .A2(new_n414), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G87), .ZN(new_n463));
  OR4_X1    g0263(.A1(KEYINPUT22), .A2(new_n244), .A3(G20), .A4(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n352), .B1(new_n347), .B2(new_n349), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n219), .B(G87), .C1(new_n465), .C2(new_n243), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT88), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT22), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n466), .B2(KEYINPUT22), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT24), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n350), .A2(G116), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G20), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n219), .B2(G107), .ZN(new_n475));
  INV_X1    g0275(.A(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(KEYINPUT23), .A3(G20), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n470), .A2(new_n471), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n471), .B1(new_n470), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n272), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n283), .A2(G33), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n288), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n308), .A2(KEYINPUT25), .A3(new_n476), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT25), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n293), .B2(G107), .ZN(new_n486));
  AOI22_X1  g0286(.A1(G107), .A2(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n259), .A2(G1), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT5), .B(G41), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n254), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G264), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n489), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n257), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n249), .A2(new_n251), .A3(G250), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G257), .A2(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n394), .A2(new_n498), .B1(G294), .B2(new_n350), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n492), .B(new_n495), .C1(new_n499), .C2(new_n396), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n265), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(G179), .B2(new_n500), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n488), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT89), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n488), .A2(KEYINPUT89), .A3(new_n503), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n488), .ZN(new_n509));
  INV_X1    g0309(.A(G190), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(G200), .B2(new_n500), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n491), .A2(G257), .B1(new_n494), .B2(new_n257), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  OAI211_X1 g0316(.A(G250), .B(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n517));
  NAND2_X1  g0317(.A1(KEYINPUT4), .A2(G244), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n516), .B(new_n517), .C1(new_n252), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(new_n390), .C1(new_n465), .C2(new_n243), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(G190), .B(new_n515), .C1(new_n522), .C2(new_n396), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n520), .ZN(new_n525));
  INV_X1    g0325(.A(new_n519), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n254), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(G190), .A4(new_n515), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n476), .B1(new_n351), .B2(new_n356), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(KEYINPUT6), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(KEYINPUT81), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  AND2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n534), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(KEYINPUT6), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(G97), .A4(new_n476), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n219), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n277), .A2(new_n307), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n532), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT82), .B1(new_n545), .B2(new_n384), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n539), .A2(new_n542), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n547), .B2(G20), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT7), .B1(new_n244), .B2(new_n219), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n368), .B2(new_n352), .ZN(new_n551));
  OAI21_X1  g0351(.A(G107), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT82), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n272), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT83), .ZN(new_n556));
  INV_X1    g0356(.A(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n293), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n556), .B(new_n558), .C1(new_n483), .C2(new_n557), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n288), .B2(new_n482), .ZN(new_n560));
  INV_X1    g0360(.A(new_n558), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT83), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n546), .A2(new_n555), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n515), .B1(new_n522), .B2(new_n396), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n531), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n489), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n567), .A2(G250), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n396), .A2(new_n568), .B1(new_n257), .B2(new_n489), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(G1698), .C1(new_n465), .C2(new_n243), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT85), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT85), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n394), .A2(new_n573), .A3(G244), .A4(G1698), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n394), .A2(G238), .A3(new_n390), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n472), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n570), .B1(new_n576), .B2(new_n254), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n267), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n219), .B(G68), .C1(new_n465), .C2(new_n243), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n219), .B1(new_n422), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT86), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n537), .A2(new_n463), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(new_n219), .C1(new_n422), .C2(new_n580), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n580), .B1(new_n274), .B2(new_n557), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n272), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n483), .A2(new_n304), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n308), .A2(new_n305), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n578), .B(new_n592), .C1(G169), .C2(new_n577), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n576), .A2(new_n254), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n569), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n483), .A2(G87), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n589), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n577), .B2(G190), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n559), .A2(new_n562), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n554), .B1(new_n553), .B2(new_n272), .ZN(new_n602));
  AOI211_X1 g0402(.A(KEYINPUT82), .B(new_n384), .C1(new_n548), .C2(new_n552), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n564), .A2(new_n265), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n396), .B1(new_n525), .B2(new_n526), .ZN(new_n606));
  INV_X1    g0406(.A(new_n515), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n267), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n566), .A2(new_n593), .A3(new_n600), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n394), .A2(G264), .A3(G1698), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n394), .A2(G257), .A3(new_n390), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n244), .A2(G303), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n254), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n493), .A2(new_n396), .A3(G270), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n495), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n293), .A2(G116), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT87), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n516), .B(new_n219), .C1(G33), .C2(new_n557), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n272), .C1(new_n219), .C2(G116), .ZN(new_n626));
  XOR2_X1   g0426(.A(new_n626), .B(KEYINPUT20), .Z(new_n627));
  NAND2_X1  g0427(.A1(new_n483), .A2(G116), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n621), .B(new_n630), .C1(new_n510), .C2(new_n620), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n620), .A3(G169), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT21), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n267), .B(new_n618), .C1(new_n615), .C2(new_n254), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n629), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n629), .A2(new_n620), .A3(KEYINPUT21), .A4(G169), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n631), .A2(new_n634), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NOR4_X1   g0438(.A1(new_n462), .A2(new_n514), .A3(new_n611), .A4(new_n638), .ZN(G372));
  NAND2_X1  g0439(.A1(new_n336), .A2(new_n338), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n459), .A2(new_n460), .B1(new_n443), .B2(new_n314), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n411), .A2(new_n412), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n401), .A2(new_n406), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n296), .ZN(new_n646));
  INV_X1    g0446(.A(new_n592), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n595), .B2(new_n265), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n578), .B1(new_n596), .B2(new_n599), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n610), .A2(KEYINPUT91), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT91), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n604), .A2(new_n652), .A3(new_n605), .A4(new_n609), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n594), .A2(G190), .A3(new_n569), .ZN(new_n655));
  INV_X1    g0455(.A(new_n598), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n577), .A2(new_n317), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n592), .B1(new_n577), .B2(G169), .ZN(new_n659));
  AOI211_X1 g0459(.A(G179), .B(new_n570), .C1(new_n576), .C2(new_n254), .ZN(new_n660));
  OAI22_X1  g0460(.A1(new_n657), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n661), .B2(new_n610), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n654), .A2(new_n662), .A3(new_n593), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT92), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n654), .A2(new_n662), .A3(KEYINPUT92), .A4(new_n593), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n611), .B1(new_n509), .B2(new_n512), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT90), .B1(new_n488), .B2(new_n503), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  AOI211_X1 g0470(.A(new_n670), .B(new_n502), .C1(new_n481), .C2(new_n487), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n645), .B(new_n646), .C1(new_n462), .C2(new_n673), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n283), .A2(new_n219), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n668), .A2(new_n630), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n630), .A2(new_n681), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n638), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n514), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n509), .B2(new_n681), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n488), .A2(new_n503), .A3(new_n680), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n668), .A2(new_n680), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n669), .A2(new_n671), .A3(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n689), .A2(new_n693), .ZN(G399));
  NOR2_X1   g0494(.A1(new_n583), .A2(G116), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n215), .A2(new_n258), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n221), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n673), .A2(new_n680), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n506), .A2(new_n507), .A3(new_n668), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n667), .ZN(new_n702));
  INV_X1    g0502(.A(new_n610), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n649), .A2(new_n651), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n593), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(KEYINPUT26), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n680), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  MUX2_X1   g0509(.A(new_n700), .B(new_n709), .S(KEYINPUT29), .Z(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n680), .A2(KEYINPUT31), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n492), .B1(new_n499), .B2(new_n396), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n564), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n635), .A3(new_n577), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n714), .A2(new_n635), .A3(KEYINPUT30), .A4(new_n577), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT93), .ZN(new_n720));
  INV_X1    g0520(.A(new_n500), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n608), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n500), .B(KEYINPUT93), .C1(new_n606), .C2(new_n607), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n620), .A2(new_n267), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n577), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n712), .B1(new_n719), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  INV_X1    g0529(.A(new_n723), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT93), .B1(new_n564), .B2(new_n500), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n595), .A2(new_n267), .A3(new_n620), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n724), .A2(new_n726), .A3(KEYINPUT94), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n717), .A4(new_n718), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n680), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n728), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n611), .A2(new_n638), .A3(new_n680), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(new_n506), .A3(new_n507), .A4(new_n513), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n711), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n710), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n699), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(new_n685), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n219), .A2(G13), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n283), .B1(new_n746), .B2(G45), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n696), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G330), .B2(new_n684), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n418), .A2(new_n215), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n215), .ZN(new_n754));
  INV_X1    g0554(.A(new_n394), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n215), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n259), .B2(new_n222), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n236), .A2(new_n259), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n218), .B1(G20), .B2(new_n265), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n749), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n219), .A2(new_n267), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n510), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n280), .A2(new_n770), .B1(new_n772), .B2(new_n344), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n510), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n219), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n557), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n767), .A2(G190), .A3(new_n317), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n418), .B1(new_n777), .B2(new_n358), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n773), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n219), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n463), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT32), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G159), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n782), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n787), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n780), .A2(new_n510), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n789), .A2(KEYINPUT32), .B1(G107), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n767), .A2(new_n784), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G77), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n779), .A2(new_n788), .A3(new_n792), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G317), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n772), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n801), .B(new_n805), .C1(G326), .C2(new_n769), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n785), .B(KEYINPUT97), .Z(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n777), .A2(new_n809), .B1(new_n793), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n775), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(G294), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n806), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n244), .B1(new_n781), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT96), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n799), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n766), .B1(new_n818), .B2(new_n763), .ZN(new_n819));
  INV_X1    g0619(.A(new_n762), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n684), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n751), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  INV_X1    g0623(.A(new_n319), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n665), .A2(new_n666), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n672), .A2(new_n667), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n824), .B(new_n681), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n312), .A2(new_n680), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n318), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n315), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n314), .A2(new_n681), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n827), .B1(new_n700), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n742), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n749), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n763), .A2(new_n760), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n748), .B1(new_n307), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n763), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n770), .A2(new_n815), .B1(new_n790), .B2(new_n463), .ZN(new_n842));
  INV_X1    g0642(.A(new_n781), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(G107), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n777), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n418), .B(new_n776), .C1(G294), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n807), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(new_n846), .C1(new_n810), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT98), .ZN(new_n849));
  INV_X1    g0649(.A(G116), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n796), .A2(new_n850), .B1(new_n800), .B2(new_n772), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n849), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G137), .A2(new_n769), .B1(new_n845), .B2(G143), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n854), .B1(new_n275), .B2(new_n772), .C1(new_n796), .C2(new_n786), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n775), .A2(new_n358), .B1(new_n790), .B2(new_n344), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n394), .B1(new_n280), .B2(new_n781), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n807), .C2(G132), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n852), .A2(new_n853), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n840), .B1(new_n841), .B2(new_n860), .C1(new_n834), .C2(new_n761), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n838), .A2(new_n861), .ZN(G384));
  OAI211_X1 g0662(.A(G116), .B(new_n220), .C1(new_n547), .C2(KEYINPUT35), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(KEYINPUT99), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(KEYINPUT99), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT36), .Z(new_n868));
  NOR3_X1   g0668(.A1(new_n359), .A2(new_n221), .A3(new_n307), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT100), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n869), .A2(new_n870), .B1(new_n280), .B2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n283), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n380), .A2(new_n272), .ZN(new_n875));
  INV_X1    g0675(.A(new_n343), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n385), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n341), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT101), .ZN(new_n879));
  INV_X1    g0679(.A(new_n678), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n881), .B(new_n341), .C1(new_n875), .C2(new_n877), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n399), .A3(new_n882), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n884), .A3(new_n409), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n404), .A2(new_n399), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n404), .A2(new_n880), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n409), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n883), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n644), .B2(new_n642), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n409), .B1(new_n388), .B2(new_n400), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n388), .A2(new_n678), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n890), .A2(new_n897), .B1(new_n413), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n898), .B2(KEYINPUT38), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n891), .A2(new_n893), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(KEYINPUT39), .A3(new_n894), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n459), .A2(new_n460), .A3(new_n681), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n644), .A2(new_n678), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n459), .A2(new_n460), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n460), .A2(new_n680), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n443), .A3(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n460), .B(new_n680), .C1(new_n459), .C2(new_n444), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n673), .A2(new_n319), .A3(new_n680), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n833), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n891), .B2(new_n893), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n909), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n908), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n645), .A2(new_n646), .ZN(new_n922));
  INV_X1    g0722(.A(new_n462), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n710), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n921), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n904), .A2(new_n894), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n737), .A2(new_n738), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n741), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n914), .A2(new_n929), .A3(new_n834), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT40), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n914), .A2(new_n929), .A3(KEYINPUT40), .A4(new_n834), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n899), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n929), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n462), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n711), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n925), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n283), .B2(new_n746), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n925), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n874), .B1(new_n941), .B2(new_n942), .ZN(G367));
  OAI221_X1 g0743(.A(new_n764), .B1(new_n215), .B2(new_n305), .C1(new_n756), .C2(new_n232), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n418), .B1(new_n275), .B2(new_n777), .C1(new_n772), .C2(new_n786), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n797), .B2(G50), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n791), .A2(G77), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n775), .A2(new_n344), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G143), .B2(new_n769), .ZN(new_n949));
  INV_X1    g0749(.A(G137), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n781), .A2(new_n358), .B1(new_n785), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT106), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT107), .Z(new_n954));
  AOI22_X1  g0754(.A1(new_n769), .A2(G311), .B1(new_n791), .B2(G97), .ZN(new_n955));
  INV_X1    g0755(.A(G294), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n955), .B1(new_n476), .B2(new_n775), .C1(new_n956), .C2(new_n772), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n797), .A2(G283), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n781), .A2(new_n850), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT46), .Z(new_n960));
  INV_X1    g0760(.A(new_n785), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n845), .A2(G303), .B1(new_n961), .B2(G317), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n958), .A2(new_n960), .A3(new_n755), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n954), .B1(new_n957), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT108), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n749), .B(new_n944), .C1(new_n966), .C2(new_n841), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n598), .A2(new_n680), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n649), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n593), .B2(new_n970), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n968), .B(new_n969), .C1(new_n820), .C2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n566), .B(new_n610), .C1(new_n563), .C2(new_n681), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n703), .A2(new_n680), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT103), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT103), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(new_n508), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n681), .B1(new_n981), .B2(new_n703), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT42), .ZN(new_n983));
  INV_X1    g0783(.A(new_n976), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n691), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT104), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n985), .B2(new_n983), .ZN(new_n987));
  NOR4_X1   g0787(.A1(new_n691), .A2(KEYINPUT104), .A3(KEYINPUT42), .A4(new_n984), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n982), .B1(new_n983), .B2(new_n985), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n689), .A2(new_n979), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT102), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT102), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n689), .A2(new_n994), .A3(new_n979), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n996), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(new_n990), .A3(new_n989), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n747), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n691), .A2(new_n692), .A3(new_n976), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT44), .B1(new_n693), .B2(new_n984), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1012), .B(new_n976), .C1(new_n691), .C2(new_n692), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n689), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n689), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n1011), .B2(new_n1013), .C1(new_n1010), .C2(new_n1009), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n687), .A2(new_n688), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n691), .B1(new_n1019), .B2(new_n690), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n745), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n743), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n743), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n696), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1006), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n973), .B1(new_n1005), .B2(new_n1027), .ZN(G387));
  NAND3_X1  g0828(.A1(new_n687), .A2(new_n688), .A3(new_n762), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n752), .A2(new_n695), .B1(G107), .B2(new_n215), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n229), .A2(new_n259), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n695), .ZN(new_n1032));
  AOI211_X1 g0832(.A(G45), .B(new_n1032), .C1(G68), .C2(G77), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n273), .A2(G50), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n756), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1030), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n749), .B1(new_n1037), .B2(new_n765), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n305), .A2(new_n775), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G159), .B2(new_n769), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n777), .A2(new_n280), .B1(new_n793), .B2(new_n344), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G150), .B2(new_n961), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n755), .B1(G97), .B2(new_n791), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n771), .A2(new_n302), .B1(new_n843), .B2(G77), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n775), .A2(new_n800), .B1(new_n781), .B2(new_n956), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G311), .A2(new_n771), .B1(new_n845), .B2(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n809), .B2(new_n770), .C1(new_n796), .C2(new_n815), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n961), .A2(G326), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n755), .B(new_n1054), .C1(new_n850), .C2(new_n790), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT110), .Z(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1045), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1038), .B1(new_n1058), .B2(new_n763), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1021), .A2(new_n1006), .B1(new_n1029), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n696), .B(KEYINPUT111), .Z(new_n1061));
  NAND2_X1  g0861(.A1(new_n1022), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1021), .A2(new_n743), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(G393));
  NAND3_X1  g0864(.A1(new_n1015), .A2(new_n1017), .A3(new_n1006), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n764), .B1(new_n557), .B2(new_n215), .C1(new_n756), .C2(new_n239), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n749), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n775), .A2(new_n307), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n772), .A2(new_n280), .B1(new_n781), .B2(new_n344), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G87), .C2(new_n791), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n770), .A2(new_n275), .B1(new_n786), .B2(new_n777), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n797), .A2(new_n302), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n755), .B1(G143), .B2(new_n961), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n781), .A2(new_n800), .B1(new_n785), .B2(new_n809), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT112), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G116), .A2(new_n812), .B1(new_n771), .B2(G303), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n244), .B1(new_n793), .B2(new_n956), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G107), .B2(new_n791), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(KEYINPUT112), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G317), .A2(new_n769), .B1(new_n845), .B2(G311), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1075), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1067), .B1(new_n1085), .B2(new_n763), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n979), .B2(new_n820), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1061), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1065), .B(new_n1087), .C1(new_n1088), .C2(new_n1089), .ZN(G390));
  NAND4_X1  g0890(.A1(new_n914), .A2(new_n929), .A3(G330), .A4(new_n834), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(KEYINPUT113), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n916), .A2(new_n907), .B1(new_n901), .B2(new_n905), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n833), .B1(new_n708), .B2(new_n830), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n914), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n907), .B(new_n899), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n827), .B2(new_n832), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n907), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n917), .A2(new_n918), .A3(new_n900), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n897), .A2(new_n890), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n413), .A2(new_n896), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n903), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT39), .B1(new_n1105), .B2(new_n894), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1099), .A2(new_n1100), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n929), .A2(G330), .A3(new_n834), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT113), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n742), .A2(new_n834), .A3(new_n914), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1107), .A2(new_n1096), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1098), .A2(new_n1006), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n906), .A2(new_n760), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n839), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n749), .B1(new_n1116), .B2(new_n302), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n476), .A2(new_n772), .B1(new_n770), .B2(new_n800), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1068), .B(new_n1118), .C1(G68), .C2(new_n791), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n797), .A2(G97), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n807), .A2(G294), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n418), .B(new_n782), .C1(G116), .C2(new_n845), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n772), .A2(new_n950), .B1(new_n790), .B2(new_n280), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n244), .B(new_n1124), .C1(G159), .C2(new_n812), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n807), .A2(G125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n796), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n781), .A2(new_n275), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G128), .A2(new_n769), .B1(new_n845), .B2(G132), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT116), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1123), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1117), .B1(new_n1134), .B2(new_n763), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1115), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1114), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT117), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1114), .A2(new_n1139), .A3(new_n1136), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n462), .A2(new_n936), .A3(new_n711), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n922), .B(new_n1142), .C1(new_n710), .C2(new_n923), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n827), .A2(new_n832), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n914), .B1(new_n742), .B2(new_n834), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT114), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1091), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(KEYINPUT114), .B(new_n914), .C1(new_n742), .C2(new_n834), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1108), .A2(new_n1095), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(new_n1094), .A3(new_n1111), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT115), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1094), .A3(KEYINPUT115), .A4(new_n1111), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1149), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1098), .A2(new_n1113), .A3(new_n1143), .A4(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n1061), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1098), .A2(new_n1113), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1141), .A2(new_n1161), .ZN(G378));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n1143), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT38), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n917), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(G330), .B1(new_n1165), .B2(new_n933), .ZN(new_n1166));
  OAI21_X1  g0966(.A(KEYINPUT120), .B1(new_n1166), .B2(new_n932), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT40), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n919), .B2(new_n930), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n711), .B1(new_n934), .B2(new_n899), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT120), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n640), .A2(new_n646), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n294), .A2(new_n880), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT55), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n1173), .B(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1167), .A2(new_n1172), .A3(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(KEYINPUT120), .C1(new_n932), .C2(new_n1166), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n921), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n921), .A3(new_n1181), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1163), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT57), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1163), .A2(new_n1184), .A3(KEYINPUT57), .A4(new_n1185), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1061), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(new_n1006), .A3(new_n1185), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n748), .B1(new_n280), .B2(new_n839), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n771), .A2(G132), .ZN(new_n1193));
  INV_X1    g0993(.A(G125), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n770), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n845), .A2(G128), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n793), .B2(new_n950), .C1(new_n781), .C2(new_n1127), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G150), .C2(new_n812), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(G33), .A2(G41), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT118), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n790), .A2(new_n786), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G124), .C2(new_n961), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n305), .A2(new_n793), .B1(new_n476), .B2(new_n777), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1207), .A2(new_n948), .A3(G41), .A4(new_n394), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n800), .B2(new_n847), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n770), .A2(new_n850), .B1(new_n781), .B2(new_n307), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n772), .A2(new_n557), .B1(new_n790), .B2(new_n358), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT58), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT58), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n280), .B(new_n1203), .C1(new_n394), .C2(G41), .ZN(new_n1215));
  AND4_X1   g1015(.A1(new_n1206), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1192), .B1(new_n841), .B2(new_n1216), .C1(new_n1178), .C2(new_n761), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1191), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1190), .A2(new_n1219), .ZN(G375));
  INV_X1    g1020(.A(new_n1143), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1155), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n1026), .A3(new_n1159), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1095), .A2(new_n760), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n749), .B1(new_n1116), .B2(G68), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n850), .A2(new_n772), .B1(new_n770), .B2(new_n956), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1039), .B(new_n1227), .C1(G97), .C2(new_n843), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n947), .B(new_n244), .C1(new_n800), .C2(new_n777), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G303), .B2(new_n807), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n476), .C2(new_n796), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT121), .Z(new_n1232));
  OAI21_X1  g1032(.A(new_n394), .B1(new_n358), .B2(new_n790), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT122), .Z(new_n1234));
  OAI22_X1  g1034(.A1(new_n772), .A2(new_n1127), .B1(new_n280), .B2(new_n775), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G159), .B2(new_n843), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n807), .A2(G128), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n777), .A2(new_n950), .B1(new_n793), .B2(new_n275), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G132), .B2(new_n769), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1232), .B1(new_n1234), .B2(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT123), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n841), .B1(new_n1241), .B2(KEYINPUT123), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1226), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1155), .A2(new_n1006), .B1(new_n1225), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1224), .A2(new_n1245), .ZN(G381));
  AND2_X1   g1046(.A1(new_n1189), .A2(new_n1061), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1218), .B1(new_n1247), .B2(new_n1188), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1138), .A2(new_n1140), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G387), .A2(new_n1250), .A3(new_n1251), .A4(G381), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  AOI21_X1  g1053(.A(new_n1249), .B1(new_n1190), .B2(new_n1219), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1186), .A2(new_n1025), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(G378), .A2(new_n1255), .A3(new_n1218), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT124), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1219), .B(new_n1249), .C1(new_n1025), .C2(new_n1186), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n679), .A2(G213), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G384), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1223), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1221), .A2(new_n1222), .A3(KEYINPUT60), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n1061), .A3(new_n1159), .A4(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n838), .A2(KEYINPUT125), .A3(new_n861), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1245), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1263), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(new_n1269), .A3(new_n1263), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1257), .A2(new_n1260), .A3(new_n1261), .A4(new_n1273), .ZN(new_n1274));
  XOR2_X1   g1074(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(G393), .B(new_n822), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1004), .B(new_n1003), .C1(new_n1279), .C2(new_n1006), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G390), .B1(new_n1280), .B2(new_n973), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G390), .B(new_n973), .C1(new_n1005), .C2(new_n1027), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G390), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G387), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n1277), .A3(new_n1282), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(KEYINPUT61), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1257), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1261), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(G2897), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT127), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1292), .A2(KEYINPUT127), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1272), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1293), .B(new_n1294), .C1(new_n1295), .C2(new_n1270), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1271), .A2(KEYINPUT127), .A3(new_n1272), .A4(new_n1292), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1290), .A2(new_n1299), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1254), .A2(new_n1256), .A3(new_n1291), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(KEYINPUT63), .A3(new_n1273), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1276), .A2(new_n1289), .A3(new_n1300), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT62), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1274), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1301), .A2(KEYINPUT62), .A3(new_n1273), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1305), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1288), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1303), .B1(new_n1309), .B2(new_n1310), .ZN(G405));
  INV_X1    g1111(.A(new_n1254), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1250), .A2(new_n1312), .A3(new_n1273), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1273), .B1(new_n1312), .B2(new_n1250), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(new_n1310), .ZN(G402));
endmodule


