//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT72), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT32), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT30), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI22_X1  g011(.A1(new_n195), .A2(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  XNOR2_X1  g013(.A(G134), .B(G137), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n198), .B(new_n199), .C1(new_n200), .C2(new_n196), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n199), .B2(new_n200), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(G143), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n207), .A2(new_n208), .A3(G128), .A4(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT65), .B1(new_n203), .B2(G143), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT64), .B(G146), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n206), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(KEYINPUT65), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n208), .B1(new_n214), .B2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n215), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n212), .B1(new_n221), .B2(KEYINPUT68), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G128), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n215), .A4(new_n218), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n202), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n209), .B1(new_n214), .B2(G143), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n228), .A2(KEYINPUT66), .A3(KEYINPUT0), .A4(G128), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n207), .A2(KEYINPUT0), .A3(G128), .A4(new_n210), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n203), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n216), .B2(new_n217), .ZN(new_n237));
  AOI211_X1 g051(.A(new_n235), .B(G143), .C1(new_n204), .C2(new_n206), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT0), .B(G128), .Z(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n200), .A2(new_n196), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n197), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(new_n196), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n194), .ZN(new_n245));
  OAI21_X1  g059(.A(G131), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n201), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n233), .A2(new_n241), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n193), .B1(new_n227), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n215), .A2(new_n218), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n220), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT68), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n226), .A3(new_n211), .ZN(new_n253));
  INV_X1    g067(.A(new_n202), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n232), .A2(new_n229), .B1(new_n239), .B2(new_n240), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n247), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(KEYINPUT69), .A2(G116), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT69), .A2(G116), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(G119), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT2), .B(G113), .Z(new_n267));
  NAND4_X1  g081(.A1(new_n262), .A2(KEYINPUT70), .A3(G119), .A4(new_n263), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n249), .A2(new_n258), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  INV_X1    g087(.A(G237), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(G210), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n276), .B(KEYINPUT27), .Z(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G101), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n253), .A2(new_n254), .B1(new_n256), .B2(new_n247), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n269), .A2(new_n270), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n272), .A2(new_n273), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n273), .B1(new_n272), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n271), .B1(new_n227), .B2(new_n248), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n255), .A2(new_n281), .A3(new_n257), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT28), .B1(new_n280), .B2(new_n281), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n279), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n192), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n272), .A2(new_n282), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT31), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n272), .A2(new_n273), .A3(new_n282), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n291), .A3(new_n192), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n191), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G472), .ZN(new_n299));
  INV_X1    g113(.A(new_n289), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  INV_X1    g115(.A(new_n290), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n279), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT29), .B1(new_n289), .B2(new_n290), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n272), .A2(new_n301), .A3(new_n288), .A4(new_n279), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT73), .B(G902), .Z(new_n308));
  AND2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n299), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n298), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n294), .A2(new_n291), .A3(new_n295), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT71), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n296), .ZN(new_n315));
  INV_X1    g129(.A(new_n189), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT32), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n187), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n220), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n211), .B1(new_n228), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G104), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G107), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n321), .A2(G107), .ZN(new_n324));
  OAI21_X1  g138(.A(G101), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n321), .B2(G107), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  INV_X1    g141(.A(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G104), .ZN(new_n329));
  INV_X1    g143(.A(G101), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n329), .A3(new_n330), .A4(new_n322), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT10), .B1(new_n320), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n326), .A2(new_n329), .A3(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G101), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n335), .A2(KEYINPUT81), .A3(new_n336), .A4(G101), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(G101), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n339), .A2(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n334), .B1(new_n256), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n247), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n333), .A2(KEYINPUT10), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n253), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n252), .A2(new_n226), .A3(new_n211), .A4(new_n332), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n320), .A2(new_n333), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT12), .B1(new_n351), .B2(new_n247), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT12), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n353), .B(new_n345), .C1(new_n349), .C2(new_n350), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G140), .ZN(new_n356));
  INV_X1    g170(.A(G227), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(G953), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n359), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n345), .B1(new_n344), .B2(new_n347), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n355), .A2(new_n359), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G469), .B1(new_n364), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n366));
  INV_X1    g180(.A(new_n359), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n348), .B(new_n367), .C1(new_n352), .C2(new_n354), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G469), .ZN(new_n371));
  AND4_X1   g185(.A1(new_n366), .A2(new_n370), .A3(new_n371), .A4(new_n308), .ZN(new_n372));
  INV_X1    g186(.A(new_n308), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n366), .B1(new_n374), .B2(new_n371), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n365), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G221), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT9), .B(G234), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G902), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G214), .B1(G237), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n266), .A2(new_n268), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n260), .ZN(new_n389));
  INV_X1    g203(.A(G113), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n333), .ZN(new_n394));
  XNOR2_X1  g208(.A(G110), .B(G122), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n339), .A2(new_n340), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n341), .A2(new_n342), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n394), .B(new_n395), .C1(new_n281), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n271), .A2(new_n343), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n395), .B1(new_n401), .B2(new_n394), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(G125), .B1(new_n222), .B2(new_n226), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n233), .A2(new_n241), .A3(G125), .ZN(new_n405));
  OAI211_X1 g219(.A(G224), .B(new_n275), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G125), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n253), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n256), .A2(G125), .ZN(new_n409));
  INV_X1    g223(.A(G224), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(G953), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g226(.A(KEYINPUT6), .B(new_n395), .C1(new_n401), .C2(new_n394), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n403), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT7), .B1(new_n410), .B2(G953), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n404), .B2(new_n405), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(new_n409), .A3(new_n415), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n395), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n393), .A2(new_n333), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n266), .A2(KEYINPUT5), .A3(new_n268), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n391), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n333), .B1(new_n392), .B2(new_n393), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n417), .A2(new_n418), .A3(new_n425), .A4(new_n399), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n380), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n386), .B1(new_n414), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n400), .A2(new_n402), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n394), .B1(new_n398), .B2(new_n281), .ZN(new_n430));
  INV_X1    g244(.A(new_n395), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n399), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n429), .A2(new_n433), .A3(new_n411), .A4(new_n406), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n434), .A2(new_n380), .A3(new_n385), .A4(new_n426), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n384), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n376), .A2(new_n382), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n321), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n274), .A2(new_n275), .A3(G214), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(G143), .ZN(new_n442));
  AND2_X1   g256(.A1(KEYINPUT18), .A2(G131), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(KEYINPUT76), .A2(G125), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(new_n203), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n407), .A2(G140), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n447), .A2(G125), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n447), .A2(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n407), .A2(G140), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT77), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT78), .B1(new_n458), .B2(new_n214), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n460), .B(new_n216), .C1(new_n454), .C2(new_n457), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n450), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT85), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT77), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT77), .B1(new_n455), .B2(new_n456), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n460), .B1(new_n466), .B2(new_n216), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n458), .A2(KEYINPUT78), .A3(new_n214), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n450), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n445), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT16), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n455), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n448), .B2(new_n473), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(new_n203), .ZN(new_n476));
  INV_X1    g290(.A(new_n442), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G131), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n442), .A2(new_n199), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(KEYINPUT17), .A3(G131), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n440), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n470), .B1(new_n469), .B2(new_n450), .ZN(new_n486));
  AOI211_X1 g300(.A(KEYINPUT85), .B(new_n449), .C1(new_n467), .C2(new_n468), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n444), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n439), .B(KEYINPUT86), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n483), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT88), .B(G475), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n472), .A2(new_n484), .A3(new_n489), .ZN(new_n495));
  MUX2_X1   g309(.A(new_n466), .B(new_n448), .S(KEYINPUT19), .Z(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n214), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n475), .A2(G146), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n478), .A2(new_n479), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n439), .B1(new_n488), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT87), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n500), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n440), .B1(new_n503), .B2(new_n472), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n491), .ZN(new_n506));
  NOR2_X1   g320(.A1(G475), .A2(G902), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n491), .ZN(new_n510));
  NOR3_X1   g324(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n494), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n262), .A2(G122), .A3(new_n263), .ZN(new_n517));
  INV_X1    g331(.A(G122), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G116), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n328), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n521), .A3(new_n519), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n262), .A2(KEYINPUT14), .A3(G122), .A4(new_n263), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G107), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT89), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n217), .B2(G128), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n220), .A2(KEYINPUT89), .A3(G143), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n528), .A2(new_n529), .B1(G128), .B2(new_n217), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(G134), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n516), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n517), .A2(new_n328), .A3(new_n519), .ZN(new_n533));
  INV_X1    g347(.A(new_n525), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n522), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n530), .B(new_n197), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(KEYINPUT90), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n530), .B1(new_n539), .B2(new_n197), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n328), .B1(new_n517), .B2(new_n519), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(new_n533), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT13), .B1(new_n528), .B2(new_n529), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n530), .A2(new_n543), .A3(new_n197), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT91), .ZN(new_n548));
  INV_X1    g362(.A(G217), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n378), .A2(new_n549), .A3(G953), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n545), .B1(new_n532), .B2(new_n537), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n547), .A2(KEYINPUT91), .A3(new_n550), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n308), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT92), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n554), .A2(new_n558), .A3(new_n308), .A4(new_n555), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n515), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n515), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G952), .ZN(new_n564));
  AOI211_X1 g378(.A(G953), .B(new_n564), .C1(G234), .C2(G237), .ZN(new_n565));
  INV_X1    g379(.A(G234), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n373), .B(G953), .C1(new_n566), .C2(new_n274), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT93), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT21), .B(G898), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT94), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n565), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n513), .A2(new_n563), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n437), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n316), .B1(new_n292), .B2(new_n297), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n190), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n310), .B1(new_n315), .B2(new_n191), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT74), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n549), .B1(new_n308), .B2(G234), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n580), .B(KEYINPUT75), .Z(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n220), .A2(G119), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT23), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n220), .A2(KEYINPUT23), .A3(G119), .ZN(new_n587));
  INV_X1    g401(.A(G110), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n259), .A2(G128), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n589), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT24), .B(G110), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n475), .A2(G146), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n469), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n591), .A2(new_n592), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n586), .A2(new_n589), .A3(new_n587), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(G110), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n475), .A2(G146), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n498), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n583), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n498), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n598), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n469), .A2(new_n594), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(KEYINPUT79), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT22), .B(G137), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n377), .A2(new_n566), .A3(G953), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n602), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n604), .A2(new_n605), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n583), .A3(new_n609), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT25), .B1(new_n614), .B2(new_n308), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT25), .ZN(new_n616));
  AOI211_X1 g430(.A(new_n616), .B(new_n373), .C1(new_n611), .C2(new_n613), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n582), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT80), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n580), .A2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n611), .A2(KEYINPUT80), .A3(new_n613), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n318), .A2(new_n575), .A3(new_n579), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  AOI21_X1  g440(.A(new_n373), .B1(new_n314), .B2(new_n296), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n576), .B1(new_n627), .B2(new_n299), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n376), .A2(new_n624), .A3(new_n382), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n556), .A2(new_n514), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n547), .A2(KEYINPUT95), .A3(new_n550), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n550), .B1(new_n547), .B2(KEYINPUT95), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT33), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n554), .A2(new_n555), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n635), .B1(new_n636), .B2(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n308), .A2(G478), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n508), .A2(KEYINPUT20), .B1(new_n510), .B2(new_n511), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n639), .B1(new_n640), .B2(new_n494), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n436), .A2(new_n573), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n631), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n509), .A2(new_n512), .ZN(new_n644));
  INV_X1    g458(.A(new_n494), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n384), .B(new_n572), .C1(new_n428), .C2(new_n435), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT96), .A4(new_n639), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n630), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT97), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  OR2_X1    g466(.A1(new_n560), .A2(new_n562), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n502), .A2(new_n506), .A3(new_n511), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n494), .B1(new_n509), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n647), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n628), .A2(new_n656), .A3(new_n629), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n612), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n621), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n618), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n660), .B1(new_n628), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n315), .A2(new_n308), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n576), .A4(new_n664), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n666), .A2(new_n669), .A3(new_n575), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NOR2_X1   g486(.A1(new_n437), .A2(new_n665), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n565), .B1(new_n568), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n653), .A2(new_n655), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n318), .A2(new_n579), .A3(new_n673), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  NAND2_X1  g494(.A1(new_n374), .A2(new_n371), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT82), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n374), .A2(new_n366), .A3(new_n371), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n381), .B1(new_n684), .B2(new_n365), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n675), .B(KEYINPUT39), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT40), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n272), .A2(new_n288), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n304), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n287), .A2(new_n288), .A3(new_n279), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n380), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n299), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n315), .B2(new_n191), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n664), .B1(new_n577), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n428), .A2(new_n435), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  OAI22_X1  g511(.A1(new_n640), .A2(new_n494), .B1(new_n560), .B2(new_n562), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n384), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n688), .A2(new_n695), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n217), .ZN(G45));
  OAI211_X1 g515(.A(new_n639), .B(new_n676), .C1(new_n640), .C2(new_n494), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n318), .A2(new_n579), .A3(new_n673), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT99), .B(G146), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G48));
  NAND2_X1  g520(.A1(new_n318), .A2(new_n579), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n374), .A2(new_n371), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n624), .A2(new_n684), .A3(new_n382), .A4(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n643), .A3(new_n648), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT41), .B(G113), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT100), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n712), .B(new_n714), .ZN(G15));
  NOR2_X1   g529(.A1(new_n656), .A2(new_n709), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n318), .A3(new_n579), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NOR2_X1   g532(.A1(new_n574), .A2(new_n665), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n684), .A2(new_n382), .A3(new_n708), .ZN(new_n720));
  INV_X1    g534(.A(new_n436), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n318), .A2(new_n579), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NOR2_X1   g538(.A1(new_n709), .A2(new_n572), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n646), .A2(KEYINPUT103), .A3(new_n653), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n721), .B1(new_n698), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n300), .A2(new_n729), .A3(new_n302), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT101), .B1(new_n289), .B2(new_n290), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n279), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n189), .B1(new_n732), .B2(new_n285), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT102), .B(G472), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n667), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n725), .A2(new_n726), .A3(new_n728), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NAND4_X1  g551(.A1(new_n722), .A2(new_n735), .A3(new_n664), .A4(new_n703), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND2_X1  g553(.A1(new_n577), .A2(new_n578), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n624), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(KEYINPUT107), .A3(new_n624), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n361), .A2(new_n363), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n355), .A2(KEYINPUT105), .A3(new_n359), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT105), .B1(new_n355), .B2(new_n359), .ZN(new_n748));
  OAI211_X1 g562(.A(G469), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(G469), .A2(G902), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT104), .Z(new_n751));
  OAI211_X1 g565(.A(new_n749), .B(new_n751), .C1(new_n372), .C2(new_n375), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n382), .A2(new_n428), .A3(new_n383), .A4(new_n435), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n754), .A2(new_n702), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n745), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n754), .A2(new_n702), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n318), .A2(new_n579), .A3(new_n758), .A4(new_n624), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n755), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NAND3_X1  g578(.A1(new_n318), .A2(new_n624), .A3(new_n579), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n677), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n653), .A2(new_n655), .A3(KEYINPUT108), .A4(new_n676), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n752), .A3(new_n753), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n197), .ZN(G36));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n513), .A2(new_n639), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n628), .A2(new_n664), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OR4_X1    g592(.A1(new_n772), .A2(new_n774), .A3(new_n777), .A4(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n696), .A2(new_n384), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n776), .B2(new_n777), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n364), .A2(KEYINPUT45), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n371), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT109), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT109), .B(G469), .C1(new_n364), .C2(KEYINPUT45), .ZN(new_n789));
  OAI211_X1 g603(.A(KEYINPUT45), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT110), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n793), .B(new_n794), .C1(KEYINPUT109), .C2(new_n787), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n751), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n799), .A3(KEYINPUT46), .A4(new_n751), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT46), .B1(new_n796), .B2(new_n751), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n798), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n801), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n684), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n382), .B(new_n686), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n785), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  OAI21_X1  g623(.A(new_n382), .B1(new_n803), .B2(new_n805), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT47), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n382), .C1(new_n803), .C2(new_n805), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n318), .A2(new_n579), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n814), .A2(new_n624), .A3(new_n702), .A4(new_n782), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  AND2_X1   g631(.A1(new_n684), .A2(new_n708), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT49), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n577), .A2(new_n624), .A3(new_n694), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n697), .A2(new_n773), .A3(new_n381), .A4(new_n384), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n811), .A2(new_n813), .B1(new_n381), .B2(new_n818), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n773), .B(KEYINPUT43), .Z(new_n824));
  NAND3_X1  g638(.A1(new_n735), .A2(new_n624), .A3(new_n565), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n782), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n697), .A2(new_n383), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n827), .A2(new_n720), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT50), .ZN(new_n834));
  INV_X1    g648(.A(new_n565), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n720), .A2(new_n782), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n820), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT118), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n646), .A2(new_n639), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n824), .A2(new_n836), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n664), .A3(new_n735), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n834), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT51), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n823), .B2(new_n829), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT119), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n745), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT48), .ZN(new_n849));
  INV_X1    g663(.A(new_n641), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n838), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n827), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n564), .B(G953), .C1(new_n852), .C2(new_n722), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n845), .B2(new_n846), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n844), .A2(new_n847), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n675), .B1(new_n618), .B2(new_n663), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n563), .A2(new_n781), .A3(new_n655), .A4(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n318), .A2(new_n579), .A3(new_n685), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n758), .A2(new_n664), .A3(new_n735), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n860), .B(new_n861), .C1(new_n765), .C2(new_n769), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n641), .B2(new_n642), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT115), .A4(new_n639), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n653), .A2(new_n647), .A3(new_n513), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n630), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n670), .A2(new_n868), .A3(new_n625), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n723), .A2(new_n736), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n710), .A2(new_n643), .A3(new_n648), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n814), .B1(new_n872), .B2(new_n716), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n717), .B1(new_n707), .B2(new_n711), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n723), .A2(new_n736), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT114), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n870), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n762), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT42), .B1(new_n759), .B2(KEYINPUT106), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n880), .A2(new_n881), .B1(new_n745), .B2(new_n756), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n679), .A2(new_n738), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n752), .A2(new_n382), .A3(new_n676), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n695), .A2(new_n885), .A3(new_n726), .A4(new_n728), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n884), .A2(KEYINPUT52), .A3(new_n704), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n679), .A2(new_n704), .A3(new_n886), .A4(new_n738), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n883), .B(new_n891), .C1(KEYINPUT116), .C2(KEYINPUT53), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n875), .A2(new_n878), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n763), .A3(new_n891), .A4(new_n870), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT53), .B1(new_n891), .B2(KEYINPUT116), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n857), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT53), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n763), .A2(new_n870), .A3(new_n878), .A4(new_n875), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n887), .A2(new_n890), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n876), .A2(new_n877), .A3(new_n898), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n891), .A2(new_n902), .A3(new_n763), .A4(new_n870), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n901), .A2(new_n857), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT117), .B1(new_n897), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n894), .A2(new_n895), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n894), .A2(new_n895), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT54), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n901), .A2(new_n857), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n856), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n822), .B1(new_n912), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n275), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n901), .A2(new_n903), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n308), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(new_n386), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n429), .A2(new_n433), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n412), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n434), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT55), .Z(new_n924));
  OAI21_X1  g738(.A(new_n916), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n920), .B2(new_n924), .ZN(G51));
  NAND2_X1  g740(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(KEYINPUT120), .B2(new_n910), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n910), .A2(KEYINPUT120), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n751), .B(KEYINPUT57), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n370), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n919), .A2(new_n795), .A3(new_n792), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n915), .B1(new_n933), .B2(new_n934), .ZN(G54));
  NAND3_X1  g749(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n502), .A2(new_n506), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n936), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n915), .ZN(G60));
  XNOR2_X1  g755(.A(new_n637), .B(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n857), .B1(new_n901), .B2(new_n903), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n904), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n949), .B2(new_n929), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT122), .B1(new_n950), .B2(new_n915), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n945), .B1(new_n928), .B2(new_n930), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n952), .A2(new_n953), .A3(new_n916), .ZN(new_n954));
  INV_X1    g768(.A(new_n944), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n911), .A2(new_n905), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n942), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n951), .A2(new_n954), .A3(new_n957), .ZN(G63));
  OAI21_X1  g772(.A(new_n916), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n918), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n962), .B2(new_n662), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n620), .A2(new_n622), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n918), .B2(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G66));
  AOI21_X1  g782(.A(new_n275), .B1(new_n570), .B2(G224), .ZN(new_n969));
  INV_X1    g783(.A(new_n869), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n893), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n972), .B2(new_n275), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n921), .B1(G898), .B2(new_n275), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT124), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  NAND3_X1  g790(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n850), .B1(new_n513), .B2(new_n653), .ZN(new_n978));
  NOR4_X1   g792(.A1(new_n765), .A2(new_n978), .A3(new_n687), .A4(new_n782), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n884), .A2(new_n704), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n700), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n808), .A3(new_n816), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n977), .B1(new_n986), .B2(G953), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n249), .A2(new_n258), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n496), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n882), .A2(new_n770), .A3(new_n980), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n745), .A2(new_n726), .A3(new_n728), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n780), .B2(new_n783), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n994), .B2(new_n806), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n990), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n994), .A2(new_n806), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n997), .A2(new_n816), .A3(KEYINPUT125), .A4(new_n992), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n996), .A2(new_n275), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n357), .A2(KEYINPUT126), .A3(G900), .ZN(new_n1000));
  OAI21_X1  g814(.A(G953), .B1(KEYINPUT126), .B2(G900), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n989), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g817(.A1(new_n987), .A2(new_n989), .B1(new_n999), .B2(new_n1003), .ZN(G72));
  NAND2_X1  g818(.A1(new_n892), .A2(new_n896), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n689), .A2(new_n304), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  NAND4_X1  g823(.A1(new_n1005), .A2(new_n1007), .A3(new_n690), .A4(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n985), .A2(new_n808), .A3(new_n816), .A4(new_n971), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1011), .A2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1010), .B1(new_n1012), .B2(new_n690), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n996), .A2(new_n971), .A3(new_n998), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1014), .A2(new_n1009), .ZN(new_n1015));
  OAI211_X1 g829(.A(KEYINPUT127), .B(new_n916), .C1(new_n1015), .C2(new_n1007), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1007), .B1(new_n1014), .B2(new_n1009), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(new_n915), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1013), .B1(new_n1016), .B2(new_n1019), .ZN(G57));
endmodule


