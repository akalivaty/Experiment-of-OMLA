

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U558 ( .A1(n542), .A2(n541), .ZN(G160) );
  XOR2_X1 U559 ( .A(n815), .B(KEYINPUT85), .Z(n525) );
  NOR2_X1 U560 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U561 ( .A1(n726), .A2(n725), .ZN(n727) );
  INV_X1 U562 ( .A(KEYINPUT90), .ZN(n687) );
  XNOR2_X1 U563 ( .A(n731), .B(KEYINPUT96), .ZN(n747) );
  NAND2_X1 U564 ( .A1(n816), .A2(n525), .ZN(n817) );
  BUF_X1 U565 ( .A(n684), .Z(G164) );
  INV_X1 U566 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U567 ( .A1(G2104), .A2(n526), .ZN(n904) );
  NAND2_X1 U568 ( .A1(n904), .A2(G126), .ZN(n527) );
  XNOR2_X1 U569 ( .A(n527), .B(KEYINPUT84), .ZN(n530) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XOR2_X2 U571 ( .A(KEYINPUT17), .B(n528), .Z(n901) );
  NAND2_X1 U572 ( .A1(G138), .A2(n901), .ZN(n529) );
  NAND2_X1 U573 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U574 ( .A1(n526), .A2(G2104), .ZN(n531) );
  XNOR2_X2 U575 ( .A(n531), .B(KEYINPUT65), .ZN(n900) );
  NAND2_X1 U576 ( .A1(G102), .A2(n900), .ZN(n533) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n905) );
  NAND2_X1 U578 ( .A1(G114), .A2(n905), .ZN(n532) );
  NAND2_X1 U579 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U580 ( .A1(n535), .A2(n534), .ZN(n684) );
  NAND2_X1 U581 ( .A1(G101), .A2(n900), .ZN(n536) );
  XOR2_X1 U582 ( .A(KEYINPUT23), .B(n536), .Z(n542) );
  NAND2_X1 U583 ( .A1(G125), .A2(n904), .ZN(n538) );
  NAND2_X1 U584 ( .A1(G113), .A2(n905), .ZN(n537) );
  AND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n540) );
  NAND2_X1 U586 ( .A1(n901), .A2(G137), .ZN(n539) );
  AND2_X1 U587 ( .A1(n540), .A2(n539), .ZN(n541) );
  INV_X1 U588 ( .A(G651), .ZN(n546) );
  NOR2_X1 U589 ( .A1(G543), .A2(n546), .ZN(n543) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n543), .Z(n644) );
  NAND2_X1 U591 ( .A1(G65), .A2(n644), .ZN(n545) );
  NOR2_X1 U592 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U593 ( .A1(G91), .A2(n650), .ZN(n544) );
  NAND2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n550) );
  XOR2_X1 U595 ( .A(KEYINPUT0), .B(G543), .Z(n641) );
  NOR2_X1 U596 ( .A1(n641), .A2(n546), .ZN(n649) );
  NAND2_X1 U597 ( .A1(G78), .A2(n649), .ZN(n548) );
  NOR2_X2 U598 ( .A1(G651), .A2(n641), .ZN(n645) );
  NAND2_X1 U599 ( .A1(G53), .A2(n645), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U601 ( .A1(n550), .A2(n549), .ZN(G299) );
  NAND2_X1 U602 ( .A1(G60), .A2(n644), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G85), .A2(n650), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U605 ( .A1(G72), .A2(n649), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G47), .A2(n645), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U608 ( .A1(n556), .A2(n555), .ZN(G290) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  NAND2_X1 U613 ( .A1(G64), .A2(n644), .ZN(n557) );
  XOR2_X1 U614 ( .A(KEYINPUT66), .B(n557), .Z(n564) );
  NAND2_X1 U615 ( .A1(G77), .A2(n649), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G90), .A2(n650), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U618 ( .A(n560), .B(KEYINPUT9), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G52), .A2(n645), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U621 ( .A1(n564), .A2(n563), .ZN(G171) );
  NAND2_X1 U622 ( .A1(n650), .A2(G89), .ZN(n565) );
  XNOR2_X1 U623 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G76), .A2(n649), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U626 ( .A(n568), .B(KEYINPUT5), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G63), .A2(n644), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G51), .A2(n645), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT6), .B(n571), .Z(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U632 ( .A(n574), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U635 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U636 ( .A(G223), .B(KEYINPUT67), .ZN(n845) );
  NAND2_X1 U637 ( .A1(n845), .A2(G567), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U639 ( .A1(G81), .A2(n650), .ZN(n577) );
  XNOR2_X1 U640 ( .A(n577), .B(KEYINPUT12), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT68), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G68), .A2(n649), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U644 ( .A(n581), .B(KEYINPUT13), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G43), .A2(n645), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n644), .A2(G56), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT14), .B(n584), .Z(n585) );
  NOR2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n985) );
  NAND2_X1 U650 ( .A1(G860), .A2(n985), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT69), .B(n587), .Z(G153) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U654 ( .A1(G92), .A2(n650), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT70), .ZN(n595) );
  NAND2_X1 U656 ( .A1(G79), .A2(n649), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G66), .A2(n644), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U659 ( .A1(G54), .A2(n645), .ZN(n591) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n591), .ZN(n592) );
  NOR2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n596), .Z(n990) );
  INV_X1 U664 ( .A(G868), .ZN(n655) );
  NAND2_X1 U665 ( .A1(n990), .A2(n655), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(G284) );
  NOR2_X1 U667 ( .A1(G286), .A2(n655), .ZN(n600) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U670 ( .A(G860), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n601), .A2(G559), .ZN(n602) );
  INV_X1 U672 ( .A(n990), .ZN(n618) );
  NAND2_X1 U673 ( .A1(n602), .A2(n618), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n603), .B(KEYINPUT72), .ZN(n604) );
  XNOR2_X1 U675 ( .A(KEYINPUT16), .B(n604), .ZN(G148) );
  NAND2_X1 U676 ( .A1(n618), .A2(G868), .ZN(n605) );
  NOR2_X1 U677 ( .A1(G559), .A2(n605), .ZN(n607) );
  AND2_X1 U678 ( .A1(n655), .A2(n985), .ZN(n606) );
  NOR2_X1 U679 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G99), .A2(n900), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G111), .A2(n905), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n904), .A2(G123), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G135), .A2(n901), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U687 ( .A(KEYINPUT73), .B(n613), .Z(n614) );
  NOR2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n930) );
  XNOR2_X1 U689 ( .A(n930), .B(G2096), .ZN(n617) );
  INV_X1 U690 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U692 ( .A1(n618), .A2(G559), .ZN(n666) );
  XOR2_X1 U693 ( .A(n985), .B(KEYINPUT74), .Z(n619) );
  XNOR2_X1 U694 ( .A(n666), .B(n619), .ZN(n620) );
  NOR2_X1 U695 ( .A1(G860), .A2(n620), .ZN(n628) );
  NAND2_X1 U696 ( .A1(G80), .A2(n649), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G67), .A2(n644), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G93), .A2(n650), .ZN(n623) );
  XNOR2_X1 U700 ( .A(KEYINPUT75), .B(n623), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n645), .A2(G55), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n657) );
  XOR2_X1 U704 ( .A(n628), .B(n657), .Z(G145) );
  NAND2_X1 U705 ( .A1(G73), .A2(n649), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n644), .A2(G61), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G86), .A2(n650), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G48), .A2(n645), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U713 ( .A(KEYINPUT77), .B(n636), .ZN(G305) );
  NAND2_X1 U714 ( .A1(G49), .A2(n645), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U717 ( .A(KEYINPUT76), .B(n639), .ZN(n640) );
  NOR2_X1 U718 ( .A1(n644), .A2(n640), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G62), .A2(n644), .ZN(n647) );
  NAND2_X1 U722 ( .A1(G50), .A2(n645), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U724 ( .A(KEYINPUT78), .B(n648), .Z(n654) );
  NAND2_X1 U725 ( .A1(n649), .A2(G75), .ZN(n652) );
  NAND2_X1 U726 ( .A1(G88), .A2(n650), .ZN(n651) );
  AND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(G303) );
  INV_X1 U729 ( .A(G303), .ZN(G166) );
  NAND2_X1 U730 ( .A1(n655), .A2(n657), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n656), .B(KEYINPUT82), .ZN(n670) );
  XNOR2_X1 U732 ( .A(G305), .B(G288), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n985), .B(G166), .ZN(n663) );
  XNOR2_X1 U734 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n657), .B(KEYINPUT79), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U737 ( .A(n660), .B(G299), .Z(n661) );
  XNOR2_X1 U738 ( .A(G290), .B(n661), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(n917) );
  XNOR2_X1 U741 ( .A(KEYINPUT81), .B(n917), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U743 ( .A1(G868), .A2(n668), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(G295) );
  INV_X1 U745 ( .A(G2072), .ZN(n961) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XOR2_X1 U749 ( .A(KEYINPUT21), .B(n673), .Z(n674) );
  NOR2_X1 U750 ( .A1(n961), .A2(n674), .ZN(n675) );
  XNOR2_X1 U751 ( .A(KEYINPUT83), .B(n675), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U755 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U756 ( .A1(G96), .A2(n678), .ZN(n849) );
  NAND2_X1 U757 ( .A1(n849), .A2(G2106), .ZN(n682) );
  NAND2_X1 U758 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U759 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U760 ( .A1(G108), .A2(n680), .ZN(n850) );
  NAND2_X1 U761 ( .A1(n850), .A2(G567), .ZN(n681) );
  NAND2_X1 U762 ( .A1(n682), .A2(n681), .ZN(n851) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U764 ( .A1(n851), .A2(n683), .ZN(n848) );
  NAND2_X1 U765 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n786) );
  INV_X1 U767 ( .A(n786), .ZN(n685) );
  NOR2_X1 U768 ( .A1(n684), .A2(G1384), .ZN(n787) );
  NAND2_X1 U769 ( .A1(n685), .A2(n787), .ZN(n686) );
  XNOR2_X2 U770 ( .A(n686), .B(KEYINPUT64), .ZN(n714) );
  INV_X1 U771 ( .A(n714), .ZN(n699) );
  INV_X1 U772 ( .A(n699), .ZN(n732) );
  NOR2_X1 U773 ( .A1(n732), .A2(G2084), .ZN(n748) );
  NAND2_X1 U774 ( .A1(n714), .A2(G8), .ZN(n733) );
  NOR2_X1 U775 ( .A1(G1966), .A2(n733), .ZN(n688) );
  XNOR2_X1 U776 ( .A(n688), .B(n687), .ZN(n750) );
  NAND2_X1 U777 ( .A1(n750), .A2(G8), .ZN(n689) );
  NOR2_X1 U778 ( .A1(n748), .A2(n689), .ZN(n690) );
  XOR2_X1 U779 ( .A(KEYINPUT30), .B(n690), .Z(n691) );
  NOR2_X1 U780 ( .A1(G168), .A2(n691), .ZN(n692) );
  XNOR2_X1 U781 ( .A(n692), .B(KEYINPUT97), .ZN(n697) );
  XOR2_X1 U782 ( .A(KEYINPUT91), .B(G1961), .Z(n1019) );
  NOR2_X1 U783 ( .A1(n1019), .A2(n699), .ZN(n694) );
  XOR2_X1 U784 ( .A(KEYINPUT25), .B(G2078), .Z(n966) );
  NOR2_X1 U785 ( .A1(n732), .A2(n966), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U787 ( .A(KEYINPUT92), .B(n695), .Z(n728) );
  OR2_X1 U788 ( .A1(n728), .A2(G171), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n698), .B(KEYINPUT31), .ZN(n746) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n699), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n714), .A2(G1348), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n717) );
  NAND2_X1 U794 ( .A1(n717), .A2(n990), .ZN(n711) );
  XNOR2_X1 U795 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n704) );
  OR2_X1 U796 ( .A1(n704), .A2(G1996), .ZN(n702) );
  NAND2_X1 U797 ( .A1(n985), .A2(n702), .ZN(n709) );
  INV_X1 U798 ( .A(G1341), .ZN(n1010) );
  NAND2_X1 U799 ( .A1(n1010), .A2(n704), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n703), .A2(n714), .ZN(n707) );
  INV_X1 U801 ( .A(G1996), .ZN(n957) );
  NOR2_X1 U802 ( .A1(n714), .A2(n957), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n714), .A2(n961), .ZN(n713) );
  XOR2_X1 U808 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n712) );
  XNOR2_X1 U809 ( .A(n713), .B(n712), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n714), .A2(G1956), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n723) );
  NOR2_X1 U812 ( .A1(G299), .A2(n723), .ZN(n719) );
  NOR2_X1 U813 ( .A1(n717), .A2(n990), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U815 ( .A(KEYINPUT95), .B(n722), .ZN(n726) );
  NAND2_X1 U816 ( .A1(G299), .A2(n723), .ZN(n724) );
  XOR2_X1 U817 ( .A(KEYINPUT28), .B(n724), .Z(n725) );
  XNOR2_X1 U818 ( .A(n727), .B(KEYINPUT29), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n728), .A2(G171), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n731) );
  INV_X1 U821 ( .A(G8), .ZN(n738) );
  NOR2_X1 U822 ( .A1(n732), .A2(G2090), .ZN(n735) );
  BUF_X1 U823 ( .A(n733), .Z(n774) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n774), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n740) );
  AND2_X1 U828 ( .A1(n747), .A2(n740), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n746), .A2(n739), .ZN(n744) );
  INV_X1 U830 ( .A(n740), .ZN(n742) );
  AND2_X1 U831 ( .A1(G286), .A2(G8), .ZN(n741) );
  OR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U834 ( .A(n745), .B(KEYINPUT32), .ZN(n771) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n752) );
  NAND2_X1 U836 ( .A1(G8), .A2(n748), .ZN(n749) );
  AND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n769) );
  NAND2_X1 U839 ( .A1(n771), .A2(n769), .ZN(n757) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n981), .A2(n753), .ZN(n754) );
  XNOR2_X1 U843 ( .A(KEYINPUT98), .B(n754), .ZN(n755) );
  INV_X1 U844 ( .A(KEYINPUT33), .ZN(n759) );
  AND2_X1 U845 ( .A1(n755), .A2(n759), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n767) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n983) );
  INV_X1 U848 ( .A(n774), .ZN(n781) );
  NAND2_X1 U849 ( .A1(n983), .A2(n781), .ZN(n758) );
  AND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n981), .A2(KEYINPUT33), .ZN(n760) );
  NOR2_X1 U852 ( .A1(n760), .A2(n774), .ZN(n763) );
  XNOR2_X1 U853 ( .A(G1981), .B(KEYINPUT99), .ZN(n761) );
  XNOR2_X1 U854 ( .A(n761), .B(G305), .ZN(n996) );
  INV_X1 U855 ( .A(n996), .ZN(n762) );
  OR2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U859 ( .A(n768), .B(KEYINPUT100), .Z(n785) );
  AND2_X1 U860 ( .A1(n769), .A2(n774), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G166), .A2(G8), .ZN(n772) );
  NOR2_X1 U863 ( .A1(G2090), .A2(n772), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n777), .B(KEYINPUT101), .ZN(n783) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U868 ( .A(n778), .B(KEYINPUT24), .Z(n779) );
  XNOR2_X1 U869 ( .A(KEYINPUT89), .B(n779), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n818) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n829) );
  NAND2_X1 U874 ( .A1(G129), .A2(n904), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G117), .A2(n905), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n900), .A2(G105), .ZN(n790) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n790), .Z(n791) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U880 ( .A1(n901), .A2(G141), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n888) );
  NAND2_X1 U882 ( .A1(G1996), .A2(n888), .ZN(n803) );
  NAND2_X1 U883 ( .A1(G119), .A2(n904), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G95), .A2(n900), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G107), .A2(n905), .ZN(n797) );
  XNOR2_X1 U887 ( .A(KEYINPUT87), .B(n797), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n901), .A2(G131), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n881) );
  NAND2_X1 U891 ( .A1(G1991), .A2(n881), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n931) );
  NAND2_X1 U893 ( .A1(n829), .A2(n931), .ZN(n821) );
  NAND2_X1 U894 ( .A1(G104), .A2(n900), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G140), .A2(n901), .ZN(n804) );
  NAND2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n806), .ZN(n811) );
  NAND2_X1 U898 ( .A1(G128), .A2(n904), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G116), .A2(n905), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n809), .Z(n810) );
  NOR2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n812), .ZN(n914) );
  XNOR2_X1 U904 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  NOR2_X1 U905 ( .A1(n914), .A2(n827), .ZN(n949) );
  NAND2_X1 U906 ( .A1(n949), .A2(n829), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n813), .B(KEYINPUT86), .ZN(n826) );
  NAND2_X1 U908 ( .A1(n821), .A2(n826), .ZN(n814) );
  XOR2_X1 U909 ( .A(KEYINPUT88), .B(n814), .Z(n816) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U911 ( .A1(n829), .A2(n987), .ZN(n815) );
  OR2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n833) );
  OR2_X1 U913 ( .A1(n888), .A2(G1996), .ZN(n935) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n881), .ZN(n932) );
  NOR2_X1 U916 ( .A1(n819), .A2(n932), .ZN(n820) );
  XOR2_X1 U917 ( .A(KEYINPUT102), .B(n820), .Z(n822) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n935), .A2(n823), .ZN(n824) );
  XOR2_X1 U920 ( .A(KEYINPUT39), .B(n824), .Z(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n914), .A2(n827), .ZN(n947) );
  NAND2_X1 U923 ( .A1(n828), .A2(n947), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U925 ( .A(KEYINPUT103), .B(n831), .Z(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT40), .ZN(n835) );
  XNOR2_X1 U928 ( .A(KEYINPUT104), .B(n835), .ZN(G329) );
  XNOR2_X1 U929 ( .A(G1341), .B(G2454), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(G2430), .ZN(n837) );
  XNOR2_X1 U931 ( .A(n837), .B(G1348), .ZN(n843) );
  XOR2_X1 U932 ( .A(G2443), .B(G2427), .Z(n839) );
  XNOR2_X1 U933 ( .A(G2438), .B(G2446), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(n841) );
  XOR2_X1 U935 ( .A(G2451), .B(G2435), .Z(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n844), .A2(G14), .ZN(n922) );
  XNOR2_X1 U939 ( .A(KEYINPUT105), .B(n922), .ZN(G401) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U942 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U944 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U946 ( .A(G120), .ZN(G236) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  INV_X1 U948 ( .A(G69), .ZN(G235) );
  NOR2_X1 U949 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U950 ( .A(G325), .ZN(G261) );
  INV_X1 U951 ( .A(n851), .ZN(G319) );
  XOR2_X1 U952 ( .A(G2100), .B(G2096), .Z(n853) );
  XNOR2_X1 U953 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2090), .Z(n855) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2678), .B(KEYINPUT106), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n861) );
  XOR2_X1 U961 ( .A(G2078), .B(G2084), .Z(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1986), .B(G1976), .Z(n863) );
  XNOR2_X1 U964 ( .A(G1966), .B(G1971), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n873) );
  XOR2_X1 U966 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U967 ( .A(G1991), .B(G2474), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U969 ( .A(G1996), .B(G1956), .Z(n867) );
  XNOR2_X1 U970 ( .A(G1981), .B(G1961), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U972 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U973 ( .A(KEYINPUT110), .B(KEYINPUT109), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U976 ( .A1(n904), .A2(G124), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G112), .A2(n905), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G100), .A2(n900), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G136), .A2(n901), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(G162) );
  XNOR2_X1 U984 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n881), .B(KEYINPUT111), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(n884), .B(KEYINPUT113), .Z(n886) );
  XNOR2_X1 U988 ( .A(G160), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U990 ( .A(n887), .B(n930), .Z(n890) );
  XOR2_X1 U991 ( .A(n888), .B(G162), .Z(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n899) );
  NAND2_X1 U993 ( .A1(G130), .A2(n904), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G118), .A2(n905), .ZN(n891) );
  NAND2_X1 U995 ( .A1(n892), .A2(n891), .ZN(n897) );
  NAND2_X1 U996 ( .A1(G106), .A2(n900), .ZN(n894) );
  NAND2_X1 U997 ( .A1(G142), .A2(n901), .ZN(n893) );
  NAND2_X1 U998 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U999 ( .A(KEYINPUT45), .B(n895), .Z(n896) );
  NOR2_X1 U1000 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U1001 ( .A(n899), .B(n898), .Z(n913) );
  NAND2_X1 U1002 ( .A1(G103), .A2(n900), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(G139), .A2(n901), .ZN(n902) );
  NAND2_X1 U1004 ( .A1(n903), .A2(n902), .ZN(n911) );
  NAND2_X1 U1005 ( .A1(G127), .A2(n904), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n905), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1008 ( .A(KEYINPUT47), .B(n908), .Z(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT112), .B(n909), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n939) );
  XNOR2_X1 U1011 ( .A(G164), .B(n939), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n916), .ZN(G395) );
  XNOR2_X1 U1015 ( .A(n917), .B(KEYINPUT115), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(G171), .B(G286), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(n990), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n921), .ZN(G397) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n922), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1028 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1040) );
  XOR2_X1 U1029 ( .A(G2084), .B(G160), .Z(n928) );
  XNOR2_X1 U1030 ( .A(KEYINPUT116), .B(n928), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n946) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G162), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(n937), .B(KEYINPUT51), .ZN(n938) );
  XOR2_X1 U1037 ( .A(KEYINPUT117), .B(n938), .Z(n944) );
  XOR2_X1 U1038 ( .A(G164), .B(G2078), .Z(n941) );
  XNOR2_X1 U1039 ( .A(n961), .B(n939), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT50), .B(n942), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n951) );
  INV_X1 U1044 ( .A(n947), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n952), .ZN(n953) );
  XOR2_X1 U1048 ( .A(KEYINPUT118), .B(n953), .Z(n955) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G29), .ZN(n1038) );
  XNOR2_X1 U1052 ( .A(G32), .B(n957), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G25), .B(G1991), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n970) );
  XNOR2_X1 U1056 ( .A(G33), .B(KEYINPUT119), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(n961), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G26), .B(G2067), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1060 ( .A(KEYINPUT120), .B(n965), .Z(n968) );
  XNOR2_X1 U1061 ( .A(n966), .B(G27), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n971), .B(KEYINPUT53), .ZN(n974) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G35), .B(G2090), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1070 ( .A(KEYINPUT55), .B(n977), .Z(n978) );
  NOR2_X1 U1071 ( .A1(G29), .A2(n978), .ZN(n1008) );
  XNOR2_X1 U1072 ( .A(KEYINPUT56), .B(G16), .ZN(n1005) );
  XNOR2_X1 U1073 ( .A(G301), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(G303), .B(G1971), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n1003) );
  INV_X1 U1076 ( .A(n981), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n984), .B(KEYINPUT123), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(G1341), .B(n985), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G299), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1348), .B(n990), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT122), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G168), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n998), .B(KEYINPUT121), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(n999), .B(KEYINPUT57), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(G11), .A2(n1006), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1035) );
  XOR2_X1 U1096 ( .A(KEYINPUT124), .B(G16), .Z(n1033) );
  XNOR2_X1 U1097 ( .A(KEYINPUT125), .B(G1966), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(G21), .ZN(n1023) );
  XNOR2_X1 U1099 ( .A(G19), .B(n1010), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G1981), .B(G6), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G20), .B(G1956), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1105 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT60), .B(n1018), .Z(n1021) );
  XNOR2_X1 U1108 ( .A(n1019), .B(G5), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1030) );
  XNOR2_X1 U1111 ( .A(G1971), .B(G22), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(G24), .B(G1986), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1027) );
  XOR2_X1 U1114 ( .A(G1976), .B(G23), .Z(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT58), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1118 ( .A(KEYINPUT61), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1121 ( .A(KEYINPUT126), .B(n1036), .Z(n1037) );
  NAND2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1123 ( .A(n1040), .B(n1039), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

