//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT27), .B(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n208), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n206), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n204), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT67), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n213), .B2(KEYINPUT23), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT25), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(G169gat), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(KEYINPUT23), .A3(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n203), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n228), .B(new_n230), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n212), .A2(new_n221), .B1(new_n227), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n214), .A2(new_n217), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n222), .B1(new_n237), .B2(KEYINPUT23), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n228), .A3(new_n231), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n230), .A2(new_n228), .A3(KEYINPUT68), .A4(new_n231), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n236), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(G113gat), .B2(G120gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(G113gat), .A2(G120gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(G127gat), .B(G134gat), .Z(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254));
  OR2_X1    g053(.A1(G113gat), .A2(G120gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n247), .A3(new_n249), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n256), .B2(new_n246), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n235), .A2(new_n245), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n251), .A2(new_n252), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n246), .A3(new_n254), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n211), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n210), .B1(new_n205), .B2(new_n206), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n221), .B(new_n203), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n234), .A2(new_n226), .A3(new_n223), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n262), .B1(new_n267), .B2(new_n244), .ZN(new_n268));
  NAND2_X1  g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT64), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n259), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G71gat), .B(G99gat), .Z(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT33), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(KEYINPUT32), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n271), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n270), .B1(new_n259), .B2(new_n268), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT34), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n271), .A2(KEYINPUT32), .ZN(new_n283));
  INV_X1    g082(.A(new_n271), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n283), .B(new_n274), .C1(new_n284), .C2(KEYINPUT33), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n280), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G228gat), .A2(G233gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT2), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT75), .B(G155gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(G162gat), .ZN(new_n290));
  INV_X1    g089(.A(G141gat), .ZN(new_n291));
  INV_X1    g090(.A(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294));
  AND2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT2), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT74), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G155gat), .B2(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI22_X1  g106(.A1(new_n290), .A2(new_n297), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G211gat), .A2(G218gat), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(G197gat), .A2(G204gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(G197gat), .A2(G204gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n309), .B(new_n312), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n309), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(new_n316), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(new_n319), .C1(new_n314), .C2(new_n313), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n308), .B1(new_n321), .B2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n287), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n297), .ZN(new_n325));
  AND2_X1   g124(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n327));
  OAI21_X1  g126(.A(G162gat), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT2), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n293), .A2(new_n288), .A3(new_n294), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n325), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT29), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n320), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n322), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  OAI221_X1 g136(.A(new_n322), .B1(new_n323), .B2(new_n287), .C1(new_n334), .C2(new_n335), .ZN(new_n338));
  AOI21_X1  g137(.A(G22gat), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(G22gat), .A3(new_n338), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT31), .ZN(new_n344));
  INV_X1    g143(.A(G50gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n340), .A2(new_n347), .A3(new_n341), .A4(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n282), .B1(new_n280), .B2(new_n285), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n286), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n297), .B1(KEYINPUT2), .B2(new_n328), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n307), .A2(new_n300), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n331), .A2(new_n306), .A3(new_n303), .A4(new_n305), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n357), .B(new_n333), .C1(new_n290), .C2(new_n297), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n258), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT5), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT4), .B1(new_n258), .B2(new_n308), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n332), .A2(new_n365), .A3(new_n262), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n363), .B2(new_n366), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n359), .B(new_n362), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT5), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n258), .A2(new_n308), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n332), .A2(new_n262), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(new_n361), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n363), .A2(new_n375), .A3(new_n366), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT76), .B(KEYINPUT4), .C1(new_n258), .C2(new_n308), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n377), .A3(new_n360), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n374), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G57gat), .ZN(new_n382));
  INV_X1    g181(.A(G85gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT78), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n379), .ZN(new_n387));
  INV_X1    g186(.A(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n369), .A2(new_n379), .A3(new_n391), .A4(new_n384), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n386), .A2(new_n389), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT83), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n389), .A2(new_n390), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT6), .B1(new_n385), .B2(KEYINPUT78), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n389), .A4(new_n392), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT72), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT29), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n235), .B2(new_n245), .ZN(new_n405));
  INV_X1    g204(.A(new_n402), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n267), .A2(new_n244), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n335), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n235), .A2(new_n245), .A3(new_n402), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n403), .B1(new_n267), .B2(new_n244), .ZN(new_n410));
  INV_X1    g209(.A(new_n335), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G64gat), .ZN(new_n414));
  INV_X1    g213(.A(G92gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n408), .A2(new_n412), .A3(KEYINPUT30), .A4(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n411), .B1(new_n409), .B2(new_n410), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n408), .A2(new_n416), .A3(new_n412), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n417), .B(new_n421), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n353), .A2(new_n400), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n386), .A2(new_n390), .A3(new_n392), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT79), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n397), .A2(new_n432), .A3(new_n392), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n389), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n427), .B1(new_n434), .B2(new_n396), .ZN(new_n435));
  NOR4_X1   g234(.A1(new_n286), .A2(new_n351), .A3(new_n352), .A4(new_n202), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n202), .A2(new_n429), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n389), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n430), .B2(KEYINPUT79), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n395), .B1(new_n439), .B2(new_n433), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n351), .B1(new_n440), .B2(new_n427), .ZN(new_n441));
  INV_X1    g240(.A(new_n351), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n359), .B1(new_n367), .B2(new_n368), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n361), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n371), .A2(new_n372), .A3(new_n360), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT39), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n447), .A3(new_n361), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n384), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(KEYINPUT82), .A2(KEYINPUT40), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n446), .A2(new_n384), .A3(new_n452), .A4(new_n448), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n427), .A2(new_n389), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT37), .B1(new_n419), .B2(new_n420), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n408), .A2(new_n456), .A3(new_n412), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n418), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT38), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n422), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT38), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n457), .A2(new_n463), .A3(new_n418), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n408), .A2(KEYINPUT84), .A3(new_n412), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(KEYINPUT37), .C1(KEYINPUT84), .C2(new_n408), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(KEYINPUT85), .A3(KEYINPUT38), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n442), .B(new_n454), .C1(new_n400), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n286), .A2(new_n352), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n286), .B2(new_n352), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n441), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n437), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G134gat), .B(G162gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT101), .ZN(new_n479));
  AND2_X1   g278(.A1(G232gat), .A2(G233gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT41), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n479), .B(new_n481), .Z(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT104), .ZN(new_n483));
  INV_X1    g282(.A(G43gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G50gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n345), .A2(G43gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT15), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT14), .ZN(new_n493));
  AND4_X1   g292(.A1(new_n487), .A2(new_n489), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT87), .B1(new_n484), .B2(G50gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n345), .A3(G43gat), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n496), .A2(new_n498), .B1(new_n484), .B2(G50gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT86), .B(KEYINPUT15), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n494), .B(new_n495), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n493), .A2(new_n489), .A3(new_n490), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n487), .C1(new_n499), .C2(new_n500), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n495), .B1(new_n502), .B2(new_n487), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT102), .B1(new_n383), .B2(new_n415), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT102), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(G85gat), .A3(G92gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT7), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT102), .B(new_n511), .C1(new_n383), .C2(new_n415), .ZN(new_n512));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513));
  AOI22_X1  g312(.A1(KEYINPUT8), .A2(new_n513), .B1(new_n383), .B2(new_n415), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(G99gat), .B(G106gat), .Z(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n516), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(new_n510), .A3(new_n512), .A4(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n506), .A2(new_n521), .B1(KEYINPUT41), .B2(new_n480), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT17), .B1(new_n501), .B2(new_n505), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT89), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT92), .B1(new_n506), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n501), .A2(new_n505), .A3(new_n527), .A4(KEYINPUT17), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n521), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n524), .A2(new_n529), .A3(KEYINPUT103), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT103), .B1(new_n524), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n522), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G190gat), .B(G218gat), .Z(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n524), .A2(new_n529), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT103), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n524), .A2(new_n529), .A3(KEYINPUT103), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n535), .B1(new_n540), .B2(new_n522), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n483), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n532), .A2(new_n533), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n522), .A3(new_n535), .ZN(new_n544));
  INV_X1    g343(.A(new_n482), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(KEYINPUT104), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G15gat), .B(G22gat), .Z(new_n549));
  INV_X1    g348(.A(G1gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT16), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(G1gat), .ZN(new_n554));
  INV_X1    g353(.A(G8gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT91), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n551), .B(new_n554), .C1(KEYINPUT90), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G8gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(KEYINPUT90), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n556), .B1(new_n549), .B2(new_n550), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n552), .B(new_n562), .C1(new_n553), .C2(G1gat), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G71gat), .B(G78gat), .Z(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n558), .B(new_n564), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT100), .Z(new_n574));
  INV_X1    g373(.A(new_n571), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT98), .B1(new_n575), .B2(KEYINPUT21), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n577), .A3(new_n572), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT99), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n576), .A2(new_n583), .A3(new_n578), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n580), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n574), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n581), .ZN(new_n590));
  INV_X1    g389(.A(new_n574), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n591), .A3(new_n585), .ZN(new_n592));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n588), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n588), .B2(new_n592), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n548), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n558), .A2(new_n564), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n526), .B2(new_n528), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n524), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n506), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n558), .A2(new_n501), .A3(new_n564), .A4(new_n505), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n606), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n605), .B(KEYINPUT13), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n602), .A2(new_n506), .A3(KEYINPUT94), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n606), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n610), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G113gat), .B(G141gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT11), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G169gat), .ZN(new_n623));
  INV_X1    g422(.A(G197gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(KEYINPUT96), .A3(new_n626), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n524), .A2(new_n603), .B1(new_n602), .B2(new_n506), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n608), .B1(new_n631), .B2(new_n605), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n626), .B1(new_n632), .B2(KEYINPUT97), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT97), .B1(new_n607), .B2(new_n609), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n613), .A2(new_n615), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n617), .A3(new_n614), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n616), .A2(KEYINPUT95), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n629), .A2(new_n630), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n225), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G204gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n571), .A2(new_n520), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n569), .A2(new_n517), .A3(new_n570), .A4(new_n519), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT10), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT106), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n648), .B2(new_n650), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n645), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n655), .B1(new_n660), .B2(new_n649), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n644), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n661), .B(KEYINPUT105), .Z(new_n664));
  NOR2_X1   g463(.A1(new_n656), .A2(new_n644), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n601), .A2(new_n640), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n477), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n440), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g470(.A1(new_n669), .A2(new_n427), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n555), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n553), .A2(new_n555), .ZN(new_n675));
  NAND2_X1  g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n669), .A2(new_n680), .A3(new_n471), .ZN(new_n681));
  INV_X1    g480(.A(new_n475), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n669), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n683), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n351), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  AOI21_X1  g486(.A(new_n548), .B1(new_n437), .B2(new_n476), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n640), .A2(new_n600), .A3(new_n667), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n491), .A3(new_n440), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(new_n689), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n695));
  INV_X1    g494(.A(new_n483), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n543), .B2(new_n544), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n441), .A2(new_n470), .A3(new_n475), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n429), .A2(new_n202), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n435), .A2(new_n436), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT44), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n694), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n440), .ZN(new_n709));
  OAI21_X1  g508(.A(G29gat), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n710), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n690), .A2(G36gat), .A3(new_n428), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n708), .B2(new_n428), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(new_n471), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n690), .A2(G43gat), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n682), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(G43gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n719), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n719), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n724), .ZN(G1330gat));
  NOR2_X1   g524(.A1(new_n442), .A2(G50gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n690), .A2(new_n727), .B1(KEYINPUT108), .B2(KEYINPUT48), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n688), .A2(new_n705), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT44), .B(new_n548), .C1(new_n437), .C2(new_n476), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n351), .B(new_n689), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT109), .B(new_n728), .C1(new_n731), .C2(G50gat), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(G50gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n728), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n732), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n735), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n737), .A2(new_n738), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n734), .A2(new_n733), .A3(new_n735), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n739), .A2(new_n744), .ZN(G1331gat));
  NAND2_X1  g544(.A1(new_n639), .A2(new_n633), .ZN(new_n746));
  INV_X1    g545(.A(new_n630), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT96), .B1(new_n620), .B2(new_n626), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n601), .A2(new_n749), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n477), .A2(new_n667), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n440), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g552(.A(new_n428), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n755), .B(new_n756), .Z(G1333gat));
  INV_X1    g556(.A(G71gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n751), .A2(new_n758), .A3(new_n471), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n751), .A2(new_n682), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n758), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT110), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n763), .B(new_n759), .C1(new_n760), .C2(new_n758), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n762), .A2(KEYINPUT50), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT50), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n351), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  INV_X1    g568(.A(new_n667), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n749), .A2(new_n600), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n688), .B2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n774), .B(new_n548), .C1(new_n437), .C2(new_n476), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n703), .A2(new_n774), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n688), .A2(KEYINPUT111), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n777), .A2(KEYINPUT51), .A3(new_n772), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n770), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n383), .A3(new_n440), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n704), .A2(new_n706), .ZN(new_n782));
  INV_X1    g581(.A(new_n772), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n770), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n440), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n383), .B2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n776), .A2(new_n779), .A3(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT112), .B(new_n771), .C1(new_n773), .C2(new_n775), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n770), .A2(G92gat), .A3(new_n428), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n782), .A2(new_n427), .A3(new_n784), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G92gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n783), .B1(new_n703), .B2(new_n774), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n797), .B2(new_n778), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n773), .A2(new_n771), .A3(new_n775), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n791), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(new_n802), .ZN(G1337gat));
  AOI21_X1  g602(.A(G99gat), .B1(new_n780), .B2(new_n471), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n782), .A2(G99gat), .A3(new_n682), .A4(new_n784), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT114), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n716), .B(new_n770), .C1(new_n776), .C2(new_n779), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n808), .B(new_n805), .C1(new_n809), .C2(G99gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1338gat));
  NOR3_X1   g610(.A1(new_n770), .A2(G106gat), .A3(new_n442), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n789), .A2(new_n790), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n782), .A2(new_n351), .A3(new_n784), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n812), .B1(new_n798), .B2(new_n799), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n812), .C1(new_n798), .C2(new_n799), .ZN(new_n821));
  XNOR2_X1  g620(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n819), .A2(new_n815), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n817), .A2(new_n823), .ZN(G1339gat));
  OAI22_X1  g623(.A1(new_n631), .A2(new_n605), .B1(new_n614), .B2(new_n635), .ZN(new_n825));
  INV_X1    g624(.A(new_n625), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n746), .A2(new_n667), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n651), .B2(new_n652), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n648), .A2(new_n650), .A3(KEYINPUT117), .A4(new_n655), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n656), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n654), .A2(new_n833), .A3(new_n658), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n644), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(new_n838), .B1(new_n664), .B2(new_n665), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT55), .A4(new_n644), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n548), .B(new_n828), .C1(new_n640), .C2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n746), .A2(new_n839), .A3(new_n840), .A4(new_n827), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n600), .B1(new_n843), .B2(new_n698), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n842), .A2(new_n844), .B1(new_n750), .B2(new_n770), .ZN(new_n845));
  INV_X1    g644(.A(new_n353), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n709), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n428), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n640), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n640), .A2(G113gat), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT118), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1340gat));
  INV_X1    g653(.A(new_n848), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n667), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n600), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(G127gat), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n698), .A2(new_n428), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT120), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT56), .Z(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n848), .B2(new_n548), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1343gat));
  NOR2_X1   g666(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n868));
  AND2_X1   g667(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT57), .B1(new_n845), .B2(new_n442), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n629), .A2(new_n630), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n841), .B1(new_n871), .B2(new_n746), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n828), .A2(new_n548), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n844), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n750), .A2(new_n770), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n351), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n709), .A2(new_n427), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n870), .A2(new_n878), .A3(new_n475), .A4(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n640), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n475), .A2(new_n351), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT121), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n876), .A2(new_n440), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n291), .A3(new_n428), .A4(new_n749), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n868), .B(new_n869), .C1(new_n881), .C2(new_n885), .ZN(new_n886));
  AND4_X1   g685(.A1(KEYINPUT122), .A2(new_n881), .A3(KEYINPUT58), .A4(new_n885), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(G1344gat));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n880), .A2(new_n770), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n889), .B(G148gat), .C1(new_n880), .C2(new_n770), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n884), .A2(new_n428), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n667), .A2(new_n292), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n891), .A2(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1345gat));
  INV_X1    g695(.A(new_n600), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n600), .A2(new_n289), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT123), .Z(new_n900));
  OAI22_X1  g699(.A1(new_n898), .A2(new_n289), .B1(new_n880), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n880), .B2(new_n548), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n884), .A2(new_n302), .A3(new_n863), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n440), .A2(new_n428), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n471), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT124), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n876), .A2(new_n908), .A3(new_n442), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n640), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n845), .A2(new_n440), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n427), .A3(new_n353), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n749), .A2(new_n224), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1348gat));
  OAI21_X1  g713(.A(G176gat), .B1(new_n909), .B2(new_n770), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n667), .A2(new_n225), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n912), .B2(new_n916), .ZN(G1349gat));
  OAI21_X1  g716(.A(G183gat), .B1(new_n909), .B2(new_n897), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n600), .A2(new_n205), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n920), .B(new_n921), .Z(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n909), .B2(new_n548), .ZN(new_n923));
  NOR2_X1   g722(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n698), .A2(new_n206), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n927));
  OAI221_X1 g726(.A(new_n925), .B1(new_n912), .B2(new_n926), .C1(new_n923), .C2(new_n927), .ZN(G1351gat));
  AND2_X1   g727(.A1(new_n870), .A2(new_n475), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n878), .A3(new_n906), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n624), .A3(new_n640), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n882), .A2(new_n428), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n911), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n749), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n931), .A2(new_n935), .ZN(G1352gat));
  NOR3_X1   g735(.A1(new_n933), .A2(G204gat), .A3(new_n770), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT62), .ZN(new_n938));
  OAI21_X1  g737(.A(G204gat), .B1(new_n930), .B2(new_n770), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n310), .A3(new_n600), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n929), .A2(new_n600), .A3(new_n878), .A4(new_n906), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(G1354gat));
  OAI21_X1  g745(.A(new_n311), .B1(new_n933), .B2(new_n548), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n930), .A2(new_n311), .A3(new_n548), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(G1355gat));
endmodule


