//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT64), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(new_n192), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n193), .A2(new_n197), .B1(new_n191), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(KEYINPUT67), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n188), .A2(new_n205), .A3(KEYINPUT1), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n194), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  AND4_X1   g022(.A1(new_n208), .A2(new_n188), .A3(new_n190), .A4(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n201), .B1(G125), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT88), .B(G224), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G953), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI221_X1 g028(.A(new_n201), .B1(G953), .B2(new_n212), .C1(G125), .C2(new_n210), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT81), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n217), .A2(new_n224), .A3(new_n218), .A4(G104), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(new_n221), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n222), .B2(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n218), .A2(KEYINPUT82), .A3(G104), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n223), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT84), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT68), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n240), .A3(G119), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n241), .A2(KEYINPUT69), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT69), .B1(new_n241), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT5), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(G113), .B1(new_n243), .B2(KEYINPUT5), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n243), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n236), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n241), .A2(KEYINPUT69), .A3(new_n243), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n251), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n253), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n225), .A2(new_n223), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n222), .A2(G107), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n224), .B1(new_n262), .B2(new_n217), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n260), .B(G101), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(G101), .B1(new_n261), .B2(new_n263), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n254), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT87), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n254), .A2(KEYINPUT87), .A3(new_n267), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G122), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n270), .A2(new_n271), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n254), .A2(KEYINPUT87), .A3(new_n267), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT87), .B1(new_n254), .B2(new_n267), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(new_n273), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n266), .A2(new_n264), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n252), .B1(new_n246), .B2(new_n248), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n259), .B1(new_n280), .B2(new_n236), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n273), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT6), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n216), .B(new_n275), .C1(new_n278), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT89), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n274), .B1(new_n281), .B2(KEYINPUT87), .ZN(new_n286));
  OAI211_X1 g100(.A(KEYINPUT6), .B(new_n282), .C1(new_n286), .C2(new_n276), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n216), .A4(new_n275), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n232), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n241), .A2(KEYINPUT5), .A3(new_n243), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n252), .B1(new_n293), .B2(new_n248), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n236), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n273), .B(KEYINPUT8), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n282), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n214), .B(new_n215), .C1(KEYINPUT7), .C2(new_n213), .ZN(new_n299));
  OR3_X1    g113(.A1(new_n211), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n290), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n285), .A2(new_n289), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT90), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n302), .B1(new_n284), .B2(KEYINPUT89), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n289), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n306), .A3(new_n289), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT31), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n316));
  XNOR2_X1  g130(.A(G134), .B(G137), .ZN(new_n317));
  INV_X1    g131(.A(G131), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G134), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G137), .ZN(new_n321));
  INV_X1    g135(.A(G137), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G134), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT66), .B(G131), .C1(new_n321), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n320), .B2(G137), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n322), .A2(KEYINPUT11), .A3(G134), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(G131), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n325), .B(new_n331), .C1(new_n207), .C2(new_n209), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n318), .A2(KEYINPUT65), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n333), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n335), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n193), .A2(new_n197), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n199), .A2(new_n191), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n332), .A2(new_n340), .A3(new_n258), .A4(new_n253), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n332), .A2(KEYINPUT30), .A3(new_n340), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT30), .B1(new_n332), .B2(new_n340), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n345), .B2(new_n259), .ZN(new_n346));
  INV_X1    g160(.A(G237), .ZN(new_n347));
  INV_X1    g161(.A(G953), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(G210), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT26), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(new_n221), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n315), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n332), .A2(new_n340), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n332), .A2(new_n340), .A3(KEYINPUT30), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n259), .A3(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(new_n315), .A3(new_n353), .A4(new_n341), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n341), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n244), .A2(new_n245), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n252), .B1(new_n363), .B2(new_n251), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(KEYINPUT28), .A3(new_n340), .A4(new_n332), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n355), .A2(new_n259), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n352), .B(G101), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n360), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n314), .B1(new_n354), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT70), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT32), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n359), .A2(new_n341), .A3(new_n353), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT31), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n360), .A3(new_n369), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT70), .A3(new_n314), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(KEYINPUT32), .A3(new_n314), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n353), .B1(new_n367), .B2(KEYINPUT29), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n366), .A2(KEYINPUT71), .A3(new_n341), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT71), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n355), .A2(new_n383), .A3(new_n259), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(KEYINPUT28), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n341), .A2(KEYINPUT72), .A3(new_n361), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT72), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n362), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n381), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n346), .A2(new_n368), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n290), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n392));
  OAI21_X1  g206(.A(G472), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n379), .A2(new_n380), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n242), .B2(G128), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n202), .A2(KEYINPUT74), .A3(G119), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT73), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT23), .A2(G119), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(G128), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n202), .A2(KEYINPUT73), .A3(KEYINPUT23), .A4(G119), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G110), .ZN(new_n406));
  XOR2_X1   g220(.A(G119), .B(G128), .Z(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT24), .B(G110), .ZN(new_n408));
  INV_X1    g222(.A(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G125), .ZN(new_n410));
  INV_X1    g224(.A(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G140), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n412), .A3(KEYINPUT16), .ZN(new_n413));
  OR3_X1    g227(.A1(new_n411), .A2(KEYINPUT16), .A3(G140), .ZN(new_n414));
  AOI21_X1  g228(.A(G146), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(G146), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI221_X1 g231(.A(new_n406), .B1(new_n407), .B2(new_n408), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n407), .A2(new_n408), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n405), .B2(G110), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(new_n412), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT75), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G125), .B(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT75), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n425), .A3(new_n187), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n416), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n348), .A2(G221), .A3(G234), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT22), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(G137), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n418), .A2(new_n427), .A3(new_n431), .ZN(new_n434));
  INV_X1    g248(.A(G217), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(G234), .B2(new_n290), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G902), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n437), .B(KEYINPUT77), .Z(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT78), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n290), .A3(new_n434), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT76), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT25), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT25), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(KEYINPUT76), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n441), .B1(new_n447), .B2(new_n436), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n394), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  OAI21_X1  g265(.A(G221), .B1(new_n451), .B2(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT79), .ZN(new_n453));
  INV_X1    g267(.A(G469), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(G128), .A3(new_n206), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n191), .ZN(new_n457));
  INV_X1    g271(.A(new_n209), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n226), .A2(new_n231), .A3(new_n234), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n234), .B1(new_n226), .B2(new_n231), .ZN(new_n461));
  OAI211_X1 g275(.A(KEYINPUT10), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n337), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT10), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n203), .A2(KEYINPUT83), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n188), .A2(new_n466), .A3(KEYINPUT1), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(G128), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n209), .B1(new_n468), .B2(new_n191), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n464), .B1(new_n469), .B2(new_n232), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n266), .A2(new_n200), .A3(new_n264), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n462), .A2(new_n463), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n348), .A2(G227), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(G140), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT80), .B(G110), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n474), .B(new_n475), .Z(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n233), .A2(new_n210), .A3(new_n235), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n469), .A2(new_n232), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT12), .B1(new_n337), .B2(KEYINPUT85), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n337), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n469), .A2(new_n232), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n460), .A2(new_n461), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(new_n210), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n481), .B1(new_n486), .B2(new_n463), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n477), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n471), .A2(new_n470), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT10), .B1(new_n207), .B2(new_n209), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n233), .B2(new_n235), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n337), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n476), .B1(new_n492), .B2(new_n472), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n454), .B(new_n290), .C1(new_n488), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n482), .B1(new_n480), .B2(new_n337), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n463), .B(new_n481), .C1(new_n478), .C2(new_n479), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n472), .B(new_n476), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n472), .ZN(new_n500));
  INV_X1    g314(.A(new_n476), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n503), .A2(KEYINPUT86), .A3(new_n454), .A4(new_n290), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n487), .A2(new_n483), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n476), .B1(new_n506), .B2(new_n472), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n492), .A2(new_n472), .A3(new_n476), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n290), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G469), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n453), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(G475), .A2(G902), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n417), .B2(new_n415), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n413), .A2(new_n414), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n187), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT91), .A3(new_n416), .ZN(new_n517));
  NOR2_X1   g331(.A1(G237), .A2(G953), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(G143), .A3(G214), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(G143), .B1(new_n518), .B2(G214), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n189), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n318), .A3(new_n519), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(KEYINPUT17), .B(G131), .C1(new_n520), .C2(new_n521), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n514), .A2(new_n517), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G113), .B(G122), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n222), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n426), .B1(new_n187), .B2(new_n424), .ZN(new_n532));
  NAND2_X1  g346(.A1(KEYINPUT18), .A2(G131), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n525), .A2(new_n519), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n525), .B2(new_n519), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n529), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT19), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n423), .A2(new_n425), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n421), .A2(KEYINPUT19), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n187), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n522), .A2(new_n526), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n416), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n531), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n512), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT20), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n537), .ZN(new_n548));
  INV_X1    g362(.A(new_n531), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n529), .A2(new_n531), .A3(new_n537), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n512), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n531), .B1(new_n529), .B2(new_n537), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n290), .B1(new_n538), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n202), .A2(G143), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n320), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n189), .A2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n202), .A2(G143), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT13), .ZN(new_n565));
  XNOR2_X1  g379(.A(G128), .B(G143), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n562), .A2(new_n565), .B1(new_n320), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n238), .A2(new_n240), .A3(G122), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n237), .A2(G122), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n568), .A2(new_n218), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n218), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n451), .A2(new_n435), .A3(G953), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n563), .A2(new_n564), .A3(new_n320), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n320), .B1(new_n563), .B2(new_n564), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n563), .A2(new_n564), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G134), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n563), .A2(new_n564), .A3(new_n320), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(KEYINPUT92), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n568), .A2(new_n218), .A3(new_n569), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT14), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n568), .A2(new_n584), .A3(new_n569), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT14), .A4(G122), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n585), .A2(G107), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n572), .B(new_n573), .C1(new_n583), .C2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(G107), .A3(new_n586), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n590), .A2(new_n582), .A3(new_n581), .A4(new_n577), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n573), .B1(new_n591), .B2(new_n572), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n290), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT15), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI221_X1 g410(.A(new_n290), .B1(KEYINPUT15), .B2(new_n594), .C1(new_n589), .C2(new_n592), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(G234), .A2(G237), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n599), .A2(G952), .A3(new_n348), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(G902), .A3(G953), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT93), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT21), .B(G898), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n559), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n511), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n313), .A2(new_n449), .A3(new_n450), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  INV_X1    g422(.A(new_n450), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n591), .A2(new_n572), .ZN(new_n611));
  INV_X1    g425(.A(new_n573), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n613), .B2(new_n588), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n610), .B1(new_n614), .B2(G478), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n593), .A2(KEYINPUT94), .A3(new_n594), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n589), .B2(new_n592), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n613), .A2(KEYINPUT33), .A3(new_n588), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n620), .A3(G478), .A4(new_n290), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n555), .A2(new_n558), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n604), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n304), .A2(new_n307), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n609), .B(new_n624), .C1(new_n625), .C2(new_n312), .ZN(new_n626));
  INV_X1    g440(.A(new_n511), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n377), .A2(new_n290), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n448), .A3(new_n373), .A4(new_n378), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  AND3_X1   g448(.A1(new_n308), .A2(new_n306), .A3(new_n289), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n306), .B1(new_n308), .B2(new_n289), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n450), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n555), .A2(KEYINPUT95), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT95), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n547), .A2(new_n554), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n638), .A2(new_n558), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n641), .A2(new_n642), .A3(new_n598), .A4(new_n623), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n638), .A2(new_n558), .A3(new_n598), .A4(new_n640), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT96), .B1(new_n644), .B2(new_n604), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n631), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NAND3_X1  g464(.A1(new_n629), .A2(new_n373), .A3(new_n378), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n432), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n428), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n447), .A2(new_n436), .B1(new_n439), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n313), .A2(new_n450), .A3(new_n606), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AOI211_X1 g473(.A(new_n609), .B(new_n654), .C1(new_n625), .C2(new_n312), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n394), .A2(new_n511), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n600), .B1(new_n602), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n644), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XOR2_X1   g480(.A(new_n313), .B(KEYINPUT38), .Z(new_n667));
  XOR2_X1   g481(.A(new_n663), .B(KEYINPUT39), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n627), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT40), .Z(new_n671));
  INV_X1    g485(.A(new_n346), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n353), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n382), .A2(new_n384), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n673), .B(new_n290), .C1(new_n353), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G472), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n379), .A2(new_n380), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n379), .A2(KEYINPUT98), .A3(new_n380), .A4(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n654), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n559), .A2(new_n598), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n683), .A3(new_n609), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  OR3_X1    g499(.A1(new_n667), .A2(new_n671), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  INV_X1    g501(.A(new_n663), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n622), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n660), .A2(new_n661), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT99), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n187), .ZN(G48));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n454), .B1(new_n503), .B2(new_n290), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n496), .B2(new_n504), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(KEYINPUT100), .A3(new_n452), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT100), .B1(new_n696), .B2(new_n452), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n694), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n695), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n505), .A2(new_n452), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT100), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n696), .A2(KEYINPUT100), .A3(new_n452), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(KEYINPUT101), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n699), .A2(new_n626), .A3(new_n705), .A4(new_n449), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT41), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G113), .ZN(G15));
  NAND4_X1  g522(.A1(new_n647), .A2(new_n699), .A3(new_n449), .A4(new_n705), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NOR2_X1   g524(.A1(new_n697), .A2(new_n698), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n660), .A2(new_n711), .A3(new_n394), .A4(new_n605), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  AOI211_X1 g527(.A(new_n609), .B(new_n683), .C1(new_n625), .C2(new_n312), .ZN(new_n714));
  INV_X1    g528(.A(new_n314), .ZN(new_n715));
  INV_X1    g529(.A(new_n360), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n389), .A2(new_n368), .B1(KEYINPUT31), .B2(new_n375), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n716), .B1(new_n717), .B2(KEYINPUT102), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n389), .A2(new_n368), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n719), .B1(new_n720), .B2(new_n354), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n715), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n448), .ZN(new_n723));
  INV_X1    g537(.A(new_n629), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n604), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n699), .A2(new_n714), .A3(new_n705), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NOR2_X1   g541(.A1(new_n722), .A2(new_n724), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n660), .A2(new_n711), .A3(new_n690), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n312), .A2(new_n450), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n311), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n311), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n452), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n507), .A2(new_n508), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n740), .B1(new_n741), .B2(G469), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n738), .B1(new_n505), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n505), .A2(new_n738), .A3(new_n742), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n734), .A2(new_n449), .A3(new_n736), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n731), .B1(new_n747), .B2(new_n689), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n749));
  INV_X1    g563(.A(new_n380), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT32), .B1(new_n377), .B2(new_n314), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n371), .A2(new_n374), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(KEYINPUT106), .A3(new_n380), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n393), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n689), .A2(new_n731), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n755), .A2(new_n448), .A3(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n734), .A2(new_n757), .A3(new_n736), .A4(new_n746), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n748), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  INV_X1    g577(.A(new_n664), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n747), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n320), .ZN(G36));
  OR2_X1    g580(.A1(new_n507), .A2(new_n508), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n454), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n770));
  OAI22_X1  g584(.A1(new_n769), .A2(new_n770), .B1(new_n768), .B2(new_n767), .ZN(new_n771));
  AOI211_X1 g585(.A(KEYINPUT108), .B(new_n454), .C1(new_n767), .C2(new_n768), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n740), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n505), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n452), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n669), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n311), .A2(new_n732), .A3(new_n735), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n735), .B1(new_n311), .B2(new_n732), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n617), .A2(new_n621), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n558), .A3(new_n555), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT109), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT43), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n651), .A3(new_n682), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT110), .Z(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT111), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n778), .A2(new_n781), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  XNOR2_X1  g607(.A(new_n777), .B(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n734), .A2(new_n736), .ZN(new_n795));
  OR4_X1    g609(.A1(new_n394), .A2(new_n795), .A3(new_n448), .A4(new_n689), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  INV_X1    g612(.A(new_n711), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n681), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n448), .A3(new_n600), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT115), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n622), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n799), .A2(new_n637), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n785), .A2(new_n600), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n448), .A3(new_n728), .ZN(new_n807));
  OAI211_X1 g621(.A(G952), .B(new_n348), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n800), .A2(new_n806), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n448), .A3(new_n755), .ZN(new_n810));
  AND2_X1   g624(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n804), .B(new_n812), .C1(new_n810), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n696), .A2(new_n453), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n794), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n807), .A2(new_n795), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n559), .A2(new_n782), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n803), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n807), .A2(new_n450), .A3(new_n799), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n667), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(KEYINPUT50), .A3(new_n667), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n722), .A2(new_n724), .A3(new_n654), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n825), .A2(new_n826), .B1(new_n809), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n814), .B1(new_n819), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n821), .A2(new_n833), .A3(new_n828), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n817), .A2(new_n818), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n815), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT117), .B1(new_n836), .B2(new_n815), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n709), .A2(new_n706), .A3(new_n726), .A4(new_n712), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n496), .A2(new_n504), .B1(new_n509), .B2(G469), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n553), .B1(new_n552), .B2(new_n512), .ZN(new_n842));
  INV_X1    g656(.A(new_n512), .ZN(new_n843));
  AOI211_X1 g657(.A(KEYINPUT20), .B(new_n843), .C1(new_n550), .C2(new_n551), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n598), .B(new_n558), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n623), .B1(new_n622), .B2(new_n846), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n630), .A2(new_n841), .A3(new_n847), .A4(new_n453), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n313), .A2(new_n848), .A3(new_n450), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n607), .A2(new_n656), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n607), .A2(new_n656), .A3(new_n849), .A4(KEYINPUT112), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n840), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n682), .A2(new_n663), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n681), .A2(new_n746), .A3(new_n714), .A4(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n660), .B(new_n661), .C1(new_n664), .C2(new_n690), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n729), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n856), .A2(new_n857), .A3(new_n729), .A4(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n747), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n779), .A2(new_n780), .A3(new_n654), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n598), .A2(new_n663), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n394), .A2(new_n511), .A3(new_n641), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n745), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n452), .B1(new_n867), .B2(new_n743), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n728), .A2(new_n690), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n863), .A2(new_n664), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n762), .A2(new_n854), .A3(new_n862), .A4(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n874), .A2(KEYINPUT114), .B1(new_n875), .B2(new_n872), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(KEYINPUT114), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n870), .A2(new_n682), .A3(new_n736), .A4(new_n734), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n764), .B2(new_n747), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n781), .A2(KEYINPUT107), .A3(new_n746), .A4(new_n757), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n758), .A2(new_n759), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n748), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .A3(new_n854), .A4(new_n862), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n878), .B1(KEYINPUT54), .B2(new_n887), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n839), .A2(new_n888), .B1(G952), .B2(G953), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n723), .A2(new_n783), .A3(new_n609), .A4(new_n453), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT49), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n696), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n891), .B2(new_n696), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n667), .A2(new_n801), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n889), .A2(new_n894), .ZN(G75));
  AND2_X1   g709(.A1(new_n879), .A2(new_n886), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n290), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(G210), .ZN(new_n898));
  NOR2_X1   g712(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT55), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n287), .A2(new_n275), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n216), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT55), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n898), .A2(new_n904), .A3(new_n899), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n901), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n348), .A2(G952), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  XNOR2_X1  g723(.A(new_n887), .B(KEYINPUT54), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n740), .B(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n503), .B(KEYINPUT120), .Z(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n897), .A2(new_n773), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n908), .B1(new_n914), .B2(new_n915), .ZN(G54));
  INV_X1    g730(.A(new_n908), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n552), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n552), .B2(new_n918), .ZN(G60));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT59), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n619), .A2(new_n910), .A3(new_n620), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n888), .A2(new_n922), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n619), .A2(new_n620), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n908), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(G63));
  XNOR2_X1  g740(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT122), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n435), .A2(new_n290), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(new_n930));
  AOI21_X1  g744(.A(KEYINPUT123), .B1(new_n887), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n932));
  INV_X1    g746(.A(new_n930), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n932), .B(new_n933), .C1(new_n879), .C2(new_n886), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n653), .ZN(new_n936));
  OAI211_X1 g750(.A(KEYINPUT61), .B(new_n917), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n433), .A2(new_n434), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n939), .ZN(new_n941));
  NOR4_X1   g755(.A1(new_n931), .A2(new_n934), .A3(KEYINPUT124), .A4(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n937), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n932), .B1(new_n896), .B2(new_n933), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n887), .A2(KEYINPUT123), .A3(new_n930), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n908), .B1(new_n946), .B2(new_n653), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n939), .A3(new_n945), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT61), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT125), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n948), .B(new_n917), .C1(new_n936), .C2(new_n935), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n948), .B(KEYINPUT124), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n953), .B(new_n954), .C1(new_n955), .C2(new_n937), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n950), .A2(new_n956), .ZN(G66));
  XOR2_X1   g771(.A(new_n854), .B(KEYINPUT126), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n348), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n212), .B2(new_n603), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n902), .B1(G898), .B2(new_n348), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n540), .A2(new_n541), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n345), .B(new_n964), .Z(new_n965));
  AND2_X1   g779(.A1(new_n797), .A2(new_n792), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n686), .A2(new_n729), .A3(new_n857), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n622), .A2(new_n846), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n781), .A2(new_n449), .A3(new_n670), .A4(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n966), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n965), .B1(new_n973), .B2(new_n348), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n857), .A2(new_n729), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n714), .A2(new_n448), .A3(new_n755), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n765), .B(new_n975), .C1(new_n778), .C2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n966), .A2(new_n762), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n978), .A2(G953), .ZN(new_n979));
  INV_X1    g793(.A(new_n965), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(G900), .B2(G953), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n974), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n348), .B1(G227), .B2(G900), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n978), .B2(new_n958), .ZN(new_n987));
  INV_X1    g801(.A(new_n391), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n908), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n990));
  INV_X1    g804(.A(new_n673), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n988), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n353), .A2(new_n990), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n672), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n877), .A2(new_n992), .A3(new_n986), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n986), .B1(new_n973), .B2(new_n958), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n991), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n989), .A2(new_n995), .A3(new_n997), .ZN(G57));
endmodule


