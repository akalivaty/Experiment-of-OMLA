//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(new_n461), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n470), .B2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n471), .A2(new_n472), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n481), .B2(new_n461), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n464), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n480), .B(new_n484), .C1(G124), .C2(new_n489), .ZN(G162));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT69), .A2(G114), .ZN(new_n493));
  OAI211_X1 g068(.A(G2104), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n464), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n501), .C1(new_n472), .C2(new_n471), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G651), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n512), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n511), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n507), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n514), .A2(new_n521), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT71), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n518), .A2(new_n528), .A3(G63), .A4(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n527), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n520), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n513), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n520), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n513), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n507), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(new_n520), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n513), .A2(G43), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n507), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(new_n511), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n512), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT73), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(KEYINPUT73), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n555), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n518), .A2(G65), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n560), .B(new_n563), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n555), .A2(G91), .A3(new_n518), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n520), .A2(KEYINPUT74), .A3(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT76), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  NOR3_X1   g154(.A1(new_n578), .A2(new_n570), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n542), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT77), .A4(new_n541), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G301));
  NAND2_X1  g161(.A1(new_n536), .A2(KEYINPUT78), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G286));
  NAND4_X1  g166(.A1(new_n509), .A2(G49), .A3(G543), .A4(new_n510), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n509), .A2(G87), .A3(new_n510), .A4(new_n518), .ZN(new_n593));
  INV_X1    g168(.A(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n516), .A2(new_n594), .A3(new_n517), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n595), .A2(KEYINPUT79), .A3(G651), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT79), .B1(new_n595), .B2(G651), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n592), .B(new_n593), .C1(new_n597), .C2(new_n598), .ZN(G288));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n516), .B2(new_n517), .ZN(new_n601));
  AND2_X1   g176(.A1(G73), .A2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n509), .A2(G48), .A3(G543), .A4(new_n510), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n509), .A2(G86), .A3(new_n510), .A4(new_n518), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n520), .A2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n513), .A2(G47), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n607), .B(new_n608), .C1(new_n507), .C2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(new_n513), .A2(G54), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(new_n507), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n520), .A2(G92), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n585), .ZN(G284));
  AOI21_X1  g197(.A(new_n621), .B1(G868), .B2(new_n585), .ZN(G321));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NOR2_X1   g199(.A1(G286), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n624), .ZN(G297));
  AOI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(new_n624), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n619), .B1(new_n629), .B2(G860), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT80), .Z(G148));
  OAI21_X1  g206(.A(KEYINPUT81), .B1(new_n548), .B2(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n619), .A2(new_n629), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  MUX2_X1   g209(.A(KEYINPUT81), .B(new_n632), .S(new_n634), .Z(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n464), .A2(new_n462), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n482), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n461), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G123), .ZN(new_n644));
  OAI221_X1 g219(.A(new_n641), .B1(new_n642), .B2(new_n643), .C1(new_n488), .C2(new_n644), .ZN(new_n645));
  AOI22_X1  g220(.A1(new_n640), .A2(G2100), .B1(G2096), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n646), .B(new_n647), .C1(G2100), .C2(new_n640), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XOR2_X1   g224(.A(KEYINPUT83), .B(G2438), .Z(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT14), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT84), .Z(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n652), .B2(new_n651), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n661), .A2(new_n665), .A3(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  NOR2_X1   g248(.A1(G2072), .A2(G2078), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n442), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n671), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(KEYINPUT17), .Z(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(new_n673), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n673), .A3(new_n671), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n671), .A3(new_n672), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT18), .Z(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2100), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT89), .B(G2096), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(new_n693), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT20), .Z(new_n697));
  AOI211_X1 g272(.A(new_n695), .B(new_n697), .C1(new_n690), .C2(new_n694), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT32), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1981), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(new_n711), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n706), .A2(G23), .ZN(new_n717));
  INV_X1    g292(.A(G288), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n706), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT33), .B(G1976), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n712), .A2(new_n715), .A3(new_n716), .A4(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n706), .B1(G290), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(G290), .ZN(new_n727));
  INV_X1    g302(.A(G24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(G16), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(G1986), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(G1986), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT90), .B(G29), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(G107), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G2105), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n482), .A2(G131), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n737), .B(new_n739), .C1(G119), .C2(new_n489), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n733), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT35), .B(G1991), .Z(new_n742));
  XOR2_X1   g317(.A(new_n741), .B(new_n742), .Z(new_n743));
  NOR3_X1   g318(.A1(new_n730), .A2(new_n731), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n723), .A2(new_n724), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(KEYINPUT36), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n723), .A2(new_n747), .A3(new_n724), .A4(new_n744), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G16), .A2(G19), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n548), .B2(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G1341), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n733), .A2(G27), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G164), .B2(new_n733), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G32), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n489), .A2(G129), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT99), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT26), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n462), .A2(G105), .ZN(new_n764));
  INV_X1    g339(.A(G141), .ZN(new_n765));
  OR3_X1    g340(.A1(new_n465), .A2(KEYINPUT98), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT98), .B1(new_n465), .B2(new_n765), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n763), .B(new_n764), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n759), .B1(new_n770), .B2(new_n758), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT27), .B(G1996), .Z(new_n772));
  NOR2_X1   g347(.A1(G4), .A2(G16), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n619), .B2(G16), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(G1348), .B2(new_n774), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n757), .B(new_n775), .C1(G1348), .C2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n732), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT93), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G140), .B2(new_n482), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n489), .A2(G128), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n733), .A2(G35), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n733), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2090), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n758), .A2(G33), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(new_n461), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT25), .Z(new_n801));
  AOI211_X1 g376(.A(new_n798), .B(new_n801), .C1(G139), .C2(new_n482), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n758), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2072), .ZN(new_n804));
  NAND2_X1  g379(.A1(G160), .A2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT24), .B(G34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n732), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT97), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G2084), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n751), .A2(G1341), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n795), .A2(new_n804), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n810), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n706), .A2(G5), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G171), .B2(new_n706), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n813), .B1(new_n815), .B2(G1961), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n771), .B2(new_n772), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT101), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n776), .A2(new_n791), .A3(new_n812), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n706), .A2(G21), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G168), .B2(new_n706), .ZN(new_n821));
  INV_X1    g396(.A(G1966), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT30), .B(G28), .ZN(new_n824));
  OR2_X1    g399(.A1(KEYINPUT31), .A2(G11), .ZN(new_n825));
  NAND2_X1  g400(.A1(KEYINPUT31), .A2(G11), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n824), .A2(new_n758), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n645), .B2(new_n732), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n815), .B2(G1961), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT100), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(KEYINPUT101), .B2(new_n817), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n706), .A2(G20), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n626), .B2(new_n706), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1956), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n819), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n749), .A2(new_n838), .ZN(G150));
  XNOR2_X1  g414(.A(G150), .B(KEYINPUT103), .ZN(G311));
  NAND2_X1  g415(.A1(new_n619), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT105), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT104), .B(G55), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n513), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n520), .A2(G93), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n845), .B(new_n846), .C1(new_n507), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n548), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n843), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(G860), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n848), .A2(G860), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT107), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(G145));
  NAND2_X1  g436(.A1(new_n482), .A2(G142), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n461), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  INV_X1    g439(.A(G130), .ZN(new_n865));
  OAI221_X1 g440(.A(new_n862), .B1(new_n863), .B2(new_n864), .C1(new_n488), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n740), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n639), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n494), .A2(new_n495), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n501), .B1(new_n464), .B2(new_n498), .ZN(new_n870));
  INV_X1    g445(.A(new_n502), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT108), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n500), .A2(new_n502), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n869), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n868), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n802), .B(new_n769), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n785), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n878), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(new_n645), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G160), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n883), .B2(new_n881), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g461(.A(G166), .B(G290), .ZN(new_n887));
  XOR2_X1   g462(.A(G288), .B(G305), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT42), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n579), .B1(new_n578), .B2(new_n570), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n560), .A2(new_n563), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n568), .A2(new_n569), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n893), .A2(KEYINPUT76), .A3(new_n576), .A4(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n892), .A2(new_n896), .A3(new_n619), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n619), .B1(new_n892), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n891), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n620), .B1(new_n577), .B2(new_n580), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n896), .A3(new_n619), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(KEYINPUT41), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n849), .B(new_n633), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n897), .A2(new_n898), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n890), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n890), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n848), .A2(new_n624), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(G331));
  NAND3_X1  g490(.A1(new_n587), .A2(G171), .A3(new_n589), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n583), .A2(G168), .A3(new_n584), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n849), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n848), .B(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n916), .A3(new_n917), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n919), .B(new_n922), .C1(new_n897), .C2(new_n898), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT110), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n922), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n904), .A2(new_n907), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n926), .A3(new_n889), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n889), .B1(new_n924), .B2(new_n926), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n933), .B(KEYINPUT43), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  INV_X1    g509(.A(new_n929), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n899), .A2(new_n902), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n925), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n923), .A2(KEYINPUT112), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n923), .A2(KEYINPUT112), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n889), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT113), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n945), .A3(new_n941), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n935), .A2(new_n943), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n932), .A2(new_n934), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n944), .B1(new_n929), .B2(new_n930), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n935), .A2(new_n943), .A3(new_n946), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n944), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(G397));
  INV_X1    g530(.A(new_n598), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n596), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(G1976), .A3(new_n592), .A4(new_n593), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n872), .A2(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n482), .A2(G137), .B1(G101), .B2(new_n462), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT67), .B1(new_n475), .B2(G2105), .ZN(new_n962));
  AOI211_X1 g537(.A(new_n468), .B(new_n461), .C1(new_n473), .C2(new_n474), .ZN(new_n963));
  OAI211_X1 g538(.A(G40), .B(new_n961), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n958), .B(G8), .C1(new_n960), .C2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT52), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n874), .B2(new_n869), .ZN(new_n967));
  NAND3_X1  g542(.A1(G160), .A2(new_n967), .A3(G40), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n968), .A2(new_n970), .A3(G8), .A4(new_n958), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT116), .B(G1981), .Z(new_n974));
  NAND4_X1  g549(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(KEYINPUT117), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(KEYINPUT117), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT49), .B(new_n973), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT118), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n975), .B(KEYINPUT117), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(new_n981), .A3(KEYINPUT49), .A4(new_n973), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n968), .A2(G8), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n973), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT49), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n972), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n964), .B1(new_n989), .B2(new_n960), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n959), .A4(new_n876), .ZN(new_n991));
  AOI21_X1  g566(.A(G1971), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2090), .ZN(new_n993));
  INV_X1    g568(.A(new_n964), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n871), .A2(new_n870), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n996), .B(new_n959), .C1(new_n997), .C2(new_n496), .ZN(new_n998));
  AND4_X1   g573(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(G8), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NOR3_X1   g577(.A1(G166), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n988), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1005), .ZN(new_n1008));
  INV_X1    g583(.A(new_n992), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n995), .A2(KEYINPUT114), .A3(new_n998), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n960), .A2(new_n1011), .A3(KEYINPUT50), .ZN(new_n1012));
  AOI211_X1 g587(.A(G2090), .B(new_n964), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n964), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1016), .A2(new_n1014), .A3(new_n993), .ZN(new_n1017));
  OAI211_X1 g592(.A(G8), .B(new_n1008), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1007), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(new_n810), .A3(new_n994), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n960), .A2(new_n989), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n994), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n822), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1002), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n536), .A2(G8), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT124), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT125), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1028), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT125), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1016), .A2(new_n810), .B1(new_n822), .B2(new_n1024), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1030), .B(new_n1031), .C1(new_n1032), .C2(new_n1002), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(KEYINPUT51), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1035));
  AOI211_X1 g610(.A(G2084), .B(new_n964), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1966), .B1(new_n990), .B2(new_n1023), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1031), .B1(new_n1038), .B2(new_n1030), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1019), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1020), .A2(new_n994), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1961), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1016), .A2(KEYINPUT121), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n990), .A2(new_n755), .A3(new_n991), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n877), .A2(new_n959), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n989), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n755), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1055), .B(new_n467), .C1(G2105), .C2(new_n475), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n991), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1049), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1043), .B1(new_n1058), .B2(G171), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n990), .A2(KEYINPUT53), .A3(new_n755), .A4(new_n1023), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1049), .A2(new_n1052), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1059), .B1(new_n585), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1052), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT121), .B1(new_n1020), .B2(new_n994), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1045), .B(new_n964), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1066), .B2(new_n1047), .ZN(new_n1067));
  AOI21_X1  g642(.A(G301), .B1(new_n1067), .B2(new_n1060), .ZN(new_n1068));
  AND4_X1   g643(.A1(G301), .A2(new_n1049), .A3(new_n1052), .A4(new_n1057), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1043), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1042), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT126), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT126), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1042), .A2(new_n1062), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n571), .A2(new_n576), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1956), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n995), .A2(new_n998), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n964), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n990), .A2(new_n991), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1075), .B(KEYINPUT57), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1080), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n990), .A2(new_n991), .ZN(new_n1090));
  INV_X1    g665(.A(new_n968), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1090), .A2(G1996), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n920), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1096));
  XOR2_X1   g671(.A(new_n1095), .B(new_n1096), .Z(new_n1097));
  NAND3_X1  g672(.A1(new_n1083), .A2(KEYINPUT61), .A3(new_n1086), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1089), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1046), .A2(new_n1100), .A3(new_n1048), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1091), .A2(new_n790), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1103), .A2(KEYINPUT123), .A3(new_n620), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n620), .B1(new_n1103), .B2(KEYINPUT123), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1104), .A2(new_n1105), .B1(KEYINPUT123), .B2(new_n1103), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1099), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1083), .A3(new_n619), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1086), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1072), .B(new_n1074), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1008), .B1(new_n1114), .B2(G8), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1038), .A2(G286), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n988), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT63), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n980), .B(KEYINPUT119), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n983), .A2(new_n987), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n718), .A2(new_n969), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n984), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1116), .A2(new_n1126), .A3(new_n1006), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1018), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n988), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1118), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1029), .A2(KEYINPUT51), .A3(new_n1033), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1035), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1029), .B2(KEYINPUT51), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT62), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1041), .A2(new_n1135), .A3(new_n1034), .ZN(new_n1136));
  AND4_X1   g711(.A1(new_n585), .A2(new_n1007), .A3(new_n1018), .A4(new_n1061), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT127), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1134), .A2(new_n1140), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1130), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1113), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1054), .A2(new_n964), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n769), .B(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n785), .A2(G2067), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n783), .A2(new_n790), .A3(new_n784), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n740), .A2(new_n742), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n740), .A2(new_n742), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1146), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(G290), .B(G1986), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1144), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1143), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1148), .B1(new_n1156), .B2(new_n1151), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(new_n1144), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1149), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1144), .B1(new_n1159), .B2(new_n769), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT47), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1144), .ZN(new_n1166));
  NOR4_X1   g741(.A1(new_n1054), .A2(G1986), .A3(G290), .A4(new_n964), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  AOI211_X1 g743(.A(new_n1158), .B(new_n1165), .C1(new_n1166), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1155), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g745(.A1(G227), .A2(new_n459), .ZN(new_n1172));
  AND3_X1   g746(.A1(new_n704), .A2(new_n669), .A3(new_n1172), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n1173), .A2(new_n948), .A3(new_n885), .ZN(G308));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n948), .A3(new_n885), .ZN(G225));
endmodule


