//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  XNOR2_X1  g000(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G137), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT67), .B1(new_n187), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n192), .B1(KEYINPUT11), .B2(new_n189), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n194), .B(new_n195), .C1(new_n197), .C2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n190), .A2(new_n193), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n190), .A2(new_n199), .A3(new_n203), .A4(new_n193), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(KEYINPUT68), .A3(G131), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT0), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n209), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n216), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n207), .A2(new_n208), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n215), .A2(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n205), .A2(new_n206), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n211), .A3(new_n213), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n208), .A2(new_n212), .A3(G143), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n210), .B(G146), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G131), .B1(new_n192), .B2(new_n189), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n204), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n204), .A2(KEYINPUT69), .A3(new_n227), .A4(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(G116), .B(G119), .Z(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT2), .B(G113), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n222), .A2(KEYINPUT30), .A3(new_n229), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n239), .B(KEYINPUT70), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n222), .A2(new_n229), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(G101), .ZN(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n245), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n243), .A2(KEYINPUT71), .A3(new_n248), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT31), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n243), .A2(KEYINPUT71), .A3(new_n248), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT71), .B1(new_n243), .B2(new_n248), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT31), .A3(new_n241), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n234), .A2(new_n239), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n243), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n243), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n248), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n255), .A2(new_n259), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(G472), .A2(G902), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT32), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n266), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n253), .A2(new_n254), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT31), .B1(new_n258), .B2(new_n241), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n268), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT73), .B(G902), .Z(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n222), .A2(new_n229), .ZN(new_n279));
  INV_X1    g093(.A(new_n242), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n243), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT28), .A3(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(KEYINPUT29), .A3(new_n264), .A4(new_n248), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n241), .A2(new_n243), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n248), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n265), .A2(new_n266), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n278), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n270), .A2(new_n276), .B1(G472), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n208), .A2(G119), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n208), .A2(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT74), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT24), .B(G110), .Z(new_n298));
  XNOR2_X1  g112(.A(new_n295), .B(KEYINPUT23), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n294), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT76), .B(G110), .Z(new_n301));
  OAI22_X1  g115(.A1(new_n297), .A2(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G125), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT16), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n303), .A2(KEYINPUT75), .A3(G125), .ZN(new_n307));
  XNOR2_X1  g121(.A(G125), .B(G140), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(KEYINPUT75), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT16), .ZN(new_n310));
  OAI211_X1 g124(.A(G146), .B(new_n306), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n308), .A2(new_n212), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n304), .A3(KEYINPUT75), .ZN(new_n317));
  OR3_X1    g131(.A1(new_n303), .A2(KEYINPUT75), .A3(G125), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n212), .B1(new_n319), .B2(new_n305), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n320), .A2(new_n311), .B1(G110), .B2(new_n300), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n297), .A2(new_n298), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G221), .A3(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT22), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(G137), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n314), .A2(new_n323), .A3(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI22_X1  g146(.A1(new_n332), .A2(new_n277), .B1(KEYINPUT77), .B2(KEYINPUT25), .ZN(new_n333));
  INV_X1    g147(.A(G217), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n278), .B2(G234), .ZN(new_n335));
  NOR2_X1   g149(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n278), .A3(new_n331), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n335), .A2(G902), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n330), .A2(new_n339), .A3(new_n331), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n292), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G475), .A2(G902), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n343), .B(KEYINPUT97), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT98), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(KEYINPUT20), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  INV_X1    g162(.A(G104), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT92), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n317), .A2(new_n351), .A3(new_n318), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n317), .B2(new_n318), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT19), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT94), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT19), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n308), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n358), .B(KEYINPUT19), .C1(new_n352), .C2(new_n353), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n355), .A2(new_n212), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G237), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n325), .A3(G214), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n210), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G131), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n203), .A3(new_n364), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT93), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n311), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n352), .A2(new_n353), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n313), .B1(new_n371), .B2(new_n212), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT18), .A2(G131), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n365), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n350), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n365), .A2(KEYINPUT17), .A3(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n320), .A2(new_n311), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT95), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n368), .A2(KEYINPUT17), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n320), .A2(new_n311), .A3(new_n377), .A4(KEYINPUT95), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n383), .A2(new_n350), .A3(new_n375), .ZN(new_n384));
  OAI221_X1 g198(.A(new_n347), .B1(new_n346), .B2(new_n345), .C1(new_n376), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n370), .A2(new_n375), .ZN(new_n386));
  INV_X1    g200(.A(new_n350), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT96), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n350), .A3(new_n375), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT96), .B1(new_n376), .B2(new_n384), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n344), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n385), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n383), .A2(new_n375), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT99), .B1(new_n396), .B2(new_n387), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n390), .ZN(new_n398));
  INV_X1    g212(.A(G902), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(KEYINPUT99), .A3(new_n387), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G475), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n210), .A2(KEYINPUT13), .A3(G128), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT100), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n208), .A2(G143), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n208), .A2(G143), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n405), .B(new_n406), .C1(KEYINPUT13), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G134), .ZN(new_n409));
  XNOR2_X1  g223(.A(G128), .B(G143), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n188), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT101), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G122), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G116), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(G116), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G107), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(KEYINPUT101), .A3(G134), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n413), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n418), .A2(new_n419), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT14), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n417), .B1(new_n415), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n425), .A2(KEYINPUT102), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(KEYINPUT102), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(KEYINPUT14), .C2(new_n416), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n428), .B2(G107), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n410), .B(G134), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n422), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT9), .B(G234), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n435), .A2(new_n334), .A3(G953), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n422), .A2(new_n432), .A3(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n278), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n325), .A2(G952), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G234), .B2(G237), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n325), .B(new_n278), .C1(G234), .C2(G237), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT21), .B(G898), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G214), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n215), .A2(new_n218), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n219), .A2(new_n220), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n455), .B(G125), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT88), .B1(new_n221), .B2(new_n315), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n315), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n464));
  INV_X1    g278(.A(G224), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G953), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n468));
  INV_X1    g282(.A(new_n466), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n460), .B1(new_n469), .B2(KEYINPUT7), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT3), .B1(new_n349), .B2(G107), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n419), .A3(G104), .ZN(new_n474));
  INV_X1    g288(.A(G101), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n349), .A2(G107), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n419), .A2(G104), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n349), .A2(G107), .ZN(new_n479));
  OAI21_X1  g293(.A(G101), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n237), .A2(new_n238), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT5), .ZN(new_n483));
  INV_X1    g297(.A(G119), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(G116), .ZN(new_n485));
  OAI211_X1 g299(.A(G113), .B(new_n485), .C1(new_n237), .C2(new_n483), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(G110), .B(G122), .Z(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(G101), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT82), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT82), .A4(G101), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(G101), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT4), .A3(new_n477), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n239), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n487), .B(new_n489), .C1(new_n496), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n486), .A2(new_n482), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n477), .A2(new_n480), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT89), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n487), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n488), .B(KEYINPUT8), .Z(new_n505));
  NAND4_X1  g319(.A1(new_n481), .A2(KEYINPUT89), .A3(new_n486), .A4(new_n482), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n467), .A2(new_n471), .A3(new_n500), .A4(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n487), .B1(new_n496), .B2(new_n499), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n488), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT6), .A3(new_n500), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n468), .A2(new_n466), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n458), .A2(new_n459), .A3(new_n462), .A4(new_n469), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n515), .A3(new_n488), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n508), .A2(new_n517), .A3(new_n399), .ZN(new_n518));
  OAI21_X1  g332(.A(G210), .B1(G237), .B2(G902), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT91), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n508), .A2(new_n517), .A3(new_n399), .A4(new_n519), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n454), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n403), .A2(new_n445), .A3(new_n452), .A4(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G221), .B1(new_n435), .B2(G902), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT78), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n205), .A2(new_n206), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT85), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n221), .A2(new_n498), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT83), .B1(new_n496), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n494), .A2(new_n495), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT83), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n498), .A4(new_n221), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT10), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n481), .A2(new_n227), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n461), .B2(new_n502), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n530), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  AOI211_X1 g358(.A(KEYINPUT85), .B(new_n542), .C1(new_n532), .C2(new_n535), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n529), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n542), .B1(new_n532), .B2(new_n535), .ZN(new_n548));
  INV_X1    g362(.A(new_n529), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT86), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n551), .B(new_n529), .C1(new_n544), .C2(new_n545), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT80), .B(G140), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n325), .A2(G227), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT79), .B(G110), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n461), .B(new_n502), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n529), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n562), .A2(new_n563), .B1(new_n548), .B2(new_n549), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n529), .A2(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT12), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(KEYINPUT87), .A3(new_n558), .A4(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n529), .A2(new_n563), .A3(new_n561), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n550), .A2(new_n566), .A3(new_n558), .A4(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT87), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G469), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n278), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n547), .A2(new_n558), .A3(new_n550), .A4(new_n552), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n564), .A2(new_n566), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n559), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(G469), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(G469), .A2(G902), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n528), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n342), .A2(new_n525), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  AOI211_X1 g399(.A(new_n528), .B(new_n341), .C1(new_n576), .C2(new_n582), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n274), .A2(new_n278), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n587), .A2(G472), .B1(new_n268), .B2(new_n274), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n395), .A2(new_n402), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT33), .B1(new_n436), .B2(KEYINPUT104), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n422), .A2(new_n432), .A3(new_n436), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n436), .B1(new_n422), .B2(new_n432), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n591), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n438), .A2(new_n439), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n596), .A3(new_n278), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G478), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n440), .A2(new_n442), .A3(new_n278), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n453), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n519), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n518), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n522), .A2(new_n603), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n452), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n589), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  XNOR2_X1  g427(.A(new_n393), .B(new_n394), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n444), .A3(new_n402), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n609), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n589), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  NOR2_X1   g433(.A1(new_n329), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n324), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n339), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n338), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n528), .B(new_n624), .C1(new_n576), .C2(new_n582), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n525), .A3(new_n588), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT37), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G110), .ZN(G12));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n447), .B1(new_n448), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n615), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n608), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n270), .A2(new_n276), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n291), .A2(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n625), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  NAND2_X1  g451(.A1(new_n590), .A2(new_n444), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n630), .B(KEYINPUT39), .Z(new_n639));
  NAND2_X1  g453(.A1(new_n583), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n454), .B(new_n638), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n521), .A2(new_n522), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT38), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n640), .ZN(new_n646));
  INV_X1    g460(.A(new_n641), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n283), .A2(new_n266), .A3(new_n284), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n253), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n650), .B2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n633), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n623), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n642), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  INV_X1    g470(.A(new_n630), .ZN(new_n657));
  AND4_X1   g471(.A1(KEYINPUT106), .A2(new_n590), .A3(new_n601), .A4(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n600), .B1(new_n395), .B2(new_n402), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT106), .B1(new_n659), .B2(new_n657), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n625), .A3(new_n635), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT107), .B(G146), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G48));
  AOI21_X1  g478(.A(new_n572), .B1(new_n553), .B2(new_n559), .ZN(new_n665));
  OAI21_X1  g479(.A(G469), .B1(new_n665), .B2(new_n277), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n576), .A2(new_n666), .A3(new_n526), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n667), .A2(new_n292), .A3(new_n341), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n610), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT41), .B(G113), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G15));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n616), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G116), .ZN(G18));
  INV_X1    g487(.A(new_n667), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n590), .A2(new_n444), .A3(new_n451), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n635), .A3(new_n675), .A4(new_n623), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G119), .ZN(G21));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT109), .B(G472), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n267), .B2(new_n277), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n268), .B(KEYINPUT108), .Z(new_n681));
  NOR2_X1   g495(.A1(new_n272), .A2(new_n273), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n248), .B1(new_n285), .B2(new_n264), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n678), .B1(new_n685), .B2(new_n341), .ZN(new_n686));
  INV_X1    g500(.A(new_n341), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n680), .A2(new_n684), .A3(new_n687), .A4(KEYINPUT110), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n667), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n638), .B2(new_n632), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n590), .A2(new_n608), .A3(KEYINPUT111), .A4(new_n444), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n451), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  NOR2_X1   g509(.A1(new_n667), .A2(new_n632), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n685), .A2(new_n624), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n661), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  NAND3_X1  g513(.A1(new_n521), .A2(new_n522), .A3(new_n453), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n526), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n581), .B(KEYINPUT112), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n580), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n576), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n701), .B1(new_n705), .B2(KEYINPUT113), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n665), .A2(G469), .A3(new_n277), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n580), .A2(new_n703), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n526), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT114), .B(KEYINPUT42), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n342), .A3(new_n661), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n700), .B1(new_n709), .B2(new_n710), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n705), .A2(KEYINPUT113), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n342), .A3(new_n661), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT114), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n203), .ZN(G33));
  INV_X1    g536(.A(KEYINPUT115), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n712), .A2(new_n723), .A3(new_n342), .A4(new_n631), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n715), .A2(new_n342), .A3(new_n631), .A4(new_n716), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT115), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n577), .A2(new_n579), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT45), .B1(new_n577), .B2(new_n579), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n732), .A2(new_n575), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n703), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n729), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n730), .B(new_n731), .ZN(new_n737));
  OAI211_X1 g551(.A(KEYINPUT46), .B(new_n703), .C1(new_n737), .C2(new_n575), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n738), .A3(new_n576), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n526), .A3(new_n639), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n403), .A2(KEYINPUT43), .A3(new_n601), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n601), .A2(new_n395), .A3(new_n402), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n588), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n623), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n700), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n740), .B(new_n749), .C1(new_n748), .C2(new_n747), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n526), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n739), .A2(KEYINPUT47), .A3(new_n526), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n292), .A2(new_n701), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n341), .A3(new_n661), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  INV_X1    g573(.A(new_n447), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n667), .A2(new_n760), .A3(new_n700), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n652), .A2(new_n341), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n403), .A2(new_n761), .A3(new_n762), .A4(new_n600), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n686), .A2(new_n688), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n760), .B1(new_n741), .B2(new_n744), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n667), .A2(new_n644), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(KEYINPUT50), .A3(new_n454), .A4(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n454), .A3(new_n767), .A4(new_n765), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n763), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n761), .A2(new_n697), .A3(new_n745), .ZN(new_n773));
  INV_X1    g587(.A(new_n755), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT47), .B1(new_n739), .B2(new_n526), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n576), .A2(new_n666), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n527), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT121), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n774), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n766), .A2(new_n701), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n772), .B(new_n773), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n446), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n761), .A2(new_n762), .A3(new_n659), .ZN(new_n785));
  INV_X1    g599(.A(new_n777), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n754), .A2(new_n755), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n781), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n773), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n790), .B(new_n763), .C1(new_n768), .C2(new_n771), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n791), .A3(KEYINPUT122), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT122), .B1(new_n789), .B2(new_n791), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n784), .B(new_n785), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n761), .A2(new_n342), .A3(new_n745), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT48), .Z(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n766), .A2(new_n696), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n789), .A2(new_n791), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n792), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n801), .A3(new_n785), .A4(new_n784), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT123), .B1(new_n807), .B2(new_n799), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n292), .A2(new_n700), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n614), .A2(new_n402), .A3(new_n657), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n625), .A2(new_n809), .A3(new_n445), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n714), .A2(new_n720), .A3(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n625), .B(new_n635), .C1(new_n661), .C2(new_n631), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n691), .A2(new_n692), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n630), .B(KEYINPUT118), .Z(new_n816));
  NOR2_X1   g630(.A1(new_n623), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n652), .A3(new_n705), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n698), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n814), .A2(new_n818), .A3(new_n698), .A4(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n661), .A2(new_n715), .A3(new_n697), .A4(new_n716), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n724), .B2(new_n726), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n694), .A2(new_n669), .A3(new_n672), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n523), .A2(new_n452), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n602), .B1(new_n445), .B2(new_n590), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n586), .A2(new_n588), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n676), .A3(new_n626), .A4(new_n584), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n813), .A2(new_n823), .A3(new_n825), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT53), .B1(new_n823), .B2(KEYINPUT117), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT54), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT119), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(KEYINPUT54), .C1(new_n834), .C2(new_n835), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(KEYINPUT53), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n714), .A2(new_n720), .A3(new_n812), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n676), .A2(new_n626), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n689), .A2(new_n693), .B1(new_n668), .B2(new_n610), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n583), .A2(new_n828), .A3(new_n687), .A4(new_n588), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n292), .A2(new_n524), .A3(new_n341), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n845), .A2(new_n827), .B1(new_n846), .B2(new_n583), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n844), .A3(new_n847), .A4(new_n672), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n823), .A4(new_n825), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n841), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT120), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n855), .B(KEYINPUT54), .C1(new_n841), .C2(new_n851), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n802), .A2(new_n808), .A3(new_n840), .A4(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(G952), .A2(G953), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR4_X1    g674(.A1(new_n528), .A2(new_n742), .A3(new_n341), .A4(new_n454), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n644), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n776), .B(KEYINPUT49), .Z(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n653), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n860), .A2(new_n866), .ZN(G75));
  NOR2_X1   g681(.A1(new_n852), .A2(new_n278), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT56), .B1(new_n868), .B2(new_n605), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n511), .A2(new_n516), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(new_n514), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT55), .Z(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g688(.A(KEYINPUT56), .B(new_n872), .C1(new_n868), .C2(new_n520), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n325), .A2(G952), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G51));
  XNOR2_X1  g691(.A(new_n852), .B(new_n853), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n703), .A2(KEYINPUT57), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n703), .A2(KEYINPUT57), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n574), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n868), .A2(new_n734), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(G54));
  NAND3_X1  g698(.A1(new_n868), .A2(KEYINPUT58), .A3(G475), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n391), .A2(new_n392), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n887), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n876), .ZN(G60));
  INV_X1    g704(.A(new_n876), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n594), .A2(new_n596), .ZN(new_n892));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n878), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n840), .B2(new_n857), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n891), .B(new_n896), .C1(new_n897), .C2(new_n892), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT60), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n841), .A2(new_n851), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n332), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n841), .A2(new_n851), .A3(new_n621), .A4(new_n901), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(KEYINPUT61), .A3(new_n891), .A4(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n904), .A2(KEYINPUT124), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(KEYINPUT124), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n891), .A3(new_n903), .A4(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n908), .A2(KEYINPUT125), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT125), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(G66));
  OAI21_X1  g726(.A(G953), .B1(new_n450), .B2(new_n465), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n831), .B2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n870), .B1(G898), .B2(new_n325), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G69));
  NAND2_X1  g730(.A1(G227), .A2(G900), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n325), .A2(G900), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n758), .A2(new_n750), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n814), .A2(new_n698), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n815), .A2(new_n342), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n740), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n721), .B1(new_n726), .B2(new_n724), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n918), .B1(new_n925), .B2(new_n325), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n236), .A2(new_n240), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(G953), .B(new_n917), .C1(new_n928), .C2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n926), .A2(new_n927), .ZN(new_n934));
  AOI211_X1 g748(.A(KEYINPUT126), .B(new_n918), .C1(new_n925), .C2(new_n325), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n917), .A2(G953), .ZN(new_n937));
  INV_X1    g751(.A(new_n920), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n655), .A2(new_n938), .A3(KEYINPUT62), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT62), .B1(new_n655), .B2(new_n938), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n646), .A2(new_n342), .A3(new_n701), .A4(new_n828), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n919), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n932), .B1(new_n945), .B2(G953), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n936), .A2(new_n937), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n933), .A2(new_n947), .ZN(G72));
  INV_X1    g762(.A(new_n288), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n919), .A2(new_n831), .A3(new_n923), .A4(new_n924), .ZN(new_n950));
  NAND2_X1  g764(.A1(G472), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT63), .Z(new_n952));
  AOI211_X1 g766(.A(new_n248), .B(new_n949), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n944), .B2(new_n848), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n248), .A3(new_n949), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n891), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n253), .B1(new_n288), .B2(new_n248), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n952), .B(new_n957), .C1(new_n834), .C2(new_n835), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n953), .B(new_n956), .C1(new_n960), .C2(new_n961), .ZN(G57));
endmodule


