

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600;

  NOR2_X1 U328 ( .A1(n514), .A2(n489), .ZN(n583) );
  XNOR2_X1 U329 ( .A(n334), .B(n333), .ZN(n376) );
  INV_X1 U330 ( .A(G36GAT), .ZN(n331) );
  XNOR2_X1 U331 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U332 ( .A(n338), .B(n450), .ZN(n339) );
  XOR2_X1 U333 ( .A(KEYINPUT38), .B(n468), .Z(n520) );
  NOR2_X1 U334 ( .A1(n536), .A2(n538), .ZN(n381) );
  XOR2_X1 U335 ( .A(G113GAT), .B(KEYINPUT0), .Z(n355) );
  XNOR2_X1 U336 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n487) );
  INV_X1 U337 ( .A(n430), .ZN(n303) );
  XNOR2_X1 U338 ( .A(n332), .B(n331), .ZN(n334) );
  XNOR2_X1 U339 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U340 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U341 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U342 ( .A(KEYINPUT123), .B(KEYINPUT55), .ZN(n491) );
  XNOR2_X1 U343 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U344 ( .A(n467), .B(n466), .ZN(n590) );
  XNOR2_X1 U345 ( .A(n340), .B(n339), .ZN(n344) );
  NOR2_X1 U346 ( .A1(n538), .A2(n493), .ZN(n579) );
  XOR2_X1 U347 ( .A(KEYINPUT41), .B(n477), .Z(n565) );
  XOR2_X1 U348 ( .A(n315), .B(n380), .Z(n547) );
  XNOR2_X1 U349 ( .A(n494), .B(G176GAT), .ZN(n495) );
  XNOR2_X1 U350 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U351 ( .A(n496), .B(n495), .ZN(G1349GAT) );
  XNOR2_X1 U352 ( .A(n472), .B(n471), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U354 ( .A(G134GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n308) );
  XOR2_X1 U356 ( .A(G99GAT), .B(n355), .Z(n299) );
  XOR2_X1 U357 ( .A(G120GAT), .B(G71GAT), .Z(n463) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(n463), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n299), .B(n298), .ZN(n306) );
  XOR2_X1 U360 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n301) );
  NAND2_X1 U361 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U362 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(n302), .ZN(n304) );
  XOR2_X1 U364 ( .A(G15GAT), .B(G127GAT), .Z(n430) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n315) );
  XOR2_X1 U366 ( .A(G183GAT), .B(KEYINPUT87), .Z(n310) );
  XNOR2_X1 U367 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U369 ( .A(KEYINPUT88), .B(KEYINPUT18), .Z(n312) );
  XNOR2_X1 U370 ( .A(KEYINPUT19), .B(KEYINPUT89), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n380) );
  INV_X1 U373 ( .A(KEYINPUT10), .ZN(n319) );
  XOR2_X1 U374 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n317) );
  XNOR2_X1 U375 ( .A(KEYINPUT75), .B(KEYINPUT64), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n321) );
  NAND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n324) );
  INV_X1 U380 ( .A(n324), .ZN(n322) );
  NAND2_X1 U381 ( .A1(n322), .A2(KEYINPUT11), .ZN(n326) );
  INV_X1 U382 ( .A(KEYINPUT11), .ZN(n323) );
  NAND2_X1 U383 ( .A1(n324), .A2(n323), .ZN(n325) );
  NAND2_X1 U384 ( .A1(n326), .A2(n325), .ZN(n336) );
  INV_X1 U385 ( .A(KEYINPUT77), .ZN(n327) );
  NAND2_X1 U386 ( .A1(G92GAT), .A2(n327), .ZN(n330) );
  INV_X1 U387 ( .A(G92GAT), .ZN(n328) );
  NAND2_X1 U388 ( .A1(n328), .A2(KEYINPUT77), .ZN(n329) );
  NAND2_X1 U389 ( .A1(n330), .A2(n329), .ZN(n332) );
  XNOR2_X1 U390 ( .A(G190GAT), .B(G218GAT), .ZN(n333) );
  XOR2_X1 U391 ( .A(n376), .B(KEYINPUT73), .Z(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n340) );
  XNOR2_X1 U393 ( .A(G50GAT), .B(G162GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n337), .B(G106GAT), .ZN(n395) );
  XOR2_X1 U395 ( .A(G134GAT), .B(KEYINPUT76), .Z(n354) );
  XNOR2_X1 U396 ( .A(n395), .B(n354), .ZN(n338) );
  XOR2_X1 U397 ( .A(G99GAT), .B(G85GAT), .Z(n450) );
  XOR2_X1 U398 ( .A(KEYINPUT7), .B(KEYINPUT65), .Z(n342) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(G29GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U401 ( .A(KEYINPUT8), .B(n343), .ZN(n448) );
  XOR2_X1 U402 ( .A(n344), .B(n448), .Z(n573) );
  XNOR2_X1 U403 ( .A(KEYINPUT78), .B(n573), .ZN(n498) );
  XNOR2_X1 U404 ( .A(KEYINPUT36), .B(KEYINPUT107), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n498), .B(n345), .ZN(n597) );
  XOR2_X1 U406 ( .A(KEYINPUT1), .B(KEYINPUT98), .Z(n347) );
  XNOR2_X1 U407 ( .A(G148GAT), .B(KEYINPUT4), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U409 ( .A(G155GAT), .B(G162GAT), .Z(n349) );
  XNOR2_X1 U410 ( .A(G127GAT), .B(G120GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n368) );
  XOR2_X1 U413 ( .A(KEYINPUT96), .B(G57GAT), .Z(n353) );
  XNOR2_X1 U414 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n359) );
  XOR2_X1 U416 ( .A(G85GAT), .B(n354), .Z(n357) );
  XNOR2_X1 U417 ( .A(G29GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U419 ( .A(n359), .B(n358), .Z(n361) );
  NAND2_X1 U420 ( .A1(G225GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n362), .B(KEYINPUT5), .Z(n366) );
  XOR2_X1 U423 ( .A(KEYINPUT92), .B(KEYINPUT3), .Z(n364) );
  XNOR2_X1 U424 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n393) );
  XNOR2_X1 U426 ( .A(n393), .B(KEYINPUT6), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U428 ( .A(n368), .B(n367), .Z(n534) );
  XOR2_X1 U429 ( .A(G8GAT), .B(KEYINPUT79), .Z(n426) );
  XOR2_X1 U430 ( .A(KEYINPUT99), .B(n426), .Z(n370) );
  NAND2_X1 U431 ( .A1(G226GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n373) );
  XOR2_X1 U433 ( .A(KEYINPUT70), .B(G64GAT), .Z(n372) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G204GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n459) );
  XOR2_X1 U436 ( .A(n373), .B(n459), .Z(n378) );
  XOR2_X1 U437 ( .A(G211GAT), .B(KEYINPUT21), .Z(n375) );
  XNOR2_X1 U438 ( .A(G197GAT), .B(KEYINPUT91), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n394) );
  XNOR2_X1 U440 ( .A(n394), .B(n376), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U442 ( .A(n380), .B(n379), .Z(n517) );
  INV_X1 U443 ( .A(n517), .ZN(n536) );
  INV_X1 U444 ( .A(n547), .ZN(n538) );
  XOR2_X1 U445 ( .A(KEYINPUT102), .B(n381), .Z(n400) );
  XOR2_X1 U446 ( .A(KEYINPUT22), .B(KEYINPUT94), .Z(n383) );
  NAND2_X1 U447 ( .A1(G228GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U449 ( .A(KEYINPUT95), .B(n384), .ZN(n391) );
  XOR2_X1 U450 ( .A(G204GAT), .B(KEYINPUT23), .Z(n386) );
  XNOR2_X1 U451 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n385) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U453 ( .A(n387), .B(KEYINPUT90), .Z(n389) );
  XOR2_X1 U454 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  XNOR2_X1 U455 ( .A(n425), .B(G218GAT), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n399) );
  XOR2_X1 U458 ( .A(G78GAT), .B(KEYINPUT69), .Z(n392) );
  XOR2_X1 U459 ( .A(G148GAT), .B(n392), .Z(n458) );
  XOR2_X1 U460 ( .A(n458), .B(n393), .Z(n397) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n490) );
  NAND2_X1 U464 ( .A1(n400), .A2(n490), .ZN(n401) );
  XOR2_X1 U465 ( .A(KEYINPUT25), .B(n401), .Z(n405) );
  XNOR2_X1 U466 ( .A(n517), .B(KEYINPUT27), .ZN(n408) );
  NOR2_X1 U467 ( .A1(n547), .A2(n490), .ZN(n402) );
  XOR2_X1 U468 ( .A(KEYINPUT26), .B(n402), .Z(n403) );
  XNOR2_X1 U469 ( .A(KEYINPUT101), .B(n403), .ZN(n582) );
  NAND2_X1 U470 ( .A1(n408), .A2(n582), .ZN(n404) );
  NAND2_X1 U471 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U472 ( .A1(n534), .A2(n406), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n407), .B(KEYINPUT103), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT28), .B(n490), .Z(n519) );
  INV_X1 U475 ( .A(n519), .ZN(n541) );
  INV_X1 U476 ( .A(n534), .ZN(n514) );
  NAND2_X1 U477 ( .A1(n408), .A2(n514), .ZN(n409) );
  XOR2_X1 U478 ( .A(KEYINPUT100), .B(n409), .Z(n561) );
  NAND2_X1 U479 ( .A1(n541), .A2(n561), .ZN(n549) );
  NOR2_X1 U480 ( .A1(n549), .A2(n547), .ZN(n410) );
  NOR2_X1 U481 ( .A1(n411), .A2(n410), .ZN(n497) );
  NOR2_X1 U482 ( .A1(n597), .A2(n497), .ZN(n433) );
  XOR2_X1 U483 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n417) );
  XNOR2_X1 U484 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n412) );
  XNOR2_X1 U485 ( .A(n412), .B(KEYINPUT66), .ZN(n437) );
  XOR2_X1 U486 ( .A(KEYINPUT15), .B(KEYINPUT83), .Z(n414) );
  XNOR2_X1 U487 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n413) );
  XNOR2_X1 U488 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U489 ( .A(n437), .B(n415), .ZN(n416) );
  XNOR2_X1 U490 ( .A(n417), .B(n416), .ZN(n424) );
  XOR2_X1 U491 ( .A(KEYINPUT80), .B(G64GAT), .Z(n419) );
  XNOR2_X1 U492 ( .A(G211GAT), .B(G78GAT), .ZN(n418) );
  XNOR2_X1 U493 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U494 ( .A(G57GAT), .B(KEYINPUT13), .Z(n451) );
  XOR2_X1 U495 ( .A(n420), .B(n451), .Z(n422) );
  XNOR2_X1 U496 ( .A(G183GAT), .B(G71GAT), .ZN(n421) );
  XNOR2_X1 U497 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U498 ( .A(n424), .B(n423), .Z(n432) );
  XOR2_X1 U499 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U500 ( .A1(G231GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U501 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U502 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U503 ( .A(n432), .B(n431), .Z(n577) );
  INV_X1 U504 ( .A(n577), .ZN(n594) );
  NAND2_X1 U505 ( .A1(n433), .A2(n594), .ZN(n434) );
  XNOR2_X1 U506 ( .A(n434), .B(KEYINPUT37), .ZN(n533) );
  XOR2_X1 U507 ( .A(G141GAT), .B(G197GAT), .Z(n436) );
  XNOR2_X1 U508 ( .A(G113GAT), .B(G22GAT), .ZN(n435) );
  XNOR2_X1 U509 ( .A(n436), .B(n435), .ZN(n447) );
  XOR2_X1 U510 ( .A(G50GAT), .B(G36GAT), .Z(n439) );
  XNOR2_X1 U511 ( .A(G15GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U512 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U513 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n441) );
  NAND2_X1 U514 ( .A1(G229GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U515 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U516 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U517 ( .A(G169GAT), .B(G8GAT), .Z(n444) );
  XNOR2_X1 U518 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U519 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U520 ( .A(n449), .B(n448), .ZN(n575) );
  INV_X1 U521 ( .A(n575), .ZN(n585) );
  XOR2_X1 U522 ( .A(n451), .B(n450), .Z(n453) );
  NAND2_X1 U523 ( .A1(G230GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U524 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U525 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n455) );
  XNOR2_X1 U526 ( .A(KEYINPUT32), .B(KEYINPUT68), .ZN(n454) );
  XNOR2_X1 U527 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U528 ( .A(n457), .B(n456), .Z(n467) );
  XOR2_X1 U529 ( .A(n459), .B(n458), .Z(n465) );
  XOR2_X1 U530 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n461) );
  XNOR2_X1 U531 ( .A(G106GAT), .B(G92GAT), .ZN(n460) );
  XNOR2_X1 U532 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U533 ( .A(n463), .B(n462), .ZN(n464) );
  INV_X1 U534 ( .A(n590), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n585), .A2(n477), .ZN(n501) );
  NAND2_X1 U536 ( .A1(n533), .A2(n501), .ZN(n468) );
  NAND2_X1 U537 ( .A1(n547), .A2(n520), .ZN(n472) );
  XOR2_X1 U538 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n470) );
  XNOR2_X1 U539 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n469) );
  NOR2_X1 U540 ( .A1(n594), .A2(n597), .ZN(n474) );
  INV_X1 U541 ( .A(KEYINPUT45), .ZN(n473) );
  XNOR2_X1 U542 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U543 ( .A1(n475), .A2(n477), .ZN(n476) );
  NAND2_X1 U544 ( .A1(n476), .A2(n585), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n565), .A2(n575), .ZN(n478) );
  XNOR2_X1 U546 ( .A(KEYINPUT46), .B(n478), .ZN(n479) );
  NAND2_X1 U547 ( .A1(n479), .A2(n594), .ZN(n480) );
  NOR2_X1 U548 ( .A1(n573), .A2(n480), .ZN(n481) );
  XOR2_X1 U549 ( .A(KEYINPUT47), .B(n481), .Z(n482) );
  XNOR2_X1 U550 ( .A(n482), .B(KEYINPUT115), .ZN(n483) );
  NAND2_X1 U551 ( .A1(n484), .A2(n483), .ZN(n545) );
  XNOR2_X1 U552 ( .A(n545), .B(KEYINPUT48), .ZN(n486) );
  XOR2_X1 U553 ( .A(KEYINPUT121), .B(n517), .Z(n485) );
  NAND2_X1 U554 ( .A1(n486), .A2(n485), .ZN(n488) );
  NAND2_X1 U555 ( .A1(n490), .A2(n583), .ZN(n492) );
  NAND2_X1 U556 ( .A1(n579), .A2(n565), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n494) );
  NOR2_X1 U558 ( .A1(n594), .A2(n498), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT16), .B(n499), .Z(n500) );
  NOR2_X1 U560 ( .A1(n497), .A2(n500), .ZN(n522) );
  NAND2_X1 U561 ( .A1(n501), .A2(n522), .ZN(n510) );
  NOR2_X1 U562 ( .A1(n534), .A2(n510), .ZN(n503) );
  XNOR2_X1 U563 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U565 ( .A(G1GAT), .B(n504), .Z(G1324GAT) );
  NOR2_X1 U566 ( .A1(n536), .A2(n510), .ZN(n505) );
  XOR2_X1 U567 ( .A(G8GAT), .B(n505), .Z(G1325GAT) );
  NOR2_X1 U568 ( .A1(n510), .A2(n538), .ZN(n509) );
  XOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n507) );
  XNOR2_X1 U570 ( .A(G15GAT), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  NOR2_X1 U573 ( .A1(n541), .A2(n510), .ZN(n511) );
  XOR2_X1 U574 ( .A(G22GAT), .B(n511), .Z(G1327GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n513) );
  XNOR2_X1 U576 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n516) );
  NAND2_X1 U578 ( .A1(n520), .A2(n514), .ZN(n515) );
  XOR2_X1 U579 ( .A(n516), .B(n515), .Z(G1328GAT) );
  NAND2_X1 U580 ( .A1(n520), .A2(n517), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n521), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U584 ( .A1(n585), .A2(n565), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n532), .A2(n522), .ZN(n528) );
  NOR2_X1 U586 ( .A1(n534), .A2(n528), .ZN(n523) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n523), .Z(n524) );
  XNOR2_X1 U588 ( .A(KEYINPUT42), .B(n524), .ZN(G1332GAT) );
  NOR2_X1 U589 ( .A1(n536), .A2(n528), .ZN(n525) );
  XOR2_X1 U590 ( .A(G64GAT), .B(n525), .Z(G1333GAT) );
  NOR2_X1 U591 ( .A1(n538), .A2(n528), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT112), .B(n526), .Z(n527) );
  XNOR2_X1 U593 ( .A(G71GAT), .B(n527), .ZN(G1334GAT) );
  NOR2_X1 U594 ( .A1(n541), .A2(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT43), .B(KEYINPUT113), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U597 ( .A(G78GAT), .B(n531), .Z(G1335GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n540) );
  NOR2_X1 U599 ( .A1(n534), .A2(n540), .ZN(n535) );
  XOR2_X1 U600 ( .A(G85GAT), .B(n535), .Z(G1336GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n540), .ZN(n537) );
  XOR2_X1 U602 ( .A(G92GAT), .B(n537), .Z(G1337GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n540), .ZN(n539) );
  XOR2_X1 U604 ( .A(G99GAT), .B(n539), .Z(G1338GAT) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U606 ( .A(KEYINPUT114), .B(KEYINPUT44), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U608 ( .A(G106GAT), .B(n544), .Z(G1339GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT48), .B(n545), .Z(n563) );
  INV_X1 U610 ( .A(n563), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n575), .A2(n558), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n550), .B(KEYINPUT116), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G113GAT), .B(n551), .ZN(G1340GAT) );
  XOR2_X1 U616 ( .A(G120GAT), .B(KEYINPUT49), .Z(n553) );
  NAND2_X1 U617 ( .A1(n558), .A2(n565), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1341GAT) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n555) );
  NAND2_X1 U621 ( .A1(n558), .A2(n577), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1342GAT) );
  XOR2_X1 U624 ( .A(G134GAT), .B(KEYINPUT51), .Z(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n498), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1343GAT) );
  NAND2_X1 U627 ( .A1(n582), .A2(n561), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n572), .A2(n575), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G141GAT), .B(n564), .ZN(G1344GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n567) );
  NAND2_X1 U632 ( .A1(n572), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U634 ( .A(G148GAT), .B(KEYINPUT52), .Z(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1345GAT) );
  NAND2_X1 U636 ( .A1(n577), .A2(n572), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT120), .ZN(n571) );
  XNOR2_X1 U638 ( .A(G155GAT), .B(n571), .ZN(G1346GAT) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U641 ( .A1(n575), .A2(n579), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U643 ( .A1(n577), .A2(n579), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U645 ( .A1(n579), .A2(n498), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT58), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT124), .B(n584), .ZN(n596) );
  NOR2_X1 U650 ( .A1(n596), .A2(n585), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  NOR2_X1 U655 ( .A1(n596), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(G204GAT), .B(n593), .ZN(G1353GAT) );
  NOR2_X1 U659 ( .A1(n594), .A2(n596), .ZN(n595) );
  XOR2_X1 U660 ( .A(G211GAT), .B(n595), .Z(G1354GAT) );
  XNOR2_X1 U661 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n599) );
  NOR2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U663 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U664 ( .A(G218GAT), .B(n600), .ZN(G1355GAT) );
endmodule

