//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT64), .B1(new_n190), .B2(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G146), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n195), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n190), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  OAI21_X1  g016(.A(G128), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n196), .A2(new_n198), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n200), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n207), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G224), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n214), .B(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(new_n217), .B(KEYINPUT85), .Z(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n219), .A2(KEYINPUT3), .A3(G107), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT78), .A2(G104), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT78), .A2(G104), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G107), .ZN(new_n229));
  NOR4_X1   g043(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT79), .A4(new_n221), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n225), .B(new_n226), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n224), .B1(G104), .B2(new_n221), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT81), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT68), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n239), .A3(G119), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n236), .B2(G119), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G113), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n236), .A2(G119), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(new_n244), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n243), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT81), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n231), .A2(new_n250), .A3(new_n233), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n235), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n225), .B1(new_n229), .B2(new_n230), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G101), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n241), .B(new_n242), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n257), .A3(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n252), .A2(new_n259), .A3(KEYINPUT84), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G122), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n252), .A2(new_n259), .A3(new_n264), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT6), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n264), .B1(new_n260), .B2(new_n261), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT6), .A3(new_n263), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n218), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n206), .A2(KEYINPUT87), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n206), .A2(KEYINPUT87), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n213), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT88), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT7), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n276), .A2(new_n277), .B1(new_n215), .B2(G224), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n276), .B2(new_n277), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n214), .B1(G224), .B2(new_n215), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n275), .A2(new_n279), .B1(new_n280), .B2(KEYINPUT7), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(new_n267), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n252), .A2(KEYINPUT86), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n264), .B(KEYINPUT8), .ZN(new_n284));
  INV_X1    g098(.A(new_n252), .ZN(new_n285));
  INV_X1    g099(.A(new_n234), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT86), .B1(new_n286), .B2(new_n249), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n189), .B1(new_n272), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n218), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n270), .A2(KEYINPUT6), .A3(new_n263), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n270), .A2(new_n263), .B1(KEYINPUT6), .B2(new_n267), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n282), .B2(new_n288), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n188), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT89), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G125), .B(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n193), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n301), .B(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n304), .B2(new_n193), .ZN(new_n305));
  NOR2_X1   g119(.A1(G237), .A2(G953), .ZN(new_n306));
  AOI21_X1  g120(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT18), .A2(G131), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n309), .ZN(new_n312));
  OAI211_X1 g126(.A(KEYINPUT18), .B(G131), .C1(new_n312), .C2(new_n307), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n305), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G113), .B(G122), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(new_n219), .ZN(new_n316));
  OAI21_X1  g130(.A(G131), .B1(new_n312), .B2(new_n307), .ZN(new_n317));
  INV_X1    g131(.A(G131), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n308), .A2(new_n318), .A3(new_n309), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT17), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n301), .A2(KEYINPUT16), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n193), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(G146), .A3(new_n323), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT17), .B(G131), .C1(new_n312), .C2(new_n307), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n321), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n314), .A2(new_n316), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n329), .A2(KEYINPUT91), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT91), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n314), .A2(new_n328), .A3(new_n331), .A4(new_n316), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n326), .B(KEYINPUT75), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n301), .B(KEYINPUT90), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT19), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT19), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n301), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n193), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n317), .A2(new_n319), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n334), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n341), .A2(new_n314), .ZN(new_n342));
  OAI22_X1  g156(.A1(new_n330), .A2(new_n333), .B1(new_n342), .B2(new_n316), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n344));
  INV_X1    g158(.A(G475), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n290), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n316), .B1(new_n341), .B2(new_n314), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n329), .A2(KEYINPUT91), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n332), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n290), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT20), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n314), .A2(new_n328), .ZN(new_n353));
  INV_X1    g167(.A(new_n316), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n330), .B2(new_n333), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n290), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n348), .A2(new_n332), .B1(new_n354), .B2(new_n353), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT92), .B1(new_n359), .B2(G902), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n360), .A3(G475), .ZN(new_n361));
  NAND2_X1  g175(.A1(G234), .A2(G237), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G952), .A3(new_n215), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n363), .B(KEYINPUT98), .Z(new_n364));
  AND3_X1   g178(.A1(new_n362), .A2(G902), .A3(G953), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT21), .B(G898), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n352), .A2(new_n361), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G478), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT15), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G134), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n197), .A2(G143), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT13), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n190), .A2(G128), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n197), .A2(G143), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT13), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(KEYINPUT93), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT93), .B1(new_n377), .B2(new_n380), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(new_n379), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G134), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n237), .A2(new_n239), .A3(G122), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n236), .A2(G122), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n221), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n221), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT94), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n392), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n386), .B1(new_n395), .B2(new_n390), .ZN(new_n396));
  INV_X1    g210(.A(new_n383), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n381), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT94), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n388), .A2(new_n403), .A3(new_n389), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G107), .B1(new_n388), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n388), .A2(new_n403), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n408), .A2(KEYINPUT95), .A3(G107), .A4(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n385), .A2(G134), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n391), .B1(new_n387), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT9), .B(G234), .Z(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT77), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n415), .A2(new_n416), .A3(G953), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n401), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n417), .B1(new_n401), .B2(new_n413), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n290), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT96), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n384), .A2(new_n393), .A3(KEYINPUT94), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n399), .B1(new_n396), .B2(new_n398), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n413), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n417), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n401), .A2(new_n413), .A3(new_n417), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT96), .A3(new_n290), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n373), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n420), .A2(new_n372), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT97), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT96), .B1(new_n429), .B2(new_n290), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n421), .B(G902), .C1(new_n427), .C2(new_n428), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n372), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n437));
  INV_X1    g251(.A(new_n432), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n370), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(KEYINPUT89), .B(new_n189), .C1(new_n272), .C2(new_n291), .ZN(new_n441));
  AND4_X1   g255(.A1(new_n187), .A2(new_n300), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n444));
  INV_X1    g258(.A(new_n212), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n258), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n255), .A2(KEYINPUT80), .A3(new_n445), .A4(new_n258), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n231), .A2(new_n250), .A3(new_n233), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n250), .B1(new_n231), .B2(new_n233), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT10), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n204), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n203), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(new_n196), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n198), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n286), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n452), .A2(new_n454), .B1(new_n459), .B2(new_n453), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT11), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n374), .B2(G137), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n374), .A2(G137), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT11), .A3(G134), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G131), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n462), .A2(new_n465), .A3(new_n318), .A4(new_n463), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n449), .A2(new_n460), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n215), .A2(G227), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n470), .B1(new_n449), .B2(new_n460), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n204), .B1(new_n450), .B2(new_n451), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n480), .A2(KEYINPUT82), .B1(new_n286), .B2(new_n458), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(new_n204), .C1(new_n450), .C2(new_n451), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n479), .B(new_n470), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n459), .A3(new_n483), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT12), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n471), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n478), .B1(new_n488), .B2(new_n474), .ZN(new_n489));
  OAI21_X1  g303(.A(G469), .B1(new_n489), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(KEYINPUT83), .B(G469), .C1(new_n489), .C2(G902), .ZN(new_n493));
  INV_X1    g307(.A(G469), .ZN(new_n494));
  INV_X1    g308(.A(new_n487), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n486), .A2(KEYINPUT12), .A3(new_n469), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n476), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n477), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n475), .B1(new_n498), .B2(new_n471), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n494), .B(new_n290), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n493), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n442), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n442), .A2(new_n501), .A3(KEYINPUT99), .A4(new_n502), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT31), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT65), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n212), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT65), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n469), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n374), .A2(G137), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n464), .A2(G134), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n468), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT66), .B1(new_n204), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n203), .A2(new_n200), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n457), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n468), .A4(new_n515), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n512), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT67), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT67), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n516), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n519), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n445), .A2(new_n469), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n445), .A2(new_n469), .A3(KEYINPUT69), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n530), .A2(KEYINPUT30), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n525), .A2(new_n256), .A3(new_n527), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n256), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n530), .A2(new_n537), .A3(new_n533), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n306), .A2(G210), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n540), .B(KEYINPUT27), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT26), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n226), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n508), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n536), .A2(KEYINPUT31), .A3(new_n538), .A4(new_n543), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n537), .A2(new_n531), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n516), .B(KEYINPUT70), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n204), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT71), .B(new_n548), .C1(new_n549), .C2(new_n551), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n522), .A2(new_n256), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n538), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT28), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n543), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n547), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n563));
  OR3_X1    g377(.A1(new_n563), .A2(G472), .A3(G902), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(G472), .B2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(KEYINPUT73), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n560), .B1(new_n545), .B2(new_n546), .ZN(new_n569));
  INV_X1    g383(.A(new_n566), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT74), .B(KEYINPUT32), .Z(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n539), .A2(new_n543), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n554), .A2(new_n555), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n533), .A2(new_n534), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n256), .B1(new_n551), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n538), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(KEYINPUT28), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n543), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n556), .A2(new_n559), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT29), .ZN(new_n584));
  OAI221_X1 g398(.A(new_n290), .B1(new_n575), .B2(KEYINPUT29), .C1(new_n582), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G472), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT32), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n569), .A2(new_n587), .A3(new_n570), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n573), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(G119), .B2(new_n197), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT23), .B1(new_n197), .B2(G119), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT24), .B(G110), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(G119), .B(G128), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n594), .A2(G110), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n334), .A2(new_n302), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n325), .A2(new_n326), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n594), .A2(G110), .B1(new_n596), .B2(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT22), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G137), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n603), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT76), .Z(new_n608));
  INV_X1    g422(.A(G234), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n609), .B2(G217), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G217), .B1(new_n609), .B2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n607), .A2(new_n290), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(KEYINPUT25), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(KEYINPUT25), .B2(new_n613), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n590), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n507), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  NAND2_X1  g433(.A1(new_n501), .A2(new_n502), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n567), .A2(new_n571), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n562), .A2(new_n622), .A3(new_n290), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT100), .B1(new_n569), .B2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(G472), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n621), .A2(new_n616), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n292), .A2(new_n298), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n187), .ZN(new_n629));
  AOI21_X1  g443(.A(G478), .B1(new_n422), .B2(new_n430), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n425), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT33), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n429), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n427), .A2(new_n632), .A3(KEYINPUT33), .A4(new_n428), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n371), .A2(G902), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n352), .A2(new_n361), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n629), .A2(new_n368), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n627), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(new_n639), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n645), .A2(new_n433), .A3(new_n439), .A4(new_n369), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n627), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NAND2_X1  g464(.A1(new_n621), .A2(new_n625), .ZN(new_n651));
  INV_X1    g465(.A(new_n606), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n603), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n610), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n615), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n507), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NOR2_X1   g475(.A1(new_n629), .A2(new_n657), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n501), .A2(new_n662), .A3(new_n502), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n433), .A2(new_n439), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n365), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n364), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n664), .A2(new_n645), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n590), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XOR2_X1   g486(.A(new_n667), .B(KEYINPUT39), .Z(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n620), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT40), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n433), .A2(new_n439), .A3(new_n187), .A4(new_n639), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n656), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT103), .Z(new_n679));
  AOI21_X1  g493(.A(new_n544), .B1(new_n536), .B2(new_n538), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n290), .B1(new_n579), .B2(new_n543), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT102), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n573), .A2(new_n589), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n300), .A2(new_n441), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT38), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n679), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n676), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  INV_X1    g504(.A(new_n640), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n590), .A2(new_n691), .A3(new_n668), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n663), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n193), .ZN(G48));
  NOR2_X1   g508(.A1(new_n497), .A2(new_n499), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n502), .A3(new_n500), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n641), .A2(new_n590), .A3(new_n616), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  AND4_X1   g514(.A1(new_n616), .A2(new_n590), .A3(new_n647), .A4(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n236), .ZN(G18));
  INV_X1    g516(.A(new_n629), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n440), .A2(new_n656), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n590), .A2(new_n697), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  OAI21_X1  g520(.A(G472), .B1(new_n569), .B2(G902), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n547), .B1(new_n543), .B2(new_n580), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n566), .B(KEYINPUT104), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n616), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n677), .B1(new_n292), .B2(new_n298), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n697), .A2(new_n711), .A3(new_n712), .A4(new_n369), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  OAI211_X1 g528(.A(new_n639), .B(new_n668), .C1(new_n630), .C2(new_n637), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT105), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n638), .A2(new_n717), .A3(new_n639), .A4(new_n668), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n710), .A2(new_n656), .A3(new_n707), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n719), .A2(new_n697), .A3(new_n703), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n490), .A2(new_n725), .A3(new_n500), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(new_n490), .B2(new_n500), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n502), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT107), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n502), .C1(new_n726), .C2(new_n727), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n686), .A2(new_n187), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n617), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n716), .A2(new_n718), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n724), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT32), .B1(new_n562), .B2(new_n566), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT108), .B1(new_n736), .B2(new_n588), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n586), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n736), .A2(new_n588), .A3(KEYINPUT108), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n616), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n740), .A2(new_n724), .A3(new_n734), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n731), .A3(new_n729), .A4(new_n732), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  INV_X1    g558(.A(new_n669), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n733), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n374), .ZN(G36));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  OAI21_X1  g562(.A(G469), .B1(new_n489), .B2(KEYINPUT45), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n750), .B(new_n478), .C1(new_n474), .C2(new_n488), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT46), .B(new_n748), .C1(new_n749), .C2(new_n751), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n500), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n502), .ZN(new_n757));
  INV_X1    g571(.A(new_n732), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n674), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n638), .A2(new_n645), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT43), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n651), .B2(new_n656), .ZN(new_n764));
  AOI211_X1 g578(.A(KEYINPUT109), .B(new_n657), .C1(new_n621), .C2(new_n625), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT44), .B(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n759), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  NOR2_X1   g585(.A1(new_n616), .A2(new_n715), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n732), .A2(new_n772), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n773), .A2(KEYINPUT111), .A3(new_n590), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT111), .B1(new_n773), .B2(new_n590), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n757), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n757), .A2(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n776), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  INV_X1    g597(.A(new_n760), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n616), .A3(new_n502), .A4(new_n187), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT112), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n696), .A2(new_n500), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT49), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n786), .A2(new_n685), .A3(new_n687), .A4(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT113), .Z(new_n790));
  NOR2_X1   g604(.A1(new_n761), .A2(new_n364), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n711), .ZN(new_n792));
  INV_X1    g606(.A(new_n697), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n187), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n687), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT50), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n792), .A2(KEYINPUT117), .A3(new_n687), .A4(new_n794), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT118), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n798), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n781), .A2(new_n780), .ZN(new_n805));
  INV_X1    g619(.A(new_n787), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n502), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n732), .B(new_n792), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n758), .A2(new_n793), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n721), .A3(new_n791), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT119), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT119), .ZN(new_n812));
  INV_X1    g626(.A(new_n364), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n616), .A2(new_n809), .A3(new_n813), .A4(new_n685), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n638), .A2(new_n639), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n811), .A2(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n804), .A2(KEYINPUT51), .A3(new_n808), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  INV_X1    g632(.A(new_n803), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n799), .A3(new_n801), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n808), .A2(new_n816), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n823));
  OR2_X1    g637(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n809), .A2(new_n791), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n740), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n814), .A2(new_n691), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n825), .A2(new_n740), .A3(new_n823), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n215), .A2(G952), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n793), .A2(new_n629), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n792), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n817), .A2(new_n822), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n734), .A2(new_n720), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n729), .A2(new_n835), .A3(new_n731), .ZN(new_n836));
  INV_X1    g650(.A(new_n620), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n431), .A2(new_n432), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n657), .A2(new_n639), .A3(new_n667), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n590), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n758), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n746), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n505), .B(new_n506), .C1(new_n617), .C2(new_n658), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n300), .A2(new_n441), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n838), .A2(new_n639), .A3(new_n368), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n844), .A2(new_n845), .A3(new_n187), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n187), .A3(new_n369), .A4(new_n691), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n300), .A2(new_n846), .A3(new_n187), .A4(new_n441), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n701), .B1(new_n627), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n698), .A2(new_n705), .A3(new_n713), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n843), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n842), .A2(new_n743), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n722), .B1(new_n663), .B2(new_n670), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n693), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n656), .A2(new_n667), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n728), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n727), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n490), .A2(new_n725), .A3(new_n500), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(KEYINPUT115), .A3(new_n502), .A4(new_n859), .ZN(new_n865));
  INV_X1    g679(.A(new_n712), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n685), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT52), .B1(new_n857), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n834), .B1(new_n855), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n857), .A2(new_n868), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n857), .A2(new_n868), .A3(KEYINPUT52), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n843), .A2(new_n852), .A3(new_n853), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n746), .A3(new_n841), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT53), .A4(new_n743), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n881), .B1(new_n872), .B2(new_n880), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(KEYINPUT116), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n884), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n882), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n833), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(G952), .A2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n790), .B1(new_n889), .B2(new_n890), .ZN(G75));
  AOI21_X1  g705(.A(new_n290), .B1(new_n872), .B2(new_n880), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n892), .B2(G210), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n294), .A2(new_n295), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT121), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n293), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n893), .A2(new_n897), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n215), .A2(G952), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(new_n695), .B(KEYINPUT122), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n883), .A2(new_n884), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n748), .B(KEYINPUT57), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n749), .A2(new_n751), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n892), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n900), .B1(new_n905), .B2(new_n907), .ZN(G54));
  AND2_X1   g722(.A1(KEYINPUT58), .A2(G475), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n892), .A2(new_n343), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n343), .B1(new_n892), .B2(new_n909), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n910), .A2(new_n911), .A3(new_n900), .ZN(G60));
  INV_X1    g726(.A(new_n900), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n634), .A2(new_n635), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT59), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n903), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n914), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n888), .A2(new_n885), .A3(new_n916), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(new_n872), .A2(new_n880), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n654), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(KEYINPUT123), .A3(new_n913), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n913), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n924), .B1(new_n872), .B2(new_n880), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n608), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n927), .B(KEYINPUT61), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n929), .A2(new_n608), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n900), .B1(new_n929), .B2(new_n654), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n932), .B(new_n933), .C1(KEYINPUT123), .C2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n931), .A2(new_n935), .ZN(G66));
  NAND2_X1  g750(.A1(new_n878), .A2(new_n215), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT124), .ZN(new_n938));
  INV_X1    g752(.A(G224), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n366), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n895), .B1(G898), .B2(new_n215), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  NAND2_X1  g757(.A1(G227), .A2(G900), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n770), .A2(new_n857), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n770), .A2(new_n947), .A3(new_n857), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n746), .ZN(new_n950));
  OR4_X1    g764(.A1(new_n674), .A2(new_n757), .A3(new_n866), .A4(new_n740), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n743), .A2(new_n782), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n949), .A2(KEYINPUT127), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT127), .B1(new_n949), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n215), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n665), .A2(G953), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT125), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n525), .A2(new_n527), .A3(new_n535), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n336), .A2(new_n338), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(new_n962));
  OAI211_X1 g776(.A(G953), .B(new_n944), .C1(new_n959), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n944), .A2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n689), .A2(new_n857), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n838), .A2(new_n639), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n758), .B1(new_n640), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n617), .A3(new_n675), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n782), .A2(new_n970), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n967), .A2(new_n770), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n962), .B1(new_n972), .B2(G953), .ZN(new_n973));
  INV_X1    g787(.A(new_n958), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975));
  INV_X1    g789(.A(new_n948), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n947), .B1(new_n770), .B2(new_n857), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n975), .B1(new_n978), .B2(new_n952), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n949), .A2(KEYINPUT127), .A3(new_n953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n974), .B1(new_n981), .B2(new_n215), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n964), .B(new_n973), .C1(new_n982), .C2(new_n962), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n963), .A2(new_n983), .ZN(G72));
  INV_X1    g798(.A(new_n680), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  NAND4_X1  g801(.A1(new_n922), .A2(new_n575), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n967), .A2(new_n770), .A3(new_n854), .A4(new_n971), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n989), .A2(new_n987), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n913), .B(new_n988), .C1(new_n990), .C2(new_n985), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n979), .A2(new_n854), .A3(new_n980), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n575), .B1(new_n992), .B2(new_n987), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n991), .A2(new_n993), .ZN(G57));
endmodule


