

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(KEYINPUT25), .B(KEYINPUT96), .ZN(n455) );
  XNOR2_X1 U325 ( .A(n342), .B(n341), .ZN(n576) );
  XNOR2_X1 U326 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U327 ( .A(n456), .B(n455), .ZN(n465) );
  XNOR2_X1 U328 ( .A(n332), .B(n331), .ZN(n334) );
  XNOR2_X1 U329 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U330 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U331 ( .A(n478), .B(n477), .ZN(n504) );
  XNOR2_X1 U332 ( .A(n386), .B(n385), .ZN(n524) );
  XOR2_X1 U333 ( .A(G106GAT), .B(G92GAT), .Z(n292) );
  XNOR2_X1 U334 ( .A(KEYINPUT76), .B(KEYINPUT74), .ZN(n293) );
  INV_X1 U335 ( .A(KEYINPUT121), .ZN(n388) );
  INV_X1 U336 ( .A(KEYINPUT94), .ZN(n462) );
  XNOR2_X1 U337 ( .A(n388), .B(KEYINPUT54), .ZN(n389) );
  XNOR2_X1 U338 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U339 ( .A(n298), .B(n293), .ZN(n300) );
  XNOR2_X1 U340 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U341 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n370) );
  XNOR2_X1 U342 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U343 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U344 ( .A(n378), .B(n292), .ZN(n304) );
  XNOR2_X1 U345 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n475) );
  XNOR2_X1 U346 ( .A(n440), .B(n377), .ZN(n382) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U348 ( .A(n476), .B(n475), .ZN(n520) );
  XNOR2_X1 U349 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n477) );
  INV_X1 U350 ( .A(G50GAT), .ZN(n479) );
  INV_X1 U351 ( .A(G36GAT), .ZN(n482) );
  XNOR2_X1 U352 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U353 ( .A(n479), .B(KEYINPUT106), .ZN(n480) );
  XNOR2_X1 U354 ( .A(n482), .B(KEYINPUT104), .ZN(n483) );
  XNOR2_X1 U355 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XNOR2_X1 U356 ( .A(n481), .B(n480), .ZN(G1331GAT) );
  INV_X1 U357 ( .A(KEYINPUT65), .ZN(n414) );
  XNOR2_X1 U358 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n294) );
  XNOR2_X1 U359 ( .A(n294), .B(KEYINPUT8), .ZN(n353) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U361 ( .A(n295), .B(KEYINPUT72), .ZN(n336) );
  XOR2_X1 U362 ( .A(n353), .B(n336), .Z(n307) );
  XOR2_X1 U363 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n297) );
  XNOR2_X1 U364 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n296) );
  XNOR2_X1 U365 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U366 ( .A(G43GAT), .B(G134GAT), .Z(n445) );
  XOR2_X1 U367 ( .A(G50GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U368 ( .A(n445), .B(n415), .ZN(n299) );
  NAND2_X1 U369 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U370 ( .A(n302), .B(n301), .ZN(n305) );
  XNOR2_X1 U371 ( .A(G36GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U372 ( .A(n303), .B(G218GAT), .ZN(n378) );
  XNOR2_X1 U373 ( .A(n307), .B(n306), .ZN(n544) );
  XNOR2_X1 U374 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n308) );
  XNOR2_X1 U375 ( .A(n544), .B(n308), .ZN(n584) );
  XOR2_X1 U376 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n310) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U378 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U379 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n312) );
  XNOR2_X1 U380 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n311) );
  XNOR2_X1 U381 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U382 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U383 ( .A(G22GAT), .B(G155GAT), .Z(n419) );
  XOR2_X1 U384 ( .A(KEYINPUT78), .B(G64GAT), .Z(n316) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U386 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U387 ( .A(n419), .B(n317), .ZN(n318) );
  XNOR2_X1 U388 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U389 ( .A(G211GAT), .B(G71GAT), .Z(n321) );
  XNOR2_X1 U390 ( .A(G183GAT), .B(G127GAT), .ZN(n320) );
  XNOR2_X1 U391 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U392 ( .A(n323), .B(n322), .Z(n325) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n349) );
  XOR2_X1 U394 ( .A(KEYINPUT13), .B(G57GAT), .Z(n330) );
  XNOR2_X1 U395 ( .A(n349), .B(n330), .ZN(n324) );
  XOR2_X1 U396 ( .A(n325), .B(n324), .Z(n560) );
  NOR2_X1 U397 ( .A1(n584), .A2(n560), .ZN(n326) );
  XNOR2_X1 U398 ( .A(KEYINPUT45), .B(n326), .ZN(n362) );
  XOR2_X1 U399 ( .A(G64GAT), .B(G92GAT), .Z(n328) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(G204GAT), .ZN(n327) );
  XNOR2_X1 U401 ( .A(n328), .B(n327), .ZN(n384) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XNOR2_X1 U403 ( .A(n384), .B(n442), .ZN(n332) );
  NAND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U405 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n333) );
  XNOR2_X1 U406 ( .A(n334), .B(n333), .ZN(n342) );
  XNOR2_X1 U407 ( .A(G106GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U408 ( .A(n335), .B(G148GAT), .ZN(n416) );
  XNOR2_X1 U409 ( .A(n416), .B(n336), .ZN(n340) );
  XOR2_X1 U410 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n338) );
  XNOR2_X1 U411 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n337) );
  XOR2_X1 U412 ( .A(n338), .B(n337), .Z(n339) );
  XOR2_X1 U413 ( .A(KEYINPUT68), .B(G22GAT), .Z(n344) );
  XNOR2_X1 U414 ( .A(G141GAT), .B(G197GAT), .ZN(n343) );
  XNOR2_X1 U415 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U416 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n346) );
  XNOR2_X1 U417 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n345) );
  XNOR2_X1 U418 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U419 ( .A(n348), .B(n347), .ZN(n360) );
  XOR2_X1 U420 ( .A(G113GAT), .B(G43GAT), .Z(n351) );
  XOR2_X1 U421 ( .A(G169GAT), .B(G8GAT), .Z(n376) );
  XNOR2_X1 U422 ( .A(n376), .B(n349), .ZN(n350) );
  XNOR2_X1 U423 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U424 ( .A(n352), .B(G36GAT), .Z(n358) );
  XOR2_X1 U425 ( .A(n353), .B(KEYINPUT67), .Z(n355) );
  NAND2_X1 U426 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U427 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U428 ( .A(n356), .B(G50GAT), .ZN(n357) );
  XNOR2_X1 U429 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U430 ( .A(n360), .B(n359), .Z(n551) );
  INV_X1 U431 ( .A(n551), .ZN(n573) );
  AND2_X1 U432 ( .A1(n576), .A2(n551), .ZN(n361) );
  AND2_X1 U433 ( .A1(n362), .A2(n361), .ZN(n369) );
  INV_X1 U434 ( .A(n544), .ZN(n563) );
  INV_X1 U435 ( .A(n560), .ZN(n581) );
  XNOR2_X1 U436 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n364) );
  XNOR2_X1 U437 ( .A(n576), .B(KEYINPUT41), .ZN(n553) );
  AND2_X1 U438 ( .A1(n573), .A2(n553), .ZN(n363) );
  XNOR2_X1 U439 ( .A(n364), .B(n363), .ZN(n365) );
  NOR2_X1 U440 ( .A1(n581), .A2(n365), .ZN(n366) );
  NAND2_X1 U441 ( .A1(n563), .A2(n366), .ZN(n367) );
  XNOR2_X1 U442 ( .A(n367), .B(KEYINPUT47), .ZN(n368) );
  NOR2_X1 U443 ( .A1(n369), .A2(n368), .ZN(n371) );
  XNOR2_X1 U444 ( .A(n371), .B(n370), .ZN(n532) );
  XOR2_X1 U445 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n373) );
  XNOR2_X1 U446 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n372) );
  XNOR2_X1 U447 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U448 ( .A(KEYINPUT19), .B(n374), .Z(n440) );
  XOR2_X1 U449 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n375) );
  XOR2_X1 U450 ( .A(n378), .B(KEYINPUT88), .Z(n380) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U452 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U453 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U454 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n383) );
  XNOR2_X1 U455 ( .A(n383), .B(G211GAT), .ZN(n427) );
  XNOR2_X1 U456 ( .A(n427), .B(n384), .ZN(n385) );
  XNOR2_X1 U457 ( .A(n524), .B(KEYINPUT120), .ZN(n387) );
  NOR2_X1 U458 ( .A1(n532), .A2(n387), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n412) );
  XOR2_X1 U460 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(G134GAT), .ZN(n391) );
  XNOR2_X1 U462 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U463 ( .A(G57GAT), .B(G148GAT), .Z(n394) );
  XNOR2_X1 U464 ( .A(G120GAT), .B(G155GAT), .ZN(n393) );
  XNOR2_X1 U465 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U466 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U467 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n398) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U469 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U470 ( .A(KEYINPUT87), .B(n399), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U472 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n403) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(KEYINPUT86), .ZN(n402) );
  XNOR2_X1 U474 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U475 ( .A(n405), .B(n404), .Z(n411) );
  XOR2_X1 U476 ( .A(G127GAT), .B(KEYINPUT0), .Z(n407) );
  XNOR2_X1 U477 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n406) );
  XNOR2_X1 U478 ( .A(n407), .B(n406), .ZN(n444) );
  XOR2_X1 U479 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n409) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n444), .B(n428), .ZN(n410) );
  XNOR2_X1 U483 ( .A(n411), .B(n410), .ZN(n521) );
  NAND2_X1 U484 ( .A1(n412), .A2(n521), .ZN(n413) );
  XNOR2_X1 U485 ( .A(n414), .B(n413), .ZN(n570) );
  XOR2_X1 U486 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U489 ( .A(n420), .B(n419), .Z(n422) );
  XNOR2_X1 U490 ( .A(G218GAT), .B(KEYINPUT22), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U492 ( .A(G204GAT), .B(KEYINPUT23), .Z(n424) );
  XNOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT84), .ZN(n423) );
  XNOR2_X1 U494 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U495 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U496 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U497 ( .A(n430), .B(n429), .ZN(n458) );
  NOR2_X1 U498 ( .A1(n570), .A2(n458), .ZN(n432) );
  INV_X1 U499 ( .A(KEYINPUT55), .ZN(n431) );
  XNOR2_X1 U500 ( .A(n432), .B(n431), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT82), .B(G176GAT), .Z(n434) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U503 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U504 ( .A(n435), .B(KEYINPUT20), .Z(n439) );
  XOR2_X1 U505 ( .A(G99GAT), .B(G190GAT), .Z(n437) );
  XNOR2_X1 U506 ( .A(G169GAT), .B(G15GAT), .ZN(n436) );
  XNOR2_X1 U507 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U508 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U510 ( .A(n447), .B(n446), .Z(n457) );
  INV_X1 U511 ( .A(n457), .ZN(n470) );
  NAND2_X1 U512 ( .A1(n448), .A2(n470), .ZN(n449) );
  XOR2_X1 U513 ( .A(KEYINPUT122), .B(n449), .Z(n566) );
  NAND2_X1 U514 ( .A1(n566), .A2(n544), .ZN(n452) );
  XOR2_X1 U515 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n450) );
  XOR2_X1 U516 ( .A(n458), .B(KEYINPUT28), .Z(n533) );
  NAND2_X1 U517 ( .A1(n573), .A2(n576), .ZN(n491) );
  NOR2_X1 U518 ( .A1(n524), .A2(n457), .ZN(n453) );
  XOR2_X1 U519 ( .A(KEYINPUT95), .B(n453), .Z(n454) );
  NOR2_X1 U520 ( .A1(n458), .A2(n454), .ZN(n456) );
  XOR2_X1 U521 ( .A(KEYINPUT93), .B(KEYINPUT26), .Z(n460) );
  NAND2_X1 U522 ( .A1(n458), .A2(n457), .ZN(n459) );
  XOR2_X1 U523 ( .A(n460), .B(n459), .Z(n549) );
  INV_X1 U524 ( .A(n549), .ZN(n571) );
  XOR2_X1 U525 ( .A(n524), .B(KEYINPUT27), .Z(n461) );
  XNOR2_X1 U526 ( .A(KEYINPUT91), .B(n461), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n571), .A2(n468), .ZN(n463) );
  NAND2_X1 U528 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n521), .A2(n466), .ZN(n467) );
  XOR2_X1 U530 ( .A(KEYINPUT97), .B(n467), .Z(n473) );
  NOR2_X1 U531 ( .A1(n521), .A2(n468), .ZN(n469) );
  XOR2_X1 U532 ( .A(KEYINPUT92), .B(n469), .Z(n531) );
  NOR2_X1 U533 ( .A1(n470), .A2(n531), .ZN(n471) );
  NAND2_X1 U534 ( .A1(n533), .A2(n471), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n473), .A2(n472), .ZN(n489) );
  NAND2_X1 U536 ( .A1(n560), .A2(n489), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n474), .A2(n584), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n491), .A2(n520), .ZN(n478) );
  NOR2_X1 U539 ( .A1(n533), .A2(n504), .ZN(n481) );
  NOR2_X1 U540 ( .A1(n524), .A2(n504), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1329GAT) );
  NAND2_X1 U542 ( .A1(n566), .A2(n553), .ZN(n487) );
  XOR2_X1 U543 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(G176GAT), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1349GAT) );
  NOR2_X1 U546 ( .A1(n544), .A2(n560), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT16), .ZN(n490) );
  NAND2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n510) );
  OR2_X1 U549 ( .A1(n491), .A2(n510), .ZN(n499) );
  NOR2_X1 U550 ( .A1(n521), .A2(n499), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT98), .B(KEYINPUT34), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U553 ( .A(G1GAT), .B(n494), .Z(G1324GAT) );
  NOR2_X1 U554 ( .A1(n524), .A2(n499), .ZN(n495) );
  XOR2_X1 U555 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  NOR2_X1 U556 ( .A1(n457), .A2(n499), .ZN(n497) );
  XNOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U559 ( .A(G15GAT), .B(n498), .Z(G1326GAT) );
  NOR2_X1 U560 ( .A1(n533), .A2(n499), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT100), .B(n500), .Z(n501) );
  XNOR2_X1 U562 ( .A(G22GAT), .B(n501), .ZN(G1327GAT) );
  NOR2_X1 U563 ( .A1(n504), .A2(n521), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n504), .A2(n457), .ZN(n506) );
  XNOR2_X1 U567 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n509) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n551), .A2(n553), .ZN(n519) );
  OR2_X1 U574 ( .A1(n519), .A2(n510), .ZN(n516) );
  NOR2_X1 U575 ( .A1(n521), .A2(n516), .ZN(n511) );
  XOR2_X1 U576 ( .A(n512), .B(n511), .Z(G1332GAT) );
  NOR2_X1 U577 ( .A1(n524), .A2(n516), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n457), .A2(n516), .ZN(n515) );
  XOR2_X1 U581 ( .A(G71GAT), .B(n515), .Z(G1334GAT) );
  NOR2_X1 U582 ( .A1(n533), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  OR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n521), .A2(n527), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT110), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n527), .ZN(n525) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n457), .A2(n527), .ZN(n526) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n533), .A2(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n550) );
  NAND2_X1 U598 ( .A1(n533), .A2(n550), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n457), .A2(n534), .ZN(n535) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(n535), .Z(n545) );
  NAND2_X1 U601 ( .A1(n545), .A2(n573), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT114), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U605 ( .A1(n545), .A2(n553), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n542) );
  NAND2_X1 U609 ( .A1(n545), .A2(n581), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n562) );
  NOR2_X1 U617 ( .A1(n551), .A2(n562), .ZN(n552) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  INV_X1 U619 ( .A(n553), .ZN(n554) );
  NOR2_X1 U620 ( .A1(n554), .A2(n562), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT52), .B(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n562), .ZN(n561) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n573), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n581), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n575) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(n572), .Z(n585) );
  INV_X1 U639 ( .A(n585), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n580), .A2(n573), .ZN(n574) );
  XOR2_X1 U641 ( .A(n575), .B(n574), .Z(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n578) );
  OR2_X1 U643 ( .A1(n585), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT127), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

