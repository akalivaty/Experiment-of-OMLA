

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746;

  XNOR2_X1 U368 ( .A(n384), .B(KEYINPUT0), .ZN(n592) );
  XNOR2_X1 U369 ( .A(n389), .B(KEYINPUT94), .ZN(n591) );
  XNOR2_X1 U370 ( .A(n429), .B(n428), .ZN(n369) );
  AND2_X2 U371 ( .A1(n410), .A2(n400), .ZN(n702) );
  AND2_X1 U372 ( .A1(n376), .A2(n377), .ZN(n346) );
  INV_X1 U373 ( .A(n537), .ZN(n670) );
  NOR2_X2 U374 ( .A1(n556), .A2(n442), .ZN(n384) );
  XNOR2_X2 U375 ( .A(n546), .B(KEYINPUT40), .ZN(n745) );
  NOR2_X1 U376 ( .A1(n673), .A2(n589), .ZN(n590) );
  XNOR2_X1 U377 ( .A(n398), .B(n397), .ZN(n576) );
  NOR2_X1 U378 ( .A1(n743), .A2(n584), .ZN(n586) );
  XNOR2_X1 U379 ( .A(n380), .B(KEYINPUT35), .ZN(n743) );
  NAND2_X1 U380 ( .A1(n512), .A2(n576), .ZN(n585) );
  NAND2_X1 U381 ( .A1(n347), .A2(n364), .ZN(n380) );
  XNOR2_X1 U382 ( .A(n382), .B(KEYINPUT42), .ZN(n746) );
  INV_X1 U383 ( .A(n589), .ZN(n371) );
  XNOR2_X1 U384 ( .A(n563), .B(n436), .ZN(n556) );
  XNOR2_X1 U385 ( .A(n496), .B(n495), .ZN(n537) );
  XOR2_X1 U386 ( .A(n692), .B(KEYINPUT59), .Z(n693) );
  XNOR2_X1 U387 ( .A(G104), .B(G110), .ZN(n420) );
  XNOR2_X1 U388 ( .A(n424), .B(n367), .ZN(n492) );
  XNOR2_X1 U389 ( .A(KEYINPUT3), .B(G119), .ZN(n424) );
  XNOR2_X1 U390 ( .A(n368), .B(G116), .ZN(n367) );
  INV_X1 U391 ( .A(G113), .ZN(n368) );
  XOR2_X1 U392 ( .A(G137), .B(KEYINPUT71), .Z(n725) );
  INV_X1 U393 ( .A(KEYINPUT76), .ZN(n421) );
  NAND2_X1 U394 ( .A1(n589), .A2(KEYINPUT34), .ZN(n366) );
  INV_X1 U395 ( .A(G234), .ZN(n395) );
  XOR2_X1 U396 ( .A(G146), .B(G125), .Z(n443) );
  NOR2_X1 U397 ( .A1(n375), .A2(n373), .ZN(n569) );
  INV_X1 U398 ( .A(n548), .ZN(n387) );
  AND2_X1 U399 ( .A1(n510), .A2(G221), .ZN(n388) );
  INV_X1 U400 ( .A(KEYINPUT66), .ZN(n428) );
  XNOR2_X1 U401 ( .A(G143), .B(G128), .ZN(n459) );
  XNOR2_X1 U402 ( .A(n443), .B(KEYINPUT10), .ZN(n500) );
  XOR2_X1 U403 ( .A(KEYINPUT72), .B(G134), .Z(n726) );
  XNOR2_X1 U404 ( .A(n492), .B(n490), .ZN(n386) );
  XNOR2_X1 U405 ( .A(n492), .B(n427), .ZN(n714) );
  INV_X1 U406 ( .A(KEYINPUT80), .ZN(n425) );
  XNOR2_X1 U407 ( .A(KEYINPUT16), .B(G122), .ZN(n426) );
  XNOR2_X1 U408 ( .A(n504), .B(n415), .ZN(n505) );
  XNOR2_X1 U409 ( .A(G119), .B(G110), .ZN(n502) );
  XNOR2_X1 U410 ( .A(G113), .B(G122), .ZN(n444) );
  XOR2_X1 U411 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n448) );
  XNOR2_X1 U412 ( .A(G143), .B(G104), .ZN(n450) );
  XNOR2_X1 U413 ( .A(n500), .B(n477), .ZN(n724) );
  XNOR2_X1 U414 ( .A(KEYINPUT15), .B(G902), .ZN(n614) );
  NAND2_X1 U415 ( .A1(n371), .A2(n372), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n561), .B(n381), .ZN(n582) );
  INV_X1 U417 ( .A(KEYINPUT90), .ZN(n381) );
  INV_X1 U418 ( .A(KEYINPUT105), .ZN(n536) );
  INV_X1 U419 ( .A(KEYINPUT108), .ZN(n531) );
  XNOR2_X1 U420 ( .A(n457), .B(n456), .ZN(n580) );
  XNOR2_X1 U421 ( .A(n511), .B(KEYINPUT25), .ZN(n397) );
  NAND2_X1 U422 ( .A1(n399), .A2(n494), .ZN(n398) );
  INV_X1 U423 ( .A(n614), .ZN(n400) );
  XNOR2_X1 U424 ( .A(n476), .B(n475), .ZN(n478) );
  INV_X1 U425 ( .A(G237), .ZN(n433) );
  XOR2_X1 U426 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n488) );
  XOR2_X1 U427 ( .A(KEYINPUT75), .B(KEYINPUT24), .Z(n503) );
  NAND2_X1 U428 ( .A1(n348), .A2(n392), .ZN(n501) );
  NAND2_X1 U429 ( .A1(n732), .A2(n393), .ZN(n392) );
  NOR2_X1 U430 ( .A1(n462), .A2(n395), .ZN(n393) );
  XNOR2_X1 U431 ( .A(KEYINPUT86), .B(KEYINPUT48), .ZN(n570) );
  INV_X1 U432 ( .A(KEYINPUT73), .ZN(n383) );
  AND2_X1 U433 ( .A1(n666), .A2(n387), .ZN(n519) );
  XNOR2_X1 U434 ( .A(n441), .B(KEYINPUT92), .ZN(n442) );
  INV_X1 U435 ( .A(G953), .ZN(n707) );
  XOR2_X1 U436 ( .A(G122), .B(G116), .Z(n464) );
  XOR2_X1 U437 ( .A(G107), .B(G134), .Z(n458) );
  XNOR2_X1 U438 ( .A(n474), .B(n725), .ZN(n475) );
  XNOR2_X1 U439 ( .A(n480), .B(n479), .ZN(n493) );
  XNOR2_X1 U440 ( .A(n431), .B(n432), .ZN(n624) );
  XNOR2_X1 U441 ( .A(n480), .B(n714), .ZN(n431) );
  XNOR2_X1 U442 ( .A(n543), .B(KEYINPUT39), .ZN(n544) );
  NAND2_X1 U443 ( .A1(n435), .A2(n652), .ZN(n563) );
  NAND2_X1 U444 ( .A1(n535), .A2(n390), .ZN(n389) );
  NOR2_X1 U445 ( .A1(n576), .A2(n391), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n509), .B(n508), .ZN(n703) );
  XNOR2_X1 U447 ( .A(n453), .B(n452), .ZN(n692) );
  INV_X1 U448 ( .A(G210), .ZN(n409) );
  NOR2_X1 U449 ( .A1(n557), .A2(n684), .ZN(n382) );
  OR2_X1 U450 ( .A1(n365), .A2(n685), .ZN(n364) );
  XNOR2_X1 U451 ( .A(n361), .B(KEYINPUT32), .ZN(n744) );
  NOR2_X1 U452 ( .A1(n582), .A2(n363), .ZN(n362) );
  NAND2_X1 U453 ( .A1(n583), .A2(n576), .ZN(n363) );
  XNOR2_X1 U454 ( .A(n691), .B(n690), .ZN(n385) );
  AND2_X1 U455 ( .A1(n370), .A2(n355), .ZN(n347) );
  XNOR2_X1 U456 ( .A(n388), .B(KEYINPUT21), .ZN(n666) );
  INV_X1 U457 ( .A(n666), .ZN(n391) );
  AND2_X1 U458 ( .A1(n396), .A2(n394), .ZN(n348) );
  XOR2_X1 U459 ( .A(n491), .B(n386), .Z(n349) );
  AND2_X1 U460 ( .A1(n378), .A2(n377), .ZN(n350) );
  OR2_X1 U461 ( .A1(n687), .A2(n686), .ZN(n351) );
  INV_X1 U462 ( .A(n576), .ZN(n667) );
  AND2_X1 U463 ( .A1(n405), .A2(n404), .ZN(n352) );
  OR2_X1 U464 ( .A1(n542), .A2(n548), .ZN(n353) );
  AND2_X1 U465 ( .A1(n434), .A2(G210), .ZN(n354) );
  AND2_X1 U466 ( .A1(n366), .A2(n581), .ZN(n355) );
  XOR2_X1 U467 ( .A(KEYINPUT74), .B(G469), .Z(n356) );
  XOR2_X1 U468 ( .A(n578), .B(n577), .Z(n357) );
  INV_X1 U469 ( .A(KEYINPUT34), .ZN(n372) );
  XOR2_X1 U470 ( .A(n624), .B(n623), .Z(n358) );
  XNOR2_X1 U471 ( .A(KEYINPUT62), .B(n615), .ZN(n359) );
  INV_X1 U472 ( .A(n547), .ZN(n407) );
  NOR2_X1 U473 ( .A1(n614), .A2(n456), .ZN(n360) );
  AND2_X1 U474 ( .A1(n618), .A2(n617), .ZN(n706) );
  INV_X1 U475 ( .A(n706), .ZN(n377) );
  NAND2_X1 U476 ( .A1(n403), .A2(n547), .ZN(n374) );
  INV_X1 U477 ( .A(n703), .ZN(n399) );
  XNOR2_X1 U478 ( .A(n505), .B(n506), .ZN(n509) );
  XNOR2_X1 U479 ( .A(n520), .B(n383), .ZN(n527) );
  NAND2_X1 U480 ( .A1(n600), .A2(n362), .ZN(n361) );
  XNOR2_X2 U481 ( .A(n379), .B(n357), .ZN(n685) );
  XNOR2_X2 U482 ( .A(n730), .B(n430), .ZN(n480) );
  XNOR2_X2 U483 ( .A(n369), .B(n459), .ZN(n730) );
  NAND2_X1 U484 ( .A1(n685), .A2(KEYINPUT34), .ZN(n370) );
  NOR2_X1 U485 ( .A1(n374), .A2(n745), .ZN(n373) );
  NAND2_X1 U486 ( .A1(n352), .A2(n406), .ZN(n375) );
  XNOR2_X1 U487 ( .A(n591), .B(n536), .ZN(n541) );
  NAND2_X1 U488 ( .A1(n624), .A2(n614), .ZN(n401) );
  XNOR2_X1 U489 ( .A(n616), .B(n359), .ZN(n376) );
  XNOR2_X1 U490 ( .A(n625), .B(n358), .ZN(n378) );
  NOR2_X1 U491 ( .A1(n540), .A2(n353), .ZN(n412) );
  NAND2_X1 U492 ( .A1(n471), .A2(n592), .ZN(n473) );
  NAND2_X1 U493 ( .A1(n585), .A2(n586), .ZN(n587) );
  NOR2_X1 U494 ( .A1(n572), .A2(n644), .ZN(n546) );
  NAND2_X1 U495 ( .A1(n588), .A2(n597), .ZN(n379) );
  NOR2_X2 U496 ( .A1(n664), .A2(n663), .ZN(n588) );
  NOR2_X1 U497 ( .A1(n527), .A2(n537), .ZN(n529) );
  NOR2_X1 U498 ( .A1(n385), .A2(n706), .ZN(G54) );
  INV_X1 U499 ( .A(n618), .ZN(n732) );
  NAND2_X1 U500 ( .A1(n462), .A2(n395), .ZN(n394) );
  NAND2_X1 U501 ( .A1(n618), .A2(n462), .ZN(n396) );
  XNOR2_X2 U502 ( .A(G953), .B(KEYINPUT64), .ZN(n618) );
  NAND2_X1 U503 ( .A1(n410), .A2(n360), .ZN(n694) );
  NAND2_X1 U504 ( .A1(n410), .A2(n411), .ZN(n616) );
  NOR2_X1 U505 ( .A1(n410), .A2(n351), .ZN(n688) );
  AND2_X2 U506 ( .A1(n613), .A2(n612), .ZN(n410) );
  INV_X1 U507 ( .A(n435), .ZN(n551) );
  XNOR2_X2 U508 ( .A(n401), .B(n354), .ZN(n435) );
  INV_X1 U509 ( .A(n592), .ZN(n589) );
  XNOR2_X2 U510 ( .A(n534), .B(KEYINPUT1), .ZN(n663) );
  NAND2_X1 U511 ( .A1(n410), .A2(n408), .ZN(n625) );
  XNOR2_X2 U512 ( .A(n605), .B(n604), .ZN(n708) );
  OR2_X2 U513 ( .A1(n402), .A2(G902), .ZN(n484) );
  XNOR2_X1 U514 ( .A(n402), .B(n689), .ZN(n690) );
  XNOR2_X1 U515 ( .A(n482), .B(n483), .ZN(n402) );
  INV_X1 U516 ( .A(n746), .ZN(n403) );
  INV_X1 U517 ( .A(n555), .ZN(n404) );
  NAND2_X1 U518 ( .A1(n746), .A2(n407), .ZN(n405) );
  NAND2_X1 U519 ( .A1(n745), .A2(n407), .ZN(n406) );
  NOR2_X1 U520 ( .A1(n614), .A2(n409), .ZN(n408) );
  NOR2_X1 U521 ( .A1(n614), .A2(n495), .ZN(n411) );
  NOR2_X1 U522 ( .A1(n541), .A2(n540), .ZN(n414) );
  NAND2_X1 U523 ( .A1(n413), .A2(n412), .ZN(n545) );
  INV_X1 U524 ( .A(n541), .ZN(n413) );
  NAND2_X1 U525 ( .A1(n414), .A2(n553), .ZN(n554) );
  NOR2_X1 U526 ( .A1(n609), .A2(n575), .ZN(n606) );
  XNOR2_X1 U527 ( .A(n571), .B(n570), .ZN(n609) );
  XNOR2_X2 U528 ( .A(n473), .B(n472), .ZN(n600) );
  XOR2_X1 U529 ( .A(n503), .B(n502), .Z(n415) );
  INV_X1 U530 ( .A(KEYINPUT8), .ZN(n462) );
  INV_X1 U531 ( .A(KEYINPUT104), .ZN(n577) );
  INV_X1 U532 ( .A(KEYINPUT28), .ZN(n528) );
  INV_X1 U533 ( .A(KEYINPUT82), .ZN(n481) );
  INV_X1 U534 ( .A(KEYINPUT45), .ZN(n604) );
  XNOR2_X1 U535 ( .A(n532), .B(n531), .ZN(n557) );
  XNOR2_X1 U536 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U537 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U538 ( .A(n443), .B(KEYINPUT18), .Z(n419) );
  INV_X1 U539 ( .A(G224), .ZN(n416) );
  OR2_X1 U540 ( .A1(n618), .A2(n416), .ZN(n417) );
  XNOR2_X1 U541 ( .A(n417), .B(KEYINPUT17), .ZN(n418) );
  XNOR2_X1 U542 ( .A(n419), .B(n418), .ZN(n423) );
  XNOR2_X1 U543 ( .A(n420), .B(G107), .ZN(n715) );
  XNOR2_X1 U544 ( .A(n421), .B(KEYINPUT77), .ZN(n422) );
  XNOR2_X1 U545 ( .A(n715), .B(n422), .ZN(n476) );
  XNOR2_X1 U546 ( .A(n423), .B(n476), .ZN(n432) );
  XNOR2_X1 U547 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X2 U548 ( .A(KEYINPUT70), .B(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U549 ( .A(KEYINPUT68), .B(G101), .ZN(n430) );
  INV_X1 U550 ( .A(G902), .ZN(n494) );
  NAND2_X1 U551 ( .A1(n494), .A2(n433), .ZN(n434) );
  NAND2_X1 U552 ( .A1(n434), .A2(G214), .ZN(n652) );
  INV_X1 U553 ( .A(KEYINPUT19), .ZN(n436) );
  NAND2_X1 U554 ( .A1(G234), .A2(G237), .ZN(n437) );
  XNOR2_X1 U555 ( .A(n437), .B(KEYINPUT14), .ZN(n438) );
  AND2_X1 U556 ( .A1(G952), .A2(n438), .ZN(n680) );
  NAND2_X1 U557 ( .A1(n680), .A2(n707), .ZN(n514) );
  NAND2_X1 U558 ( .A1(n438), .A2(G902), .ZN(n439) );
  XNOR2_X1 U559 ( .A(n439), .B(KEYINPUT91), .ZN(n515) );
  NOR2_X1 U560 ( .A1(G898), .A2(n707), .ZN(n718) );
  NAND2_X1 U561 ( .A1(n515), .A2(n718), .ZN(n440) );
  AND2_X1 U562 ( .A1(n514), .A2(n440), .ZN(n441) );
  XNOR2_X1 U563 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n455) );
  XOR2_X1 U564 ( .A(G131), .B(G140), .Z(n477) );
  XOR2_X1 U565 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n445) );
  XNOR2_X1 U566 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U567 ( .A(n724), .B(n446), .ZN(n453) );
  NOR2_X1 U568 ( .A1(G953), .A2(G237), .ZN(n486) );
  NAND2_X1 U569 ( .A1(G214), .A2(n486), .ZN(n447) );
  XNOR2_X1 U570 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U571 ( .A(n449), .B(KEYINPUT11), .Z(n451) );
  XNOR2_X1 U572 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U573 ( .A1(G902), .A2(n692), .ZN(n454) );
  XNOR2_X1 U574 ( .A(n455), .B(n454), .ZN(n457) );
  INV_X1 U575 ( .A(G475), .ZN(n456) );
  XNOR2_X1 U576 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n461) );
  XNOR2_X1 U577 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U578 ( .A(n461), .B(n460), .ZN(n466) );
  NAND2_X1 U579 ( .A1(G217), .A2(n501), .ZN(n463) );
  XNOR2_X1 U580 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U581 ( .A(n466), .B(n465), .ZN(n698) );
  NOR2_X1 U582 ( .A1(G902), .A2(n698), .ZN(n468) );
  INV_X1 U583 ( .A(G478), .ZN(n467) );
  XNOR2_X1 U584 ( .A(n468), .B(n467), .ZN(n558) );
  INV_X1 U585 ( .A(n558), .ZN(n579) );
  NAND2_X1 U586 ( .A1(n580), .A2(n579), .ZN(n656) );
  XOR2_X1 U587 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n470) );
  NAND2_X1 U588 ( .A1(G234), .A2(n614), .ZN(n469) );
  XNOR2_X1 U589 ( .A(n470), .B(n469), .ZN(n510) );
  NOR2_X1 U590 ( .A1(n656), .A2(n391), .ZN(n471) );
  XNOR2_X1 U591 ( .A(KEYINPUT79), .B(KEYINPUT22), .ZN(n472) );
  NAND2_X1 U592 ( .A1(G227), .A2(n732), .ZN(n474) );
  XOR2_X1 U593 ( .A(n478), .B(n477), .Z(n483) );
  XNOR2_X1 U594 ( .A(n726), .B(G146), .ZN(n479) );
  XNOR2_X1 U595 ( .A(n493), .B(n481), .ZN(n482) );
  XNOR2_X2 U596 ( .A(n484), .B(n356), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n600), .A2(n663), .ZN(n485) );
  XNOR2_X1 U598 ( .A(n485), .B(KEYINPUT103), .ZN(n497) );
  NAND2_X1 U599 ( .A1(n486), .A2(G210), .ZN(n487) );
  XNOR2_X1 U600 ( .A(n487), .B(n488), .ZN(n489) );
  XOR2_X1 U601 ( .A(n489), .B(KEYINPUT95), .Z(n491) );
  XNOR2_X1 U602 ( .A(G137), .B(G131), .ZN(n490) );
  XNOR2_X1 U603 ( .A(n493), .B(n349), .ZN(n615) );
  NAND2_X1 U604 ( .A1(n615), .A2(n494), .ZN(n496) );
  INV_X1 U605 ( .A(G472), .ZN(n495) );
  NAND2_X1 U606 ( .A1(n497), .A2(n537), .ZN(n498) );
  XNOR2_X1 U607 ( .A(n498), .B(KEYINPUT67), .ZN(n512) );
  XNOR2_X1 U608 ( .A(KEYINPUT23), .B(KEYINPUT81), .ZN(n499) );
  XOR2_X1 U609 ( .A(n500), .B(n499), .Z(n506) );
  NAND2_X1 U610 ( .A1(G221), .A2(n501), .ZN(n504) );
  XNOR2_X1 U611 ( .A(G128), .B(G140), .ZN(n507) );
  XNOR2_X1 U612 ( .A(n507), .B(n725), .ZN(n508) );
  NAND2_X1 U613 ( .A1(G217), .A2(n510), .ZN(n511) );
  XNOR2_X1 U614 ( .A(n585), .B(G110), .ZN(G12) );
  INV_X1 U615 ( .A(n663), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n580), .A2(n558), .ZN(n513) );
  XOR2_X1 U617 ( .A(n513), .B(KEYINPUT101), .Z(n640) );
  INV_X1 U618 ( .A(n640), .ZN(n644) );
  INV_X1 U619 ( .A(n514), .ZN(n518) );
  NAND2_X1 U620 ( .A1(n618), .A2(n515), .ZN(n516) );
  NOR2_X1 U621 ( .A1(G900), .A2(n516), .ZN(n517) );
  NOR2_X1 U622 ( .A1(n518), .A2(n517), .ZN(n548) );
  NAND2_X1 U623 ( .A1(n576), .A2(n519), .ZN(n520) );
  INV_X1 U624 ( .A(KEYINPUT6), .ZN(n521) );
  XNOR2_X1 U625 ( .A(n537), .B(n521), .ZN(n583) );
  OR2_X1 U626 ( .A1(n527), .A2(n583), .ZN(n522) );
  NOR2_X1 U627 ( .A1(n644), .A2(n522), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n562), .A2(n652), .ZN(n523) );
  NOR2_X1 U629 ( .A1(n561), .A2(n523), .ZN(n524) );
  XNOR2_X1 U630 ( .A(n524), .B(KEYINPUT43), .ZN(n526) );
  INV_X1 U631 ( .A(n551), .ZN(n525) );
  OR2_X1 U632 ( .A1(n526), .A2(n525), .ZN(n574) );
  XNOR2_X1 U633 ( .A(n574), .B(G140), .ZN(G42) );
  XNOR2_X1 U634 ( .A(n529), .B(n528), .ZN(n530) );
  NOR2_X1 U635 ( .A1(n534), .A2(n530), .ZN(n532) );
  XOR2_X1 U636 ( .A(KEYINPUT38), .B(n551), .Z(n542) );
  INV_X1 U637 ( .A(n542), .ZN(n653) );
  NAND2_X1 U638 ( .A1(n653), .A2(n652), .ZN(n657) );
  NOR2_X1 U639 ( .A1(n656), .A2(n657), .ZN(n533) );
  XNOR2_X1 U640 ( .A(n533), .B(KEYINPUT41), .ZN(n684) );
  INV_X1 U641 ( .A(n534), .ZN(n535) );
  NAND2_X1 U642 ( .A1(n652), .A2(n670), .ZN(n538) );
  XNOR2_X1 U643 ( .A(n538), .B(KEYINPUT30), .ZN(n539) );
  XNOR2_X1 U644 ( .A(KEYINPUT106), .B(n539), .ZN(n540) );
  INV_X1 U645 ( .A(KEYINPUT78), .ZN(n543) );
  XNOR2_X1 U646 ( .A(n545), .B(n544), .ZN(n572) );
  XNOR2_X1 U647 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n547) );
  INV_X1 U648 ( .A(n580), .ZN(n550) );
  NOR2_X1 U649 ( .A1(n579), .A2(n548), .ZN(n549) );
  NAND2_X1 U650 ( .A1(n550), .A2(n549), .ZN(n552) );
  NOR2_X1 U651 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U652 ( .A(KEYINPUT107), .B(n554), .ZN(n741) );
  XNOR2_X1 U653 ( .A(n741), .B(KEYINPUT84), .ZN(n555) );
  NOR2_X1 U654 ( .A1(n557), .A2(n556), .ZN(n641) );
  AND2_X1 U655 ( .A1(n580), .A2(n558), .ZN(n636) );
  NOR2_X1 U656 ( .A1(n636), .A2(n640), .ZN(n658) );
  NOR2_X1 U657 ( .A1(KEYINPUT69), .A2(n658), .ZN(n559) );
  NAND2_X1 U658 ( .A1(n641), .A2(n559), .ZN(n560) );
  XNOR2_X1 U659 ( .A(KEYINPUT47), .B(n560), .ZN(n567) );
  INV_X1 U660 ( .A(n562), .ZN(n564) );
  NOR2_X1 U661 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U662 ( .A(KEYINPUT36), .B(n565), .Z(n566) );
  NOR2_X1 U663 ( .A1(n582), .A2(n566), .ZN(n650) );
  NOR2_X1 U664 ( .A1(n567), .A2(n650), .ZN(n568) );
  NAND2_X1 U665 ( .A1(n569), .A2(n568), .ZN(n571) );
  INV_X1 U666 ( .A(n636), .ZN(n648) );
  NOR2_X1 U667 ( .A1(n648), .A2(n572), .ZN(n573) );
  XNOR2_X1 U668 ( .A(n573), .B(KEYINPUT109), .ZN(n742) );
  NAND2_X1 U669 ( .A1(n742), .A2(n574), .ZN(n608) );
  OR2_X1 U670 ( .A1(KEYINPUT85), .A2(n608), .ZN(n575) );
  INV_X1 U671 ( .A(n583), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n667), .A2(n666), .ZN(n664) );
  XNOR2_X1 U673 ( .A(KEYINPUT33), .B(KEYINPUT89), .ZN(n578) );
  NOR2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U675 ( .A(n744), .ZN(n584) );
  XNOR2_X1 U676 ( .A(n587), .B(KEYINPUT44), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n588), .A2(n670), .ZN(n673) );
  XNOR2_X1 U678 ( .A(n590), .B(KEYINPUT31), .ZN(n647) );
  NOR2_X1 U679 ( .A1(n591), .A2(n670), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n593), .A2(n371), .ZN(n630) );
  NAND2_X1 U681 ( .A1(n647), .A2(n630), .ZN(n595) );
  INV_X1 U682 ( .A(n658), .ZN(n594) );
  NAND2_X1 U683 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U684 ( .A(KEYINPUT102), .B(n596), .Z(n601) );
  NAND2_X1 U685 ( .A1(n663), .A2(n667), .ZN(n598) );
  NOR2_X1 U686 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n627) );
  OR2_X1 U688 ( .A1(n601), .A2(n627), .ZN(n602) );
  NOR2_X2 U689 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n708), .ZN(n607) );
  XNOR2_X1 U691 ( .A(n607), .B(KEYINPUT2), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n723) );
  INV_X1 U693 ( .A(KEYINPUT85), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n723), .A2(n610), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n708), .A2(n611), .ZN(n612) );
  INV_X1 U696 ( .A(G952), .ZN(n617) );
  XNOR2_X1 U697 ( .A(KEYINPUT110), .B(KEYINPUT63), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT87), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n346), .B(n620), .ZN(G57) );
  XOR2_X1 U700 ( .A(KEYINPUT88), .B(KEYINPUT54), .Z(n622) );
  XNOR2_X1 U701 ( .A(KEYINPUT55), .B(KEYINPUT83), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U703 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n350), .B(n626), .ZN(G51) );
  XNOR2_X1 U705 ( .A(G101), .B(n627), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT111), .ZN(G3) );
  NOR2_X1 U707 ( .A1(n644), .A2(n630), .ZN(n629) );
  XOR2_X1 U708 ( .A(G104), .B(n629), .Z(G6) );
  NOR2_X1 U709 ( .A1(n648), .A2(n630), .ZN(n635) );
  XOR2_X1 U710 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n632) );
  XNOR2_X1 U711 ( .A(G107), .B(KEYINPUT26), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U713 ( .A(KEYINPUT112), .B(n633), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n635), .B(n634), .ZN(G9) );
  XOR2_X1 U715 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n638) );
  NAND2_X1 U716 ( .A1(n641), .A2(n636), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U718 ( .A(G128), .B(n639), .ZN(G30) );
  XOR2_X1 U719 ( .A(G146), .B(KEYINPUT115), .Z(n643) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n643), .B(n642), .ZN(G48) );
  NOR2_X1 U722 ( .A1(n644), .A2(n647), .ZN(n645) );
  XOR2_X1 U723 ( .A(KEYINPUT116), .B(n645), .Z(n646) );
  XNOR2_X1 U724 ( .A(G113), .B(n646), .ZN(G15) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U726 ( .A(G116), .B(n649), .Z(G18) );
  XNOR2_X1 U727 ( .A(G125), .B(n650), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n651), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT117), .B(n654), .Z(n655) );
  NOR2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n660) );
  NOR2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(KEYINPUT118), .ZN(n662) );
  NOR2_X1 U735 ( .A1(n685), .A2(n662), .ZN(n678) );
  NAND2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(KEYINPUT50), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U739 ( .A(KEYINPUT49), .B(n668), .Z(n669) );
  NOR2_X1 U740 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(KEYINPUT51), .B(n675), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n684), .A2(n676), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U746 ( .A(KEYINPUT52), .B(n679), .Z(n681) );
  NAND2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U748 ( .A(KEYINPUT119), .B(n682), .ZN(n683) );
  OR2_X1 U749 ( .A1(G953), .A2(n683), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U751 ( .A(KEYINPUT53), .B(n688), .ZN(G75) );
  NAND2_X1 U752 ( .A1(n702), .A2(G469), .ZN(n691) );
  XOR2_X1 U753 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n689) );
  XNOR2_X1 U754 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X2 U755 ( .A1(n695), .A2(n706), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n696), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U757 ( .A1(n702), .A2(G478), .ZN(n700) );
  INV_X1 U758 ( .A(KEYINPUT121), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n706), .A2(n701), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n702), .A2(G217), .ZN(n704) );
  XNOR2_X1 U761 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U762 ( .A1(n706), .A2(n705), .ZN(G66) );
  NAND2_X1 U763 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U764 ( .A1(G953), .A2(G224), .ZN(n709) );
  XNOR2_X1 U765 ( .A(KEYINPUT61), .B(n709), .ZN(n710) );
  NAND2_X1 U766 ( .A1(n710), .A2(G898), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT122), .ZN(n712) );
  NAND2_X1 U768 ( .A1(n713), .A2(n712), .ZN(n722) );
  XOR2_X1 U769 ( .A(KEYINPUT123), .B(n714), .Z(n717) );
  XNOR2_X1 U770 ( .A(G101), .B(n715), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n720), .B(KEYINPUT124), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n722), .B(n721), .ZN(G69) );
  INV_X1 U775 ( .A(n723), .ZN(n731) );
  XOR2_X1 U776 ( .A(KEYINPUT125), .B(n724), .Z(n728) );
  XNOR2_X1 U777 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(n729) );
  XOR2_X1 U779 ( .A(n730), .B(n729), .Z(n735) );
  XNOR2_X1 U780 ( .A(n731), .B(n735), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U782 ( .A(KEYINPUT126), .B(n734), .ZN(n740) );
  XNOR2_X1 U783 ( .A(n735), .B(G227), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U785 ( .A1(G953), .A2(n737), .ZN(n738) );
  XOR2_X1 U786 ( .A(KEYINPUT127), .B(n738), .Z(n739) );
  NAND2_X1 U787 ( .A1(n740), .A2(n739), .ZN(G72) );
  XOR2_X1 U788 ( .A(n741), .B(G143), .Z(G45) );
  XNOR2_X1 U789 ( .A(G134), .B(n742), .ZN(G36) );
  XOR2_X1 U790 ( .A(n743), .B(G122), .Z(G24) );
  XNOR2_X1 U791 ( .A(G119), .B(n744), .ZN(G21) );
  XOR2_X1 U792 ( .A(n745), .B(G131), .Z(G33) );
  XOR2_X1 U793 ( .A(n746), .B(G137), .Z(G39) );
endmodule

