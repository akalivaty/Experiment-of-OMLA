

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802;

  OR2_X1 U371 ( .A1(n657), .A2(n724), .ZN(n606) );
  XNOR2_X1 U372 ( .A(n635), .B(KEYINPUT39), .ZN(n656) );
  AND2_X2 U373 ( .A1(n398), .A2(n663), .ZN(n390) );
  NAND2_X4 U374 ( .A1(n662), .A2(KEYINPUT65), .ZN(n397) );
  XOR2_X2 U375 ( .A(n404), .B(n683), .Z(n360) );
  XNOR2_X1 U376 ( .A(G146), .B(G125), .ZN(n457) );
  INV_X1 U377 ( .A(G902), .ZN(n367) );
  XNOR2_X1 U378 ( .A(n613), .B(n612), .ZN(n741) );
  NOR2_X1 U379 ( .A1(n757), .A2(n436), .ZN(n435) );
  AND2_X2 U380 ( .A1(n448), .A2(n450), .ZN(n447) );
  OR2_X2 U381 ( .A1(n597), .A2(n744), .ZN(n599) );
  NAND2_X2 U382 ( .A1(n428), .A2(n427), .ZN(n426) );
  INV_X2 U383 ( .A(n579), .ZN(n603) );
  AND2_X2 U384 ( .A1(n626), .A2(n690), .ZN(n402) );
  XNOR2_X2 U385 ( .A(n381), .B(KEYINPUT48), .ZN(n655) );
  XNOR2_X1 U386 ( .A(n422), .B(n499), .ZN(n517) );
  AND2_X1 U387 ( .A1(n800), .A2(n625), .ZN(n626) );
  XNOR2_X1 U388 ( .A(n604), .B(n401), .ZN(n727) );
  XNOR2_X1 U389 ( .A(n747), .B(n559), .ZN(n620) );
  INV_X1 U390 ( .A(n591), .ZN(n560) );
  XNOR2_X1 U391 ( .A(n510), .B(n509), .ZN(n558) );
  XNOR2_X1 U392 ( .A(n477), .B(n476), .ZN(n591) );
  AND2_X1 U393 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U394 ( .A(n423), .B(n517), .ZN(n785) );
  XNOR2_X1 U395 ( .A(n388), .B(G119), .ZN(n422) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n528) );
  INV_X1 U397 ( .A(KEYINPUT80), .ZN(n411) );
  INV_X2 U398 ( .A(G953), .ZN(n387) );
  XNOR2_X2 U399 ( .A(n406), .B(n407), .ZN(n405) );
  XNOR2_X1 U400 ( .A(n406), .B(n407), .ZN(n634) );
  NOR2_X1 U401 ( .A1(n393), .A2(n392), .ZN(n391) );
  NOR2_X1 U402 ( .A1(n399), .A2(n397), .ZN(n392) );
  BUF_X2 U403 ( .A(n558), .Z(n747) );
  XNOR2_X2 U404 ( .A(n589), .B(KEYINPUT110), .ZN(n607) );
  NAND2_X1 U405 ( .A1(n801), .A2(n379), .ZN(n377) );
  NAND2_X1 U406 ( .A1(n802), .A2(n379), .ZN(n378) );
  NAND2_X1 U407 ( .A1(n376), .A2(n375), .ZN(n374) );
  NOR2_X1 U408 ( .A1(n730), .A2(n653), .ZN(n384) );
  NAND2_X2 U409 ( .A1(n369), .A2(n365), .ZN(n641) );
  OR2_X1 U410 ( .A1(n704), .A2(n366), .ZN(n365) );
  NAND2_X1 U411 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U412 ( .A1(n661), .A2(n663), .ZN(n394) );
  INV_X1 U413 ( .A(KEYINPUT92), .ZN(n498) );
  NAND2_X1 U414 ( .A1(n568), .A2(n432), .ZN(n430) );
  NOR2_X1 U415 ( .A1(n568), .A2(n432), .ZN(n427) );
  XNOR2_X1 U416 ( .A(n641), .B(n563), .ZN(n597) );
  XNOR2_X1 U417 ( .A(n638), .B(KEYINPUT28), .ZN(n639) );
  XNOR2_X1 U418 ( .A(n792), .B(n492), .ZN(n704) );
  AND2_X1 U419 ( .A1(n386), .A2(G953), .ZN(n680) );
  INV_X1 U420 ( .A(G952), .ZN(n386) );
  INV_X1 U421 ( .A(KEYINPUT46), .ZN(n379) );
  XNOR2_X1 U422 ( .A(KEYINPUT91), .B(KEYINPUT15), .ZN(n470) );
  INV_X1 U423 ( .A(G237), .ZN(n497) );
  NAND2_X1 U424 ( .A1(n704), .A2(n494), .ZN(n371) );
  INV_X1 U425 ( .A(KEYINPUT86), .ZN(n432) );
  XNOR2_X1 U426 ( .A(G101), .B(G146), .ZN(n500) );
  XOR2_X1 U427 ( .A(KEYINPUT73), .B(G137), .Z(n501) );
  XOR2_X1 U428 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n503) );
  OR2_X1 U429 ( .A1(n654), .A2(n439), .ZN(n438) );
  INV_X1 U430 ( .A(n732), .ZN(n439) );
  NAND2_X1 U431 ( .A1(n547), .A2(G221), .ZN(n437) );
  XNOR2_X1 U432 ( .A(G122), .B(KEYINPUT98), .ZN(n526) );
  XNOR2_X1 U433 ( .A(G143), .B(G104), .ZN(n531) );
  XOR2_X1 U434 ( .A(G140), .B(G113), .Z(n532) );
  XNOR2_X1 U435 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n458) );
  NAND2_X1 U436 ( .A1(G237), .A2(G234), .ZN(n481) );
  INV_X1 U437 ( .A(KEYINPUT114), .ZN(n638) );
  XNOR2_X1 U438 ( .A(KEYINPUT16), .B(G122), .ZN(n515) );
  XNOR2_X1 U439 ( .A(G134), .B(G107), .ZN(n541) );
  XNOR2_X1 U440 ( .A(KEYINPUT102), .B(KEYINPUT104), .ZN(n543) );
  XOR2_X1 U441 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n544) );
  INV_X1 U442 ( .A(KEYINPUT30), .ZN(n511) );
  INV_X1 U443 ( .A(KEYINPUT19), .ZN(n569) );
  AND2_X1 U444 ( .A1(n385), .A2(G953), .ZN(n570) );
  INV_X1 U445 ( .A(G898), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n435), .B(KEYINPUT42), .ZN(n801) );
  INV_X1 U447 ( .A(KEYINPUT40), .ZN(n433) );
  NOR2_X1 U448 ( .A1(n652), .A2(n745), .ZN(n730) );
  INV_X1 U449 ( .A(KEYINPUT106), .ZN(n401) );
  XNOR2_X1 U450 ( .A(n421), .B(n420), .ZN(n700) );
  INV_X1 U451 ( .A(n699), .ZN(n420) );
  INV_X1 U452 ( .A(KEYINPUT60), .ZN(n416) );
  INV_X1 U453 ( .A(KEYINPUT56), .ZN(n418) );
  AND2_X1 U454 ( .A1(n658), .A2(KEYINPUT81), .ZN(n349) );
  AND2_X1 U455 ( .A1(n665), .A2(n349), .ZN(n350) );
  XNOR2_X1 U456 ( .A(KEYINPUT77), .B(KEYINPUT23), .ZN(n351) );
  NOR2_X1 U457 ( .A1(n755), .A2(n754), .ZN(n352) );
  AND2_X1 U458 ( .A1(n528), .A2(G214), .ZN(n353) );
  XOR2_X1 U459 ( .A(n501), .B(n500), .Z(n354) );
  AND2_X1 U460 ( .A1(n760), .A2(n759), .ZN(n355) );
  AND2_X1 U461 ( .A1(n745), .A2(n560), .ZN(n356) );
  AND2_X1 U462 ( .A1(n514), .A2(n513), .ZN(n357) );
  AND2_X1 U463 ( .A1(n350), .A2(n396), .ZN(n358) );
  AND2_X1 U464 ( .A1(n378), .A2(n377), .ZN(n359) );
  XNOR2_X1 U465 ( .A(KEYINPUT59), .B(n687), .ZN(n361) );
  XOR2_X1 U466 ( .A(KEYINPUT71), .B(KEYINPUT44), .Z(n362) );
  INV_X1 U467 ( .A(n661), .ZN(n662) );
  INV_X1 U468 ( .A(KEYINPUT65), .ZN(n663) );
  INV_X1 U469 ( .A(KEYINPUT81), .ZN(n659) );
  XOR2_X1 U470 ( .A(KEYINPUT90), .B(n680), .Z(n694) );
  XNOR2_X1 U471 ( .A(n364), .B(G134), .ZN(n488) );
  XNOR2_X1 U472 ( .A(n364), .B(n363), .ZN(n533) );
  INV_X1 U473 ( .A(KEYINPUT11), .ZN(n363) );
  XNOR2_X2 U474 ( .A(KEYINPUT69), .B(G131), .ZN(n364) );
  INV_X1 U475 ( .A(n494), .ZN(n368) );
  NAND2_X1 U476 ( .A1(n494), .A2(G902), .ZN(n370) );
  NAND2_X1 U477 ( .A1(n699), .A2(n367), .ZN(n477) );
  XNOR2_X1 U478 ( .A(n372), .B(n469), .ZN(n699) );
  XNOR2_X1 U479 ( .A(n373), .B(n437), .ZN(n372) );
  XNOR2_X1 U480 ( .A(n468), .B(n351), .ZN(n373) );
  NAND2_X1 U481 ( .A1(n359), .A2(n374), .ZN(n382) );
  INV_X1 U482 ( .A(n802), .ZN(n375) );
  NOR2_X1 U483 ( .A1(n801), .A2(n379), .ZN(n376) );
  AND2_X1 U484 ( .A1(n384), .A2(n380), .ZN(n383) );
  XNOR2_X1 U485 ( .A(n646), .B(KEYINPUT47), .ZN(n380) );
  NAND2_X1 U486 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U487 ( .A1(n350), .A2(n440), .ZN(n398) );
  NAND2_X1 U488 ( .A1(n387), .A2(G224), .ZN(n519) );
  NAND2_X1 U489 ( .A1(n387), .A2(G234), .ZN(n467) );
  NAND2_X1 U490 ( .A1(n387), .A2(G227), .ZN(n490) );
  NAND2_X1 U491 ( .A1(n387), .A2(G952), .ZN(n571) );
  NAND2_X1 U492 ( .A1(n440), .A2(n387), .ZN(n784) );
  NAND2_X1 U493 ( .A1(n794), .A2(n387), .ZN(n799) );
  XNOR2_X2 U494 ( .A(G116), .B(KEYINPUT3), .ZN(n388) );
  NAND2_X1 U495 ( .A1(n358), .A2(n440), .ZN(n395) );
  NAND2_X1 U496 ( .A1(n391), .A2(n389), .ZN(n674) );
  NAND2_X1 U497 ( .A1(n390), .A2(n399), .ZN(n389) );
  NAND2_X1 U498 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U499 ( .A(n397), .ZN(n396) );
  AND2_X2 U500 ( .A1(n443), .A2(n441), .ZN(n399) );
  XOR2_X1 U501 ( .A(G146), .B(G125), .Z(n400) );
  XNOR2_X1 U502 ( .A(n507), .B(n489), .ZN(n792) );
  NAND2_X1 U503 ( .A1(n429), .A2(n426), .ZN(n648) );
  XNOR2_X1 U504 ( .A(G143), .B(G128), .ZN(n403) );
  XNOR2_X2 U505 ( .A(n619), .B(n618), .ZN(n690) );
  XNOR2_X1 U506 ( .A(G128), .B(G110), .ZN(n459) );
  XNOR2_X2 U507 ( .A(n599), .B(n598), .ZN(n610) );
  NOR2_X2 U508 ( .A1(G953), .A2(n779), .ZN(n780) );
  XNOR2_X2 U509 ( .A(n400), .B(n458), .ZN(n791) );
  BUF_X1 U510 ( .A(n684), .Z(n404) );
  BUF_X1 U511 ( .A(n597), .Z(n745) );
  XNOR2_X2 U512 ( .A(n548), .B(KEYINPUT4), .ZN(n522) );
  NAND2_X1 U513 ( .A1(n665), .A2(n658), .ZN(n442) );
  BUF_X1 U514 ( .A(n665), .Z(n793) );
  NOR2_X2 U515 ( .A1(n684), .A2(n658), .ZN(n406) );
  AND2_X1 U516 ( .A1(n525), .A2(G210), .ZN(n407) );
  XOR2_X1 U517 ( .A(G122), .B(G116), .Z(n542) );
  NAND2_X1 U518 ( .A1(n442), .A2(n659), .ZN(n441) );
  NAND2_X1 U519 ( .A1(n738), .A2(KEYINPUT109), .ZN(n408) );
  BUF_X1 U520 ( .A(n424), .Z(n409) );
  XNOR2_X1 U521 ( .A(n425), .B(n409), .ZN(n410) );
  XNOR2_X1 U522 ( .A(n425), .B(n424), .ZN(n516) );
  XNOR2_X1 U523 ( .A(n516), .B(n515), .ZN(n423) );
  XNOR2_X1 U524 ( .A(n412), .B(n411), .ZN(n771) );
  NOR2_X2 U525 ( .A1(n793), .A2(KEYINPUT2), .ZN(n412) );
  BUF_X1 U526 ( .A(n785), .Z(n413) );
  XNOR2_X1 U527 ( .A(n415), .B(n569), .ZN(n414) );
  XNOR2_X1 U528 ( .A(n648), .B(n569), .ZN(n643) );
  NOR2_X1 U529 ( .A1(n687), .A2(G902), .ZN(n540) );
  BUF_X1 U530 ( .A(n664), .Z(n770) );
  XNOR2_X2 U531 ( .A(n624), .B(KEYINPUT32), .ZN(n800) );
  NAND2_X1 U532 ( .A1(n445), .A2(n408), .ZN(n444) );
  INV_X1 U533 ( .A(n738), .ZN(n453) );
  NAND2_X1 U534 ( .A1(n594), .A2(n747), .ZN(n595) );
  BUF_X1 U535 ( .A(n741), .Z(n764) );
  XNOR2_X1 U536 ( .A(n456), .B(n615), .ZN(n455) );
  NAND2_X1 U537 ( .A1(n741), .A2(n614), .ZN(n456) );
  NAND2_X1 U538 ( .A1(n429), .A2(n426), .ZN(n415) );
  XNOR2_X1 U539 ( .A(n417), .B(n416), .ZN(G60) );
  NAND2_X1 U540 ( .A1(n689), .A2(n694), .ZN(n417) );
  XNOR2_X1 U541 ( .A(n419), .B(n418), .ZN(G51) );
  NAND2_X1 U542 ( .A1(n686), .A2(n694), .ZN(n419) );
  BUF_X1 U543 ( .A(n596), .Z(n614) );
  NAND2_X1 U544 ( .A1(n698), .A2(G217), .ZN(n421) );
  XNOR2_X1 U545 ( .A(n518), .B(KEYINPUT17), .ZN(n521) );
  XNOR2_X2 U546 ( .A(G110), .B(G107), .ZN(n424) );
  XNOR2_X2 U547 ( .A(G104), .B(G101), .ZN(n425) );
  INV_X1 U548 ( .A(n405), .ZN(n428) );
  AND2_X2 U549 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U550 ( .A1(n634), .A2(n432), .ZN(n431) );
  INV_X1 U551 ( .A(n757), .ZN(n765) );
  XNOR2_X2 U552 ( .A(n434), .B(n433), .ZN(n802) );
  NAND2_X1 U553 ( .A1(n656), .A2(n724), .ZN(n434) );
  INV_X1 U554 ( .A(n644), .ZN(n436) );
  NOR2_X1 U555 ( .A1(n655), .A2(n654), .ZN(n669) );
  NOR2_X2 U556 ( .A1(n655), .A2(n438), .ZN(n665) );
  AND2_X2 U557 ( .A1(n608), .A2(n607), .ZN(n631) );
  INV_X1 U558 ( .A(n664), .ZN(n440) );
  NAND2_X1 U559 ( .A1(n664), .A2(n659), .ZN(n443) );
  NAND2_X1 U560 ( .A1(n447), .A2(n444), .ZN(n608) );
  NAND2_X1 U561 ( .A1(n446), .A2(n453), .ZN(n445) );
  NAND2_X1 U562 ( .A1(n726), .A2(KEYINPUT109), .ZN(n446) );
  NAND2_X1 U563 ( .A1(n449), .A2(n453), .ZN(n448) );
  AND2_X2 U564 ( .A1(n709), .A2(KEYINPUT109), .ZN(n449) );
  NAND2_X1 U565 ( .A1(n452), .A2(n451), .ZN(n450) );
  INV_X1 U566 ( .A(n726), .ZN(n451) );
  NOR2_X1 U567 ( .A1(n709), .A2(KEYINPUT109), .ZN(n452) );
  XNOR2_X2 U568 ( .A(n595), .B(KEYINPUT97), .ZN(n709) );
  NAND2_X1 U569 ( .A1(n626), .A2(n690), .ZN(n454) );
  NAND2_X1 U570 ( .A1(n454), .A2(n627), .ZN(n628) );
  NAND2_X1 U571 ( .A1(n455), .A2(n617), .ZN(n619) );
  XNOR2_X1 U572 ( .A(n405), .B(KEYINPUT38), .ZN(n734) );
  XNOR2_X2 U573 ( .A(n676), .B(n675), .ZN(n701) );
  NAND2_X1 U574 ( .A1(n674), .A2(n673), .ZN(n676) );
  XNOR2_X1 U575 ( .A(n529), .B(n353), .ZN(n530) );
  XNOR2_X1 U576 ( .A(n791), .B(n530), .ZN(n536) );
  BUF_X1 U577 ( .A(n709), .Z(n711) );
  INV_X1 U578 ( .A(n457), .ZN(n518) );
  INV_X1 U579 ( .A(n791), .ZN(n462) );
  XOR2_X1 U580 ( .A(KEYINPUT24), .B(G119), .Z(n460) );
  XNOR2_X1 U581 ( .A(n460), .B(n459), .ZN(n463) );
  INV_X1 U582 ( .A(n463), .ZN(n461) );
  NAND2_X1 U583 ( .A1(n462), .A2(n461), .ZN(n465) );
  NAND2_X1 U584 ( .A1(n463), .A2(n791), .ZN(n464) );
  NAND2_X1 U585 ( .A1(n465), .A2(n464), .ZN(n469) );
  XNOR2_X1 U586 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n466) );
  XNOR2_X1 U587 ( .A(n467), .B(n466), .ZN(n547) );
  XNOR2_X2 U588 ( .A(G140), .B(G137), .ZN(n489) );
  XNOR2_X1 U589 ( .A(n489), .B(KEYINPUT94), .ZN(n468) );
  XNOR2_X1 U590 ( .A(n470), .B(n367), .ZN(n660) );
  NAND2_X1 U591 ( .A1(n660), .A2(G234), .ZN(n471) );
  XNOR2_X1 U592 ( .A(n471), .B(KEYINPUT20), .ZN(n478) );
  NAND2_X1 U593 ( .A1(n478), .A2(G217), .ZN(n475) );
  XNOR2_X1 U594 ( .A(KEYINPUT25), .B(KEYINPUT76), .ZN(n473) );
  INV_X1 U595 ( .A(KEYINPUT75), .ZN(n472) );
  XNOR2_X1 U596 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U597 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U598 ( .A1(n478), .A2(G221), .ZN(n479) );
  XNOR2_X1 U599 ( .A(n479), .B(KEYINPUT21), .ZN(n750) );
  INV_X1 U600 ( .A(KEYINPUT14), .ZN(n480) );
  XNOR2_X1 U601 ( .A(n481), .B(n480), .ZN(n762) );
  NAND2_X1 U602 ( .A1(G953), .A2(G902), .ZN(n482) );
  NOR2_X1 U603 ( .A1(n762), .A2(n482), .ZN(n483) );
  XNOR2_X1 U604 ( .A(n483), .B(KEYINPUT113), .ZN(n484) );
  NOR2_X1 U605 ( .A1(G900), .A2(n484), .ZN(n486) );
  NOR2_X1 U606 ( .A1(n762), .A2(n571), .ZN(n485) );
  NOR2_X1 U607 ( .A1(n486), .A2(n485), .ZN(n487) );
  NOR2_X1 U608 ( .A1(n750), .A2(n487), .ZN(n561) );
  NAND2_X1 U609 ( .A1(n560), .A2(n561), .ZN(n495) );
  XNOR2_X2 U610 ( .A(G143), .B(G128), .ZN(n548) );
  XNOR2_X2 U611 ( .A(n488), .B(n522), .ZN(n507) );
  XNOR2_X1 U612 ( .A(n490), .B(G146), .ZN(n491) );
  XNOR2_X1 U613 ( .A(n410), .B(n491), .ZN(n492) );
  INV_X1 U614 ( .A(KEYINPUT70), .ZN(n493) );
  XNOR2_X1 U615 ( .A(n493), .B(G469), .ZN(n494) );
  NOR2_X1 U616 ( .A1(n495), .A2(n641), .ZN(n496) );
  XNOR2_X1 U617 ( .A(n496), .B(KEYINPUT74), .ZN(n514) );
  NAND2_X1 U618 ( .A1(n367), .A2(n497), .ZN(n525) );
  NAND2_X1 U619 ( .A1(n525), .A2(G214), .ZN(n733) );
  XNOR2_X1 U620 ( .A(n498), .B(G113), .ZN(n499) );
  INV_X1 U621 ( .A(n517), .ZN(n506) );
  NAND2_X1 U622 ( .A1(n528), .A2(G210), .ZN(n502) );
  XNOR2_X1 U623 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U624 ( .A(n354), .B(n504), .ZN(n505) );
  XNOR2_X1 U625 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U626 ( .A(n508), .B(n507), .ZN(n691) );
  NAND2_X1 U627 ( .A1(n691), .A2(n367), .ZN(n510) );
  INV_X1 U628 ( .A(G472), .ZN(n509) );
  INV_X1 U629 ( .A(n558), .ZN(n600) );
  NAND2_X1 U630 ( .A1(n733), .A2(n600), .ZN(n512) );
  XNOR2_X1 U631 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U632 ( .A(n519), .B(KEYINPUT18), .ZN(n520) );
  XNOR2_X1 U633 ( .A(n521), .B(n520), .ZN(n523) );
  XNOR2_X1 U634 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U635 ( .A(n785), .B(n524), .ZN(n684) );
  INV_X1 U636 ( .A(n660), .ZN(n658) );
  INV_X1 U637 ( .A(n405), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n357), .A2(n566), .ZN(n557) );
  XOR2_X1 U639 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n527) );
  XNOR2_X1 U640 ( .A(n527), .B(n526), .ZN(n529) );
  XNOR2_X1 U641 ( .A(n532), .B(n531), .ZN(n534) );
  XNOR2_X1 U642 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U643 ( .A(n536), .B(n535), .ZN(n687) );
  XOR2_X1 U644 ( .A(KEYINPUT101), .B(KEYINPUT13), .Z(n538) );
  XNOR2_X1 U645 ( .A(KEYINPUT100), .B(G475), .ZN(n537) );
  XNOR2_X1 U646 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U647 ( .A(n540), .B(n539), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n542), .B(n541), .ZN(n546) );
  XNOR2_X1 U649 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U650 ( .A(n546), .B(n545), .Z(n552) );
  NAND2_X1 U651 ( .A1(G217), .A2(n547), .ZN(n550) );
  XNOR2_X1 U652 ( .A(n403), .B(KEYINPUT9), .ZN(n549) );
  XNOR2_X1 U653 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U654 ( .A(n552), .B(n551), .ZN(n677) );
  NOR2_X1 U655 ( .A1(G902), .A2(n677), .ZN(n554) );
  XNOR2_X1 U656 ( .A(G478), .B(KEYINPUT105), .ZN(n553) );
  XNOR2_X1 U657 ( .A(n554), .B(n553), .ZN(n602) );
  AND2_X1 U658 ( .A1(n579), .A2(n602), .ZN(n556) );
  INV_X1 U659 ( .A(KEYINPUT112), .ZN(n555) );
  XNOR2_X1 U660 ( .A(n556), .B(n555), .ZN(n616) );
  NOR2_X1 U661 ( .A1(n557), .A2(n616), .ZN(n653) );
  XOR2_X1 U662 ( .A(G143), .B(n653), .Z(G45) );
  NOR2_X1 U663 ( .A1(n602), .A2(n603), .ZN(n724) );
  INV_X1 U664 ( .A(KEYINPUT6), .ZN(n559) );
  INV_X1 U665 ( .A(n560), .ZN(n749) );
  NAND2_X1 U666 ( .A1(n561), .A2(n749), .ZN(n637) );
  NOR2_X1 U667 ( .A1(n620), .A2(n637), .ZN(n562) );
  NAND2_X1 U668 ( .A1(n724), .A2(n562), .ZN(n647) );
  INV_X1 U669 ( .A(n733), .ZN(n568) );
  NOR2_X1 U670 ( .A1(n647), .A2(n568), .ZN(n564) );
  XNOR2_X1 U671 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n563) );
  NAND2_X1 U672 ( .A1(n564), .A2(n745), .ZN(n565) );
  XOR2_X1 U673 ( .A(KEYINPUT43), .B(n565), .Z(n567) );
  NOR2_X1 U674 ( .A1(n567), .A2(n566), .ZN(n654) );
  XOR2_X1 U675 ( .A(G140), .B(n654), .Z(G42) );
  XOR2_X1 U676 ( .A(KEYINPUT93), .B(n570), .Z(n786) );
  NAND2_X1 U677 ( .A1(n786), .A2(G902), .ZN(n572) );
  NAND2_X1 U678 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U679 ( .A(n762), .ZN(n573) );
  AND2_X1 U680 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U681 ( .A1(n643), .A2(n575), .ZN(n578) );
  XNOR2_X1 U682 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n576) );
  XNOR2_X1 U683 ( .A(n576), .B(KEYINPUT67), .ZN(n577) );
  XNOR2_X2 U684 ( .A(n578), .B(n577), .ZN(n596) );
  INV_X1 U685 ( .A(n602), .ZN(n580) );
  NAND2_X1 U686 ( .A1(n603), .A2(n580), .ZN(n736) );
  NOR2_X1 U687 ( .A1(n736), .A2(n750), .ZN(n581) );
  NAND2_X1 U688 ( .A1(n596), .A2(n581), .ZN(n583) );
  INV_X1 U689 ( .A(KEYINPUT22), .ZN(n582) );
  XNOR2_X2 U690 ( .A(n583), .B(n582), .ZN(n622) );
  AND2_X1 U691 ( .A1(n591), .A2(n747), .ZN(n584) );
  AND2_X1 U692 ( .A1(n745), .A2(n584), .ZN(n585) );
  NAND2_X1 U693 ( .A1(n622), .A2(n585), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n625), .B(G110), .ZN(G12) );
  NAND2_X1 U695 ( .A1(n622), .A2(n620), .ZN(n586) );
  XNOR2_X1 U696 ( .A(n586), .B(KEYINPUT84), .ZN(n587) );
  INV_X1 U697 ( .A(n587), .ZN(n588) );
  NAND2_X1 U698 ( .A1(n588), .A2(n356), .ZN(n589) );
  XNOR2_X1 U699 ( .A(G101), .B(KEYINPUT116), .ZN(n590) );
  XNOR2_X1 U700 ( .A(n607), .B(n590), .ZN(G3) );
  OR2_X1 U701 ( .A1(n591), .A2(n750), .ZN(n744) );
  NOR2_X1 U702 ( .A1(n641), .A2(n744), .ZN(n592) );
  NAND2_X1 U703 ( .A1(n596), .A2(n592), .ZN(n593) );
  XNOR2_X1 U704 ( .A(n593), .B(KEYINPUT95), .ZN(n594) );
  INV_X1 U705 ( .A(KEYINPUT72), .ZN(n598) );
  AND2_X1 U706 ( .A1(n610), .A2(n600), .ZN(n754) );
  NAND2_X1 U707 ( .A1(n614), .A2(n754), .ZN(n601) );
  XNOR2_X1 U708 ( .A(n601), .B(KEYINPUT31), .ZN(n726) );
  NAND2_X1 U709 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U710 ( .A(KEYINPUT107), .B(n727), .Z(n657) );
  INV_X1 U711 ( .A(KEYINPUT108), .ZN(n605) );
  XNOR2_X1 U712 ( .A(n606), .B(n605), .ZN(n645) );
  BUF_X1 U713 ( .A(n645), .Z(n738) );
  INV_X1 U714 ( .A(n620), .ZN(n609) );
  NAND2_X1 U715 ( .A1(n610), .A2(n609), .ZN(n613) );
  XNOR2_X1 U716 ( .A(KEYINPUT111), .B(KEYINPUT33), .ZN(n611) );
  XNOR2_X1 U717 ( .A(n611), .B(KEYINPUT89), .ZN(n612) );
  INV_X1 U718 ( .A(KEYINPUT34), .ZN(n615) );
  INV_X1 U719 ( .A(n616), .ZN(n617) );
  XNOR2_X1 U720 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n618) );
  NOR2_X1 U721 ( .A1(n745), .A2(n560), .ZN(n621) );
  AND2_X1 U722 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U723 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U724 ( .A1(n402), .A2(n362), .ZN(n629) );
  NOR2_X1 U725 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n627) );
  NAND2_X1 U726 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U727 ( .A1(n631), .A2(n630), .ZN(n633) );
  INV_X1 U728 ( .A(KEYINPUT45), .ZN(n632) );
  XNOR2_X2 U729 ( .A(n633), .B(n632), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n357), .A2(n734), .ZN(n635) );
  NAND2_X1 U731 ( .A1(n734), .A2(n733), .ZN(n737) );
  NOR2_X1 U732 ( .A1(n737), .A2(n736), .ZN(n636) );
  XNOR2_X1 U733 ( .A(n636), .B(KEYINPUT41), .ZN(n757) );
  NOR2_X1 U734 ( .A1(n747), .A2(n637), .ZN(n640) );
  XNOR2_X1 U735 ( .A(n640), .B(n639), .ZN(n642) );
  NOR2_X1 U736 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U737 ( .A1(n644), .A2(n414), .ZN(n722) );
  NOR2_X1 U738 ( .A1(n645), .A2(n722), .ZN(n646) );
  XNOR2_X1 U739 ( .A(n647), .B(KEYINPUT115), .ZN(n649) );
  NAND2_X1 U740 ( .A1(n649), .A2(n415), .ZN(n651) );
  XOR2_X1 U741 ( .A(KEYINPUT85), .B(KEYINPUT36), .Z(n650) );
  XNOR2_X1 U742 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U743 ( .A1(n656), .A2(n657), .ZN(n732) );
  INV_X1 U744 ( .A(KEYINPUT2), .ZN(n769) );
  NOR2_X1 U745 ( .A1(n660), .A2(n769), .ZN(n661) );
  AND2_X1 U746 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n793), .A2(n666), .ZN(n671) );
  AND2_X1 U748 ( .A1(n732), .A2(KEYINPUT2), .ZN(n667) );
  NOR2_X1 U749 ( .A1(n667), .A2(KEYINPUT78), .ZN(n668) );
  NAND2_X1 U750 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n672) );
  AND2_X1 U752 ( .A1(n440), .A2(n672), .ZN(n773) );
  INV_X1 U753 ( .A(n773), .ZN(n673) );
  INV_X1 U754 ( .A(KEYINPUT64), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n701), .A2(G478), .ZN(n679) );
  INV_X1 U756 ( .A(n677), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U758 ( .A1(n681), .A2(n694), .ZN(n682) );
  XNOR2_X1 U759 ( .A(n682), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n701), .A2(G210), .ZN(n685) );
  XOR2_X1 U761 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n683) );
  XNOR2_X1 U762 ( .A(n685), .B(n360), .ZN(n686) );
  INV_X1 U763 ( .A(n694), .ZN(n707) );
  NAND2_X1 U764 ( .A1(n701), .A2(G475), .ZN(n688) );
  XNOR2_X1 U765 ( .A(n688), .B(n361), .ZN(n689) );
  XNOR2_X1 U766 ( .A(n690), .B(G122), .ZN(G24) );
  NAND2_X1 U767 ( .A1(n701), .A2(G472), .ZN(n693) );
  XNOR2_X1 U768 ( .A(n691), .B(KEYINPUT62), .ZN(n692) );
  XNOR2_X1 U769 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U770 ( .A1(n695), .A2(n694), .ZN(n697) );
  XOR2_X1 U771 ( .A(KEYINPUT87), .B(KEYINPUT63), .Z(n696) );
  XNOR2_X1 U772 ( .A(n697), .B(n696), .ZN(G57) );
  BUF_X1 U773 ( .A(n701), .Z(n698) );
  NOR2_X1 U774 ( .A1(n700), .A2(n707), .ZN(G66) );
  NAND2_X1 U775 ( .A1(n698), .A2(G469), .ZN(n706) );
  XOR2_X1 U776 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n702) );
  XNOR2_X1 U777 ( .A(n702), .B(KEYINPUT58), .ZN(n703) );
  XNOR2_X1 U778 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U779 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U780 ( .A1(n708), .A2(n707), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n711), .A2(n724), .ZN(n710) );
  XNOR2_X1 U782 ( .A(n710), .B(G104), .ZN(G6) );
  XOR2_X1 U783 ( .A(KEYINPUT118), .B(KEYINPUT27), .Z(n713) );
  NAND2_X1 U784 ( .A1(n711), .A2(n727), .ZN(n712) );
  XNOR2_X1 U785 ( .A(n713), .B(n712), .ZN(n714) );
  XOR2_X1 U786 ( .A(n714), .B(KEYINPUT26), .Z(n716) );
  XNOR2_X1 U787 ( .A(G107), .B(KEYINPUT117), .ZN(n715) );
  XNOR2_X1 U788 ( .A(n716), .B(n715), .ZN(G9) );
  INV_X1 U789 ( .A(n727), .ZN(n717) );
  NOR2_X1 U790 ( .A1(n722), .A2(n717), .ZN(n719) );
  XNOR2_X1 U791 ( .A(KEYINPUT119), .B(KEYINPUT29), .ZN(n718) );
  XNOR2_X1 U792 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U793 ( .A(G128), .B(n720), .Z(G30) );
  INV_X1 U794 ( .A(n724), .ZN(n721) );
  NOR2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U796 ( .A(G146), .B(n723), .Z(G48) );
  NAND2_X1 U797 ( .A1(n726), .A2(n724), .ZN(n725) );
  XNOR2_X1 U798 ( .A(n725), .B(G113), .ZN(G15) );
  NAND2_X1 U799 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U800 ( .A(n728), .B(KEYINPUT120), .ZN(n729) );
  XNOR2_X1 U801 ( .A(G116), .B(n729), .ZN(G18) );
  XNOR2_X1 U802 ( .A(n730), .B(G125), .ZN(n731) );
  XNOR2_X1 U803 ( .A(n731), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U804 ( .A(G134), .B(n732), .ZN(G36) );
  NOR2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n740) );
  NOR2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U808 ( .A1(n740), .A2(n739), .ZN(n743) );
  INV_X1 U809 ( .A(n764), .ZN(n742) );
  OR2_X1 U810 ( .A1(n743), .A2(n742), .ZN(n760) );
  XNOR2_X1 U811 ( .A(KEYINPUT121), .B(KEYINPUT51), .ZN(n756) );
  NAND2_X1 U812 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U813 ( .A(n746), .B(KEYINPUT50), .ZN(n748) );
  NAND2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n753) );
  NAND2_X1 U815 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U816 ( .A(KEYINPUT49), .B(n751), .ZN(n752) );
  NOR2_X1 U817 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U818 ( .A(n756), .B(n352), .ZN(n758) );
  OR2_X1 U819 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U820 ( .A(n355), .B(KEYINPUT52), .ZN(n761) );
  NOR2_X1 U821 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U822 ( .A1(n763), .A2(G952), .ZN(n767) );
  NAND2_X1 U823 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U824 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U825 ( .A(KEYINPUT122), .B(n768), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U827 ( .A1(n772), .A2(n771), .ZN(n774) );
  NOR2_X1 U828 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U829 ( .A(n775), .B(KEYINPUT82), .ZN(n776) );
  NOR2_X1 U830 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U831 ( .A(n778), .B(KEYINPUT123), .ZN(n779) );
  XNOR2_X1 U832 ( .A(KEYINPUT53), .B(n780), .ZN(G75) );
  NAND2_X1 U833 ( .A1(G953), .A2(G224), .ZN(n781) );
  XNOR2_X1 U834 ( .A(KEYINPUT61), .B(n781), .ZN(n782) );
  NAND2_X1 U835 ( .A1(n782), .A2(G898), .ZN(n783) );
  NAND2_X1 U836 ( .A1(n784), .A2(n783), .ZN(n789) );
  XOR2_X1 U837 ( .A(KEYINPUT126), .B(n413), .Z(n787) );
  NOR2_X1 U838 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U839 ( .A(n789), .B(n788), .ZN(n790) );
  XOR2_X1 U840 ( .A(KEYINPUT127), .B(n790), .Z(G69) );
  XNOR2_X1 U841 ( .A(n792), .B(n791), .ZN(n795) );
  XNOR2_X1 U842 ( .A(n793), .B(n795), .ZN(n794) );
  XOR2_X1 U843 ( .A(G227), .B(n795), .Z(n796) );
  NAND2_X1 U844 ( .A1(n796), .A2(G900), .ZN(n797) );
  NAND2_X1 U845 ( .A1(n797), .A2(G953), .ZN(n798) );
  NAND2_X1 U846 ( .A1(n799), .A2(n798), .ZN(G72) );
  XNOR2_X1 U847 ( .A(G119), .B(n800), .ZN(G21) );
  XOR2_X1 U848 ( .A(n801), .B(G137), .Z(G39) );
  XOR2_X1 U849 ( .A(n802), .B(G131), .Z(G33) );
endmodule

