//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT67), .B1(new_n189), .B2(G116), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(G119), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n196), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n195), .B1(new_n190), .B2(new_n193), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n201), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n197), .B1(new_n209), .B2(new_n195), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n203), .A2(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT76), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT76), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT77), .B(new_n212), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(KEYINPUT76), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(G104), .ZN(new_n219));
  AOI21_X1  g033(.A(G107), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n212), .B2(G104), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n217), .B(G101), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G107), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(G104), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G107), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n218), .A3(new_n219), .ZN(new_n228));
  INV_X1    g042(.A(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n223), .A2(KEYINPUT78), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT78), .B1(new_n223), .B2(new_n230), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n211), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n205), .B1(new_n204), .B2(new_n201), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n234), .A2(new_n235), .B1(new_n204), .B2(new_n201), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n229), .B1(new_n226), .B2(new_n228), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n226), .A2(new_n228), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n230), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(KEYINPUT82), .A3(new_n239), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT82), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n230), .A2(KEYINPUT4), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(new_n245), .B2(new_n237), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n204), .A2(new_n201), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n203), .B2(new_n206), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n244), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n233), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G110), .B(G122), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n233), .A2(new_n243), .A3(new_n249), .A4(new_n251), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(KEYINPUT6), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n256), .A3(new_n252), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G146), .ZN(new_n260));
  INV_X1    g074(.A(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT65), .A3(G143), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(G146), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n260), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n261), .A2(G143), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n267), .A2(new_n269), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n259), .A2(G146), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n261), .A2(G143), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n266), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G125), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  OR2_X1    g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(new_n280), .C1(new_n272), .C2(new_n273), .ZN(new_n281));
  INV_X1    g095(.A(new_n279), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n260), .A2(new_n262), .A3(new_n282), .A4(new_n265), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G125), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G953), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G224), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n286), .B(new_n288), .Z(new_n289));
  NAND3_X1  g103(.A1(new_n255), .A2(new_n257), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT84), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT84), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n255), .A2(new_n292), .A3(new_n257), .A4(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT87), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n210), .A2(new_n297), .B1(new_n204), .B2(KEYINPUT5), .ZN(new_n298));
  OAI21_X1  g112(.A(G113), .B1(new_n207), .B2(new_n196), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT86), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n298), .A2(new_n300), .B1(new_n203), .B2(new_n206), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n231), .B2(new_n232), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n208), .A2(new_n210), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n234), .B2(new_n235), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n223), .A2(new_n230), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n251), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n296), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  AOI211_X1 g125(.A(KEYINPUT87), .B(new_n309), .C1(new_n302), .C2(new_n306), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT7), .B1(new_n288), .B2(KEYINPUT89), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(KEYINPUT89), .B2(new_n288), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n278), .A2(new_n285), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT90), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n278), .A2(new_n318), .A3(new_n285), .A4(new_n315), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT88), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n278), .A2(new_n285), .B1(KEYINPUT7), .B2(new_n288), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n317), .A2(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n321), .A2(new_n320), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n254), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n295), .B1(new_n313), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n294), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G210), .B1(G237), .B2(G902), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n294), .A2(new_n326), .A3(new_n328), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n188), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G217), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(G234), .B2(new_n295), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT66), .B(G128), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n189), .A2(G128), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT71), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n341), .A3(new_n338), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT24), .B(G110), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT72), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n340), .A2(new_n347), .A3(new_n342), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G125), .B(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT16), .ZN(new_n351));
  INV_X1    g165(.A(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G125), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n353), .A2(KEYINPUT16), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n261), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(G146), .A3(new_n354), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n189), .B2(G128), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n338), .B(new_n360), .C1(new_n337), .C2(new_n359), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G110), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n349), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n351), .A2(KEYINPUT73), .A3(new_n354), .A4(G146), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n350), .A2(new_n261), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n361), .A2(G110), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n337), .A2(new_n341), .A3(new_n338), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n341), .B1(new_n337), .B2(new_n338), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n343), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT22), .B(G137), .ZN(new_n377));
  INV_X1    g191(.A(G221), .ZN(new_n378));
  INV_X1    g192(.A(G234), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n378), .A2(new_n379), .A3(G953), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n377), .B(new_n380), .Z(new_n381));
  NAND3_X1  g195(.A1(new_n365), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n381), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n363), .B1(new_n346), .B2(new_n348), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n375), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n386), .A2(new_n387), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n335), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n390), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n382), .A2(new_n385), .A3(new_n392), .A4(new_n388), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n382), .A2(new_n385), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n334), .A2(G902), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n281), .A2(new_n283), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT11), .ZN(new_n400));
  INV_X1    g214(.A(G134), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(G137), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(G137), .ZN(new_n403));
  INV_X1    g217(.A(G137), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT11), .A3(G134), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G131), .ZN(new_n407));
  INV_X1    g221(.A(G131), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n402), .A2(new_n405), .A3(new_n408), .A4(new_n403), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n399), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n401), .A2(G137), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n404), .A2(G134), .ZN(new_n413));
  OAI21_X1  g227(.A(G131), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n267), .A2(new_n269), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n415), .A2(new_n416), .B1(new_n270), .B2(new_n265), .ZN(new_n417));
  AND4_X1   g231(.A1(new_n260), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n409), .B(new_n414), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n411), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT64), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT30), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n423));
  AOI211_X1 g237(.A(KEYINPUT64), .B(new_n423), .C1(new_n411), .C2(new_n419), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n236), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G237), .A2(G953), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G210), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT27), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(G101), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  AND4_X1   g244(.A1(KEYINPUT69), .A2(new_n248), .A3(new_n411), .A4(new_n419), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n409), .A2(new_n414), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n410), .A2(new_n399), .B1(new_n432), .B2(new_n275), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT69), .B1(new_n433), .B2(new_n248), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n425), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT31), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT31), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n425), .A2(new_n435), .A3(new_n438), .A4(new_n430), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n420), .A2(new_n236), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT28), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT69), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n420), .B2(new_n236), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT70), .B1(new_n433), .B2(new_n248), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT70), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n420), .A2(new_n445), .A3(new_n236), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n433), .A2(KEYINPUT69), .A3(new_n248), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n441), .B1(new_n448), .B2(KEYINPUT28), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n437), .B(new_n439), .C1(new_n430), .C2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G472), .A2(G902), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(KEYINPUT32), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n420), .A2(new_n236), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n443), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n441), .B1(new_n454), .B2(KEYINPUT28), .ZN(new_n455));
  INV_X1    g269(.A(new_n430), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n423), .B1(new_n433), .B2(KEYINPUT64), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT30), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n248), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n443), .A2(new_n447), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n457), .B1(new_n464), .B2(new_n430), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n456), .B(new_n441), .C1(new_n448), .C2(KEYINPUT28), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G472), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n452), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n450), .A2(new_n451), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT32), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n398), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT9), .B(G234), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n378), .B1(new_n475), .B2(new_n295), .ZN(new_n476));
  INV_X1    g290(.A(G469), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n295), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT10), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n276), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n231), .B2(new_n232), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n260), .A2(new_n265), .A3(new_n262), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT1), .ZN(new_n483));
  OAI21_X1  g297(.A(G128), .B1(new_n272), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n266), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n223), .A2(new_n486), .A3(new_n230), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n284), .B1(new_n238), .B2(new_n237), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n487), .A2(new_n479), .B1(new_n488), .B2(new_n242), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n410), .B(KEYINPUT79), .Z(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G140), .ZN(new_n492));
  INV_X1    g306(.A(G227), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(G953), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n410), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n481), .B2(new_n489), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n410), .A2(KEYINPUT80), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n231), .A2(new_n232), .A3(new_n275), .ZN(new_n502));
  INV_X1    g316(.A(new_n487), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT12), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n506), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n491), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n495), .B(KEYINPUT75), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n500), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n478), .B1(new_n511), .B2(G469), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n481), .A2(new_n489), .A3(new_n490), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n495), .B1(new_n513), .B2(new_n499), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT81), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n505), .A2(new_n496), .A3(new_n491), .A4(new_n507), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT81), .B(new_n495), .C1(new_n513), .C2(new_n499), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n477), .A3(new_n295), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n476), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n474), .A2(new_n333), .A3(G953), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n336), .A2(G143), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n259), .A2(G128), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(G134), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT93), .B(G122), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G116), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n192), .A2(G122), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G107), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n212), .A3(new_n529), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n526), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n523), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n524), .B(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G134), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n533), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n529), .A2(KEYINPUT14), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT95), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n544));
  INV_X1    g358(.A(new_n529), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n528), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G107), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n401), .B1(new_n523), .B2(new_n524), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n547), .B(new_n532), .C1(new_n526), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n522), .B1(new_n541), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n541), .A2(new_n549), .A3(new_n522), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n295), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n554), .A2(new_n559), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n426), .A2(G143), .A3(G214), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(G143), .B1(new_n426), .B2(G214), .ZN(new_n566));
  OAI21_X1  g380(.A(G131), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n568));
  INV_X1    g382(.A(G237), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n287), .A3(G214), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n259), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n408), .A3(new_n564), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT17), .B(G131), .C1(new_n565), .C2(new_n566), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n356), .A3(new_n574), .A4(new_n357), .ZN(new_n575));
  XNOR2_X1  g389(.A(G113), .B(G122), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(new_n215), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n350), .A2(new_n261), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(KEYINPUT91), .B2(new_n369), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n277), .A2(G140), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n353), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n581), .A2(KEYINPUT91), .A3(G146), .ZN(new_n582));
  AND4_X1   g396(.A1(KEYINPUT18), .A2(new_n571), .A3(G131), .A4(new_n564), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n571), .A2(new_n564), .B1(KEYINPUT18), .B2(G131), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n579), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n577), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n577), .B1(new_n575), .B2(new_n585), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n295), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G475), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT20), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n567), .A2(new_n572), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n350), .A2(KEYINPUT19), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n350), .A2(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n261), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n367), .A2(new_n592), .A3(new_n595), .A4(new_n368), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n585), .ZN(new_n597));
  INV_X1    g411(.A(new_n577), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n586), .ZN(new_n600));
  NOR2_X1   g414(.A1(G475), .A2(G902), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n591), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n601), .ZN(new_n603));
  AOI211_X1 g417(.A(KEYINPUT20), .B(new_n603), .C1(new_n599), .C2(new_n586), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n590), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT92), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n590), .B(new_n607), .C1(new_n602), .C2(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n287), .A2(G952), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n379), .B2(new_n569), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI211_X1 g427(.A(new_n295), .B(new_n287), .C1(G234), .C2(G237), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT21), .B(G898), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n563), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n332), .A2(new_n473), .A3(new_n521), .A4(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT97), .B(G101), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G3));
  NAND2_X1  g434(.A1(new_n512), .A2(new_n520), .ZN(new_n621));
  INV_X1    g435(.A(new_n476), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n391), .A2(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n438), .B1(new_n464), .B2(new_n430), .ZN(new_n625));
  INV_X1    g439(.A(new_n439), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n449), .A2(new_n430), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(G902), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G472), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n470), .B(new_n624), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT98), .B1(new_n623), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n450), .B2(new_n295), .ZN(new_n634));
  INV_X1    g448(.A(new_n451), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n627), .B2(new_n629), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n521), .A2(new_n637), .A3(new_n638), .A4(new_n624), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n330), .A2(new_n331), .ZN(new_n641));
  INV_X1    g455(.A(new_n616), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT99), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n643), .A2(KEYINPUT99), .ZN(new_n645));
  INV_X1    g459(.A(new_n552), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n550), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n551), .A2(KEYINPUT99), .A3(new_n643), .A4(new_n552), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n555), .A2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n554), .A2(new_n555), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n609), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n641), .A2(new_n187), .A3(new_n642), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n640), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  AOI21_X1  g473(.A(new_n328), .B1(new_n294), .B2(new_n326), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n329), .B(new_n325), .C1(new_n291), .C2(new_n293), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n187), .B(new_n642), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n562), .A2(new_n605), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n639), .A3(new_n633), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  OR3_X1    g482(.A1(new_n384), .A2(KEYINPUT100), .A3(new_n375), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT100), .B1(new_n384), .B2(new_n375), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(KEYINPUT36), .B2(new_n383), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n383), .A2(KEYINPUT36), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n396), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n394), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(new_n636), .A3(new_n634), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n332), .A2(new_n521), .A3(new_n678), .A4(new_n617), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  AOI21_X1  g495(.A(new_n677), .B1(new_n469), .B2(new_n472), .ZN(new_n682));
  INV_X1    g496(.A(new_n614), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n612), .B1(new_n683), .B2(G900), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT101), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n605), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n562), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n332), .A2(new_n521), .A3(new_n682), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XNOR2_X1  g503(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n641), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n685), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n521), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n521), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n464), .A2(new_n456), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n295), .B1(new_n454), .B2(new_n430), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n472), .A2(new_n452), .A3(new_n699), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n676), .A2(new_n562), .A3(new_n188), .A4(new_n609), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n694), .A2(new_n696), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n259), .ZN(G45));
  NOR3_X1   g518(.A1(new_n654), .A2(new_n609), .A3(new_n685), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n332), .A2(new_n521), .A3(new_n682), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  NAND2_X1  g521(.A1(new_n519), .A2(new_n295), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n622), .A3(new_n520), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n473), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n656), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n662), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n452), .A2(new_n468), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT32), .B1(new_n450), .B2(new_n451), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n624), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n710), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n715), .A3(new_n719), .A4(new_n655), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  NAND3_X1  g537(.A1(new_n714), .A2(new_n663), .A3(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NAND4_X1  g539(.A1(new_n332), .A2(new_n617), .A3(new_n682), .A4(new_n711), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  AOI211_X1 g541(.A(KEYINPUT106), .B(new_n631), .C1(new_n450), .C2(new_n295), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n437), .A2(new_n439), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n295), .B1(new_n730), .B2(new_n628), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n729), .B1(new_n731), .B2(G472), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n454), .A2(KEYINPUT28), .ZN(new_n733));
  INV_X1    g547(.A(new_n441), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n735), .A2(new_n456), .B1(new_n436), .B2(KEYINPUT31), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n626), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n462), .A2(new_n463), .A3(new_n456), .ZN(new_n739));
  OAI22_X1  g553(.A1(new_n739), .A2(new_n438), .B1(new_n455), .B2(new_n430), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT104), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n635), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n728), .A2(new_n732), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n624), .B(KEYINPUT107), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n709), .A2(new_n622), .A3(new_n520), .A4(new_n642), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n439), .B1(new_n740), .B2(KEYINPUT104), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n735), .A2(new_n456), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n737), .B1(new_n748), .B2(new_n437), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n743), .B(new_n451), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n562), .A2(new_n609), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n641), .A2(new_n187), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  OAI21_X1  g571(.A(KEYINPUT106), .B1(new_n630), .B2(new_n631), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n634), .A2(new_n729), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n451), .B1(new_n747), .B2(new_n749), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n758), .A2(new_n759), .B1(KEYINPUT105), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n676), .A3(new_n705), .A4(new_n750), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n332), .A2(new_n711), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G125), .ZN(G27));
  NOR3_X1   g579(.A1(new_n660), .A2(new_n661), .A3(new_n188), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n623), .A2(KEYINPUT108), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n521), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n473), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n705), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n330), .A2(new_n187), .A3(new_n331), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n521), .A2(new_n768), .ZN(new_n775));
  AOI211_X1 g589(.A(KEYINPUT108), .B(new_n476), .C1(new_n512), .C2(new_n520), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n398), .A2(KEYINPUT107), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n624), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n452), .B(new_n468), .C1(new_n717), .C2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n636), .A2(KEYINPUT109), .A3(KEYINPUT32), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n781), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n472), .A2(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n717), .A2(new_n783), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n469), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n782), .B1(new_n790), .B2(new_n781), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n777), .B(new_n705), .C1(new_n787), .C2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n773), .B1(new_n792), .B2(KEYINPUT42), .ZN(new_n793));
  XOR2_X1   g607(.A(KEYINPUT111), .B(G131), .Z(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(G33));
  INV_X1    g609(.A(new_n687), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n770), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n401), .ZN(G36));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT43), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n653), .B2(new_n609), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n653), .A2(new_n609), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(KEYINPUT43), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n801), .B1(new_n804), .B2(new_n800), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n637), .B2(new_n677), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n676), .B(KEYINPUT115), .C1(new_n634), .C2(new_n636), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n766), .B1(new_n809), .B2(KEYINPUT44), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(KEYINPUT44), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n809), .A2(KEYINPUT116), .A3(KEYINPUT44), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n692), .A2(new_n622), .ZN(new_n816));
  OAI21_X1  g630(.A(G469), .B1(new_n511), .B2(KEYINPUT45), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n511), .A2(KEYINPUT45), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(KEYINPUT112), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n821));
  INV_X1    g635(.A(new_n819), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n817), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n478), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT46), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n520), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n478), .B1(new_n820), .B2(new_n823), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(KEYINPUT46), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n828), .B1(new_n831), .B2(KEYINPUT113), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(KEYINPUT113), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n816), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n815), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G137), .ZN(G39));
  INV_X1    g651(.A(new_n834), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n622), .B1(new_n838), .B2(new_n832), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT47), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT47), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n622), .C1(new_n838), .C2(new_n832), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n705), .A2(new_n472), .A3(new_n469), .A4(new_n398), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n774), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(G140), .ZN(G42));
  AND2_X1   g660(.A1(new_n709), .A2(new_n520), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT49), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n622), .A2(new_n187), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n745), .A2(new_n700), .A3(new_n802), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n691), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n623), .A2(new_n563), .A3(new_n686), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n682), .A3(new_n766), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n770), .B2(new_n796), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n762), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n787), .A2(new_n791), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n766), .A2(new_n767), .A3(new_n705), .A4(new_n769), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT42), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n773), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n857), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n653), .A2(new_n609), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n609), .B2(new_n562), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n633), .A2(new_n639), .A3(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n714), .A2(new_n865), .B1(new_n752), .B2(new_n755), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n618), .A2(new_n726), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n617), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n187), .B(new_n521), .C1(new_n660), .C2(new_n661), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n871), .A2(new_n678), .B1(new_n665), .B2(new_n719), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n866), .A2(new_n721), .A3(new_n868), .A4(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n862), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n688), .B(new_n706), .C1(new_n762), .C2(new_n763), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n676), .A2(new_n685), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n700), .A2(new_n521), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n754), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n879), .ZN(new_n881));
  INV_X1    g695(.A(new_n870), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n682), .C1(new_n687), .C2(new_n705), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n764), .A2(new_n881), .A3(KEYINPUT52), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(KEYINPUT117), .B(new_n875), .C1(new_n876), .C2(new_n879), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n633), .A2(new_n639), .A3(new_n864), .ZN(new_n891));
  INV_X1    g705(.A(new_n746), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n761), .A2(new_n781), .A3(new_n892), .A4(new_n750), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n891), .A2(new_n662), .B1(new_n893), .B2(new_n754), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n724), .A2(new_n679), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n867), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n793), .A3(new_n721), .A4(new_n857), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n880), .A2(new_n884), .ZN(new_n898));
  OR3_X1    g712(.A1(new_n897), .A2(new_n898), .A3(new_n889), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n874), .A2(KEYINPUT53), .A3(new_n886), .A4(new_n887), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n901), .B1(KEYINPUT54), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n690), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n641), .B(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n907), .A2(new_n187), .A3(new_n710), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n805), .A2(new_n612), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n744), .A2(new_n745), .A3(new_n751), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT50), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n908), .A2(KEYINPUT50), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n909), .A2(new_n711), .A3(new_n766), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n761), .A2(new_n676), .A3(new_n750), .ZN(new_n919));
  OR3_X1    g733(.A1(new_n918), .A2(KEYINPUT118), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT118), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n624), .A2(new_n613), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n774), .A2(new_n700), .A3(new_n710), .A4(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n610), .A2(new_n653), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n920), .A2(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n840), .A2(new_n842), .B1(new_n476), .B2(new_n847), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n912), .A2(new_n766), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT51), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n926), .B(KEYINPUT51), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n611), .B1(new_n911), .B2(new_n763), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n918), .A2(new_n858), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT48), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n933), .B(new_n935), .C1(new_n655), .C2(new_n923), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n905), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(G952), .A2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n851), .B1(new_n938), .B2(new_n939), .ZN(G75));
  AOI21_X1  g754(.A(new_n295), .B1(new_n902), .B2(new_n903), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(G210), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n255), .A2(new_n257), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n289), .ZN(new_n946));
  XOR2_X1   g760(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT120), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n946), .B(new_n948), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n287), .A2(G952), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n944), .A2(new_n949), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G51));
  INV_X1    g769(.A(KEYINPUT54), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n904), .B(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n478), .B(KEYINPUT57), .Z(new_n958));
  OAI21_X1  g772(.A(new_n519), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n941), .A2(new_n823), .A3(new_n820), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(G54));
  AND2_X1   g775(.A1(KEYINPUT58), .A2(G475), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n941), .A2(new_n600), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n600), .B1(new_n941), .B2(new_n962), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n951), .ZN(G60));
  XNOR2_X1  g779(.A(new_n649), .B(KEYINPUT121), .ZN(new_n966));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT59), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n905), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n952), .B1(new_n957), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(G63));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n672), .A2(new_n674), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n904), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n902), .B2(new_n903), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n952), .B1(new_n980), .B2(new_n395), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n973), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n904), .A2(new_n977), .ZN(new_n983));
  INV_X1    g797(.A(new_n395), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n980), .B2(new_n974), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n985), .A2(new_n987), .A3(KEYINPUT123), .A4(new_n952), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n978), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n980), .A2(KEYINPUT122), .A3(new_n974), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n991), .A2(new_n985), .A3(new_n952), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n986), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n994), .ZN(G66));
  NAND2_X1  g809(.A1(G224), .A2(G953), .ZN(new_n996));
  OAI22_X1  g810(.A1(new_n873), .A2(G953), .B1(new_n615), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n945), .B1(G898), .B2(new_n287), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n997), .B(new_n998), .Z(G69));
  NOR2_X1   g813(.A1(new_n858), .A2(new_n754), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n835), .B1(new_n815), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n860), .ZN(new_n1002));
  NOR4_X1   g816(.A1(new_n1002), .A2(new_n773), .A3(new_n797), .A4(new_n876), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n845), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT124), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n845), .A2(new_n1001), .A3(new_n1003), .A4(KEYINPUT124), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1006), .A2(new_n287), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n460), .A2(new_n461), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n593), .A2(new_n594), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(G900), .B2(G953), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n693), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1014), .A2(new_n766), .A3(new_n473), .A4(new_n864), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n815), .B2(new_n835), .ZN(new_n1017));
  OAI21_X1  g831(.A(KEYINPUT62), .B1(new_n703), .B2(new_n876), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n701), .A2(new_n696), .A3(new_n700), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n907), .A2(new_n694), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1020), .A2(new_n764), .A3(new_n1021), .A4(new_n883), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n845), .A2(new_n1017), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1011), .B1(new_n1024), .B2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1013), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(G900), .ZN(new_n1027));
  OAI21_X1  g841(.A(G953), .B1(new_n493), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT125), .Z(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1013), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(G72));
  INV_X1    g847(.A(new_n697), .ZN(new_n1034));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  NAND2_X1  g850(.A1(new_n464), .A2(new_n456), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n890), .B2(new_n899), .ZN(new_n1039));
  INV_X1    g853(.A(new_n873), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n845), .A2(new_n1017), .A3(new_n1040), .A4(new_n1023), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1034), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1042));
  NOR3_X1   g856(.A1(new_n1039), .A2(new_n1042), .A3(new_n951), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1006), .A2(new_n1040), .A3(new_n1007), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n1044), .A2(new_n1036), .ZN(new_n1045));
  OAI211_X1 g859(.A(KEYINPUT126), .B(new_n1043), .C1(new_n1045), .C2(new_n1037), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT126), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1042), .A2(new_n951), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1039), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1037), .B1(new_n1044), .B2(new_n1036), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1046), .A2(new_n1052), .ZN(G57));
endmodule


