

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573;

  XNOR2_X1 U318 ( .A(n498), .B(KEYINPUT48), .ZN(n524) );
  XOR2_X1 U319 ( .A(n315), .B(n314), .Z(n286) );
  XNOR2_X1 U320 ( .A(n526), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U321 ( .A(n528), .B(n527), .ZN(n555) );
  XNOR2_X1 U322 ( .A(n316), .B(n286), .ZN(n317) );
  XNOR2_X1 U323 ( .A(n318), .B(n317), .ZN(n323) );
  XNOR2_X1 U324 ( .A(n537), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U325 ( .A(n563), .B(n460), .ZN(n539) );
  XNOR2_X1 U326 ( .A(n423), .B(n422), .ZN(n535) );
  XNOR2_X1 U327 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n435) );
  XOR2_X1 U328 ( .A(G8GAT), .B(G197GAT), .Z(n288) );
  XNOR2_X1 U329 ( .A(G141GAT), .B(G22GAT), .ZN(n287) );
  XNOR2_X1 U330 ( .A(n288), .B(n287), .ZN(n292) );
  XOR2_X1 U331 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n290) );
  XNOR2_X1 U332 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U334 ( .A(n292), .B(n291), .Z(n297) );
  XOR2_X1 U335 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n294) );
  NAND2_X1 U336 ( .A1(G229GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U338 ( .A(KEYINPUT66), .B(n295), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U340 ( .A(G36GAT), .B(G50GAT), .Z(n300) );
  XNOR2_X1 U341 ( .A(G15GAT), .B(G1GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n298), .B(KEYINPUT72), .ZN(n347) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(n347), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U345 ( .A(n302), .B(n301), .Z(n308) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(KEYINPUT70), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n303), .B(G29GAT), .ZN(n304) );
  XOR2_X1 U348 ( .A(n304), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U349 ( .A(KEYINPUT7), .B(KEYINPUT71), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n327) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(n327), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n559) );
  XOR2_X1 U353 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n310) );
  XNOR2_X1 U354 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n313) );
  XOR2_X1 U356 ( .A(KEYINPUT13), .B(G57GAT), .Z(n312) );
  XNOR2_X1 U357 ( .A(G71GAT), .B(G78GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n339) );
  XOR2_X1 U359 ( .A(n313), .B(n339), .Z(n318) );
  XOR2_X1 U360 ( .A(G106GAT), .B(G148GAT), .Z(n357) );
  XOR2_X1 U361 ( .A(G99GAT), .B(G85GAT), .Z(n329) );
  XNOR2_X1 U362 ( .A(n357), .B(n329), .ZN(n316) );
  XOR2_X1 U363 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n315) );
  NAND2_X1 U364 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XOR2_X1 U365 ( .A(KEYINPUT76), .B(G64GAT), .Z(n320) );
  XNOR2_X1 U366 ( .A(G176GAT), .B(G92GAT), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U368 ( .A(G204GAT), .B(n321), .Z(n396) );
  XNOR2_X1 U369 ( .A(n396), .B(KEYINPUT32), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n563) );
  NAND2_X1 U371 ( .A1(n559), .A2(n563), .ZN(n447) );
  XOR2_X1 U372 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n325) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n336) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n328), .B(G218GAT), .ZN(n399) );
  XOR2_X1 U378 ( .A(n399), .B(n329), .Z(n331) );
  NAND2_X1 U379 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U381 ( .A(n332), .B(G92GAT), .Z(n334) );
  XOR2_X1 U382 ( .A(G50GAT), .B(G162GAT), .Z(n361) );
  XNOR2_X1 U383 ( .A(G134GAT), .B(n361), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n487) );
  INV_X1 U386 ( .A(n487), .ZN(n551) );
  XOR2_X1 U387 ( .A(KEYINPUT12), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U388 ( .A(G127GAT), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U390 ( .A(n339), .B(KEYINPUT14), .Z(n341) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n351) );
  XOR2_X1 U394 ( .A(G8GAT), .B(G183GAT), .Z(n395) );
  XOR2_X1 U395 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n345) );
  XNOR2_X1 U396 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U398 ( .A(n395), .B(n346), .Z(n349) );
  XOR2_X1 U399 ( .A(G22GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U400 ( .A(n347), .B(n358), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n567) );
  INV_X1 U403 ( .A(n567), .ZN(n492) );
  NOR2_X1 U404 ( .A1(n551), .A2(n492), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n352), .B(KEYINPUT16), .ZN(n433) );
  XOR2_X1 U406 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n354) );
  XNOR2_X1 U407 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n387) );
  XOR2_X1 U409 ( .A(G211GAT), .B(KEYINPUT90), .Z(n356) );
  XNOR2_X1 U410 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n405) );
  XNOR2_X1 U412 ( .A(n387), .B(n405), .ZN(n372) );
  XOR2_X1 U413 ( .A(n358), .B(n357), .Z(n360) );
  NAND2_X1 U414 ( .A1(G228GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U416 ( .A(n362), .B(n361), .Z(n370) );
  XOR2_X1 U417 ( .A(KEYINPUT24), .B(G78GAT), .Z(n364) );
  XNOR2_X1 U418 ( .A(G218GAT), .B(G204GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U420 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n366) );
  XNOR2_X1 U421 ( .A(KEYINPUT92), .B(KEYINPUT89), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n529) );
  XOR2_X1 U426 ( .A(n529), .B(KEYINPUT28), .Z(n481) );
  XOR2_X1 U427 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n374) );
  XNOR2_X1 U428 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n394) );
  XOR2_X1 U430 ( .A(G85GAT), .B(G148GAT), .Z(n376) );
  XNOR2_X1 U431 ( .A(G29GAT), .B(G162GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U433 ( .A(G57GAT), .B(KEYINPUT6), .Z(n378) );
  XNOR2_X1 U434 ( .A(G1GAT), .B(G155GAT), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U436 ( .A(n380), .B(n379), .Z(n392) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G127GAT), .Z(n382) );
  XNOR2_X1 U438 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U440 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n384) );
  XNOR2_X1 U441 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U443 ( .A(n386), .B(n385), .Z(n414) );
  XOR2_X1 U444 ( .A(n387), .B(KEYINPUT94), .Z(n389) );
  NAND2_X1 U445 ( .A1(G225GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n414), .B(n390), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n556) );
  XOR2_X1 U450 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U453 ( .A(n400), .B(n399), .Z(n407) );
  XNOR2_X1 U454 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n401), .B(KEYINPUT87), .ZN(n402) );
  XOR2_X1 U456 ( .A(n402), .B(KEYINPUT88), .Z(n404) );
  XNOR2_X1 U457 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n415) );
  XNOR2_X1 U459 ( .A(n415), .B(n405), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n523) );
  XNOR2_X1 U461 ( .A(n523), .B(KEYINPUT27), .ZN(n425) );
  NAND2_X1 U462 ( .A1(n556), .A2(n425), .ZN(n513) );
  NOR2_X1 U463 ( .A1(n481), .A2(n513), .ZN(n499) );
  XOR2_X1 U464 ( .A(KEYINPUT20), .B(G183GAT), .Z(n409) );
  XNOR2_X1 U465 ( .A(G190GAT), .B(G176GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U467 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n411) );
  XNOR2_X1 U468 ( .A(G15GAT), .B(G71GAT), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U470 ( .A(n413), .B(n412), .Z(n417) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n419) );
  NAND2_X1 U474 ( .A1(G227GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n423) );
  XNOR2_X1 U477 ( .A(G43GAT), .B(G99GAT), .ZN(n422) );
  INV_X1 U478 ( .A(n535), .ZN(n501) );
  NAND2_X1 U479 ( .A1(n499), .A2(n501), .ZN(n432) );
  NOR2_X1 U480 ( .A1(n529), .A2(n535), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n424), .B(KEYINPUT26), .ZN(n557) );
  NAND2_X1 U482 ( .A1(n425), .A2(n557), .ZN(n429) );
  NAND2_X1 U483 ( .A1(n535), .A2(n523), .ZN(n426) );
  NAND2_X1 U484 ( .A1(n529), .A2(n426), .ZN(n427) );
  XOR2_X1 U485 ( .A(KEYINPUT25), .B(n427), .Z(n428) );
  NAND2_X1 U486 ( .A1(n429), .A2(n428), .ZN(n430) );
  INV_X1 U487 ( .A(n556), .ZN(n530) );
  NAND2_X1 U488 ( .A1(n430), .A2(n530), .ZN(n431) );
  NAND2_X1 U489 ( .A1(n432), .A2(n431), .ZN(n443) );
  NAND2_X1 U490 ( .A1(n433), .A2(n443), .ZN(n462) );
  NOR2_X1 U491 ( .A1(n447), .A2(n462), .ZN(n440) );
  NAND2_X1 U492 ( .A1(n440), .A2(n556), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(G1324GAT) );
  XOR2_X1 U494 ( .A(G8GAT), .B(KEYINPUT95), .Z(n437) );
  NAND2_X1 U495 ( .A1(n440), .A2(n523), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(G1325GAT) );
  XOR2_X1 U497 ( .A(G15GAT), .B(KEYINPUT35), .Z(n439) );
  NAND2_X1 U498 ( .A1(n440), .A2(n535), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(G1326GAT) );
  NAND2_X1 U500 ( .A1(n440), .A2(n481), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n441), .B(KEYINPUT96), .ZN(n442) );
  XNOR2_X1 U502 ( .A(G22GAT), .B(n442), .ZN(G1327GAT) );
  XOR2_X1 U503 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n451) );
  XNOR2_X1 U504 ( .A(n487), .B(KEYINPUT36), .ZN(n571) );
  NAND2_X1 U505 ( .A1(n492), .A2(n443), .ZN(n444) );
  NOR2_X1 U506 ( .A1(n571), .A2(n444), .ZN(n446) );
  XOR2_X1 U507 ( .A(KEYINPUT97), .B(KEYINPUT37), .Z(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n476) );
  NOR2_X1 U509 ( .A1(n476), .A2(n447), .ZN(n449) );
  XNOR2_X1 U510 ( .A(KEYINPUT98), .B(KEYINPUT38), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n458), .A2(n556), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U514 ( .A(G29GAT), .B(n452), .Z(G1328GAT) );
  NAND2_X1 U515 ( .A1(n458), .A2(n523), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n453), .B(KEYINPUT100), .ZN(n454) );
  XNOR2_X1 U517 ( .A(G36GAT), .B(n454), .ZN(G1329GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n456) );
  NAND2_X1 U519 ( .A1(n458), .A2(n535), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U521 ( .A(G43GAT), .B(n457), .ZN(G1330GAT) );
  NAND2_X1 U522 ( .A1(n458), .A2(n481), .ZN(n459) );
  XNOR2_X1 U523 ( .A(n459), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U524 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n460) );
  INV_X1 U525 ( .A(n559), .ZN(n461) );
  NAND2_X1 U526 ( .A1(n539), .A2(n461), .ZN(n475) );
  NOR2_X1 U527 ( .A1(n475), .A2(n462), .ZN(n463) );
  XNOR2_X1 U528 ( .A(KEYINPUT102), .B(n463), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n471), .A2(n556), .ZN(n464) );
  XNOR2_X1 U530 ( .A(n464), .B(KEYINPUT42), .ZN(n465) );
  XNOR2_X1 U531 ( .A(G57GAT), .B(n465), .ZN(G1332GAT) );
  XOR2_X1 U532 ( .A(G64GAT), .B(KEYINPUT103), .Z(n467) );
  NAND2_X1 U533 ( .A1(n523), .A2(n471), .ZN(n466) );
  XNOR2_X1 U534 ( .A(n467), .B(n466), .ZN(G1333GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n469) );
  NAND2_X1 U536 ( .A1(n535), .A2(n471), .ZN(n468) );
  XNOR2_X1 U537 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U538 ( .A(G71GAT), .B(n470), .ZN(G1334GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n473) );
  NAND2_X1 U540 ( .A1(n481), .A2(n471), .ZN(n472) );
  XNOR2_X1 U541 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U542 ( .A(G78GAT), .B(n474), .ZN(G1335GAT) );
  NOR2_X1 U543 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U544 ( .A(KEYINPUT107), .B(n477), .Z(n482) );
  NAND2_X1 U545 ( .A1(n556), .A2(n482), .ZN(n478) );
  XNOR2_X1 U546 ( .A(n478), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U547 ( .A1(n482), .A2(n523), .ZN(n479) );
  XNOR2_X1 U548 ( .A(n479), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U549 ( .A1(n482), .A2(n535), .ZN(n480) );
  XNOR2_X1 U550 ( .A(n480), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U551 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n483), .B(KEYINPUT44), .ZN(n484) );
  XNOR2_X1 U553 ( .A(G106GAT), .B(n484), .ZN(G1339GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT108), .B(n567), .ZN(n546) );
  INV_X1 U555 ( .A(KEYINPUT46), .ZN(n486) );
  NAND2_X1 U556 ( .A1(n559), .A2(n539), .ZN(n485) );
  XOR2_X1 U557 ( .A(n486), .B(n485), .Z(n488) );
  NAND2_X1 U558 ( .A1(n488), .A2(n487), .ZN(n489) );
  OR2_X1 U559 ( .A1(n546), .A2(n489), .ZN(n490) );
  XNOR2_X1 U560 ( .A(n490), .B(KEYINPUT109), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n491), .B(KEYINPUT47), .ZN(n497) );
  NOR2_X1 U562 ( .A1(n492), .A2(n571), .ZN(n493) );
  XOR2_X1 U563 ( .A(KEYINPUT45), .B(n493), .Z(n494) );
  NOR2_X1 U564 ( .A1(n559), .A2(n494), .ZN(n495) );
  NAND2_X1 U565 ( .A1(n495), .A2(n563), .ZN(n496) );
  NAND2_X1 U566 ( .A1(n497), .A2(n496), .ZN(n498) );
  NAND2_X1 U567 ( .A1(n524), .A2(n499), .ZN(n500) );
  NOR2_X1 U568 ( .A1(n501), .A2(n500), .ZN(n509) );
  NAND2_X1 U569 ( .A1(n509), .A2(n559), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n502), .B(KEYINPUT110), .ZN(n503) );
  XNOR2_X1 U571 ( .A(G113GAT), .B(n503), .ZN(G1340GAT) );
  XOR2_X1 U572 ( .A(G120GAT), .B(KEYINPUT49), .Z(n505) );
  NAND2_X1 U573 ( .A1(n509), .A2(n539), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n505), .B(n504), .ZN(G1341GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT111), .B(KEYINPUT50), .Z(n507) );
  NAND2_X1 U576 ( .A1(n509), .A2(n546), .ZN(n506) );
  XNOR2_X1 U577 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U578 ( .A(G127GAT), .B(n508), .ZN(G1342GAT) );
  XOR2_X1 U579 ( .A(G134GAT), .B(KEYINPUT51), .Z(n511) );
  NAND2_X1 U580 ( .A1(n509), .A2(n551), .ZN(n510) );
  XNOR2_X1 U581 ( .A(n511), .B(n510), .ZN(G1343GAT) );
  NAND2_X1 U582 ( .A1(n524), .A2(n557), .ZN(n512) );
  NOR2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n520) );
  NAND2_X1 U584 ( .A1(n520), .A2(n559), .ZN(n514) );
  XNOR2_X1 U585 ( .A(n514), .B(KEYINPUT112), .ZN(n515) );
  XNOR2_X1 U586 ( .A(G141GAT), .B(n515), .ZN(G1344GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n517) );
  NAND2_X1 U588 ( .A1(n520), .A2(n539), .ZN(n516) );
  XNOR2_X1 U589 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U590 ( .A(G148GAT), .B(n518), .ZN(G1345GAT) );
  NAND2_X1 U591 ( .A1(n520), .A2(n567), .ZN(n519) );
  XNOR2_X1 U592 ( .A(n519), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U593 ( .A(G162GAT), .B(KEYINPUT113), .Z(n522) );
  NAND2_X1 U594 ( .A1(n520), .A2(n551), .ZN(n521) );
  XNOR2_X1 U595 ( .A(n522), .B(n521), .ZN(G1347GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n533) );
  XNOR2_X1 U597 ( .A(KEYINPUT114), .B(n523), .ZN(n525) );
  NAND2_X1 U598 ( .A1(n525), .A2(n524), .ZN(n528) );
  XOR2_X1 U599 ( .A(KEYINPUT54), .B(KEYINPUT115), .Z(n526) );
  NAND2_X1 U600 ( .A1(n530), .A2(n529), .ZN(n531) );
  OR2_X1 U601 ( .A1(n555), .A2(n531), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n534), .B(KEYINPUT55), .ZN(n536) );
  NAND2_X1 U604 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U605 ( .A1(n552), .A2(n559), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n538), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U607 ( .A1(n552), .A2(n539), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n541) );
  XNOR2_X1 U609 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U611 ( .A(G176GAT), .B(KEYINPUT56), .Z(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1349GAT) );
  XOR2_X1 U614 ( .A(G183GAT), .B(KEYINPUT123), .Z(n548) );
  NAND2_X1 U615 ( .A1(n552), .A2(n546), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1350GAT) );
  XNOR2_X1 U617 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n549), .B(KEYINPUT124), .ZN(n550) );
  XOR2_X1 U619 ( .A(KEYINPUT125), .B(n550), .Z(n554) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1351GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n570) );
  INV_X1 U624 ( .A(n570), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n568), .A2(n559), .ZN(n562) );
  XOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT60), .Z(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT59), .B(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1352GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n565) );
  OR2_X1 U630 ( .A1(n570), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G204GAT), .B(n566), .ZN(G1353GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT62), .B(n572), .Z(n573) );
  XNOR2_X1 U637 ( .A(G218GAT), .B(n573), .ZN(G1355GAT) );
endmodule

