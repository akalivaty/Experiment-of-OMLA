//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT76), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G227), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT77), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n195), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G146), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n200), .B1(new_n205), .B2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n204), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G104), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(KEYINPUT78), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n216), .A2(new_n218), .A3(new_n211), .A4(G104), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n215), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(G104), .B1(new_n216), .B2(new_n218), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n214), .A2(G107), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n210), .A2(KEYINPUT79), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n224), .A2(new_n221), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT79), .B1(new_n227), .B2(new_n210), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n202), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n207), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n196), .A2(new_n198), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n207), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n204), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n226), .A2(new_n228), .B1(new_n233), .B2(new_n227), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(G137), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT11), .A3(G134), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n237), .A2(new_n240), .A3(new_n243), .A4(new_n238), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n234), .A2(KEYINPUT12), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n199), .A2(new_n201), .B1(G128), .B2(new_n208), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n224), .A2(new_n221), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n233), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n253), .A2(new_n225), .B1(new_n254), .B2(new_n252), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n242), .A2(new_n244), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n247), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n246), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n226), .B2(new_n228), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n216), .A2(new_n218), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n211), .A2(G104), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT3), .B1(new_n214), .B2(G107), .ZN(new_n263));
  OAI22_X1  g077(.A1(new_n261), .A2(new_n262), .B1(new_n223), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G101), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n266));
  INV_X1    g080(.A(new_n230), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n205), .B2(G143), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n268), .A2(new_n271), .B1(new_n206), .B2(new_n269), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n264), .A2(new_n273), .A3(G101), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n233), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n260), .A2(new_n277), .A3(new_n256), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n194), .B1(new_n258), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT10), .B1(new_n253), .B2(new_n225), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n276), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n245), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n193), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT80), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT80), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n280), .A2(new_n281), .A3(new_n245), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n246), .B2(new_n257), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n287), .B(new_n284), .C1(new_n289), .C2(new_n194), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(G469), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT12), .B1(new_n234), .B2(new_n245), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n255), .A2(new_n247), .A3(new_n256), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n278), .B(new_n283), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n278), .A2(new_n282), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n193), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n294), .B1(new_n300), .B2(new_n292), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n189), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT90), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G140), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n306), .A2(new_n308), .A3(new_n309), .A4(KEYINPUT16), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT16), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT69), .B1(new_n306), .B2(KEYINPUT16), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n308), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT19), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT19), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n313), .A2(G146), .B1(new_n319), .B2(new_n205), .ZN(new_n320));
  INV_X1    g134(.A(G237), .ZN(new_n321));
  INV_X1    g135(.A(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G214), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(new_n207), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  AOI21_X1  g139(.A(G143), .B1(new_n325), .B2(G214), .ZN(new_n326));
  OAI21_X1  g140(.A(G131), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n207), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n243), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT71), .B1(new_n231), .B2(new_n314), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n205), .A2(new_n317), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n314), .A2(G146), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(KEYINPUT18), .A2(G131), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n328), .A2(new_n329), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n328), .B2(new_n329), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n320), .A2(new_n331), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G113), .B(G122), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(new_n214), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT88), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n346));
  INV_X1    g160(.A(new_n344), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n313), .A2(G146), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n319), .A2(new_n205), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n348), .A2(new_n331), .A3(new_n349), .ZN(new_n350));
  AOI211_X1 g164(.A(new_n340), .B(new_n339), .C1(new_n335), .C2(new_n336), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n346), .B(new_n347), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT17), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n327), .A2(new_n353), .A3(new_n330), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n195), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT17), .B(G131), .C1(new_n324), .C2(new_n326), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n348), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n337), .A2(new_n341), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n344), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n345), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G475), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n293), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT89), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n304), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n357), .A2(new_n358), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n347), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n366), .B2(new_n359), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n361), .B1(new_n367), .B2(KEYINPUT91), .ZN(new_n368));
  INV_X1    g182(.A(new_n359), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n344), .B1(new_n357), .B2(new_n358), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n293), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n303), .A2(new_n364), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n187), .A2(new_n375), .A3(G953), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n207), .A2(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n202), .A2(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G134), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n236), .ZN(new_n381));
  INV_X1    g195(.A(new_n261), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G122), .ZN(new_n384));
  INV_X1    g198(.A(G122), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G116), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n383), .A2(G122), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(new_n390), .C1(new_n384), .C2(KEYINPUT14), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(G116), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n386), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT92), .B1(new_n390), .B2(KEYINPUT14), .ZN(new_n395));
  OAI211_X1 g209(.A(G107), .B(new_n391), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT13), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n202), .B2(G143), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n378), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n377), .A2(new_n398), .ZN(new_n401));
  OAI21_X1  g215(.A(G134), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n382), .A2(new_n387), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n261), .A2(new_n384), .A3(new_n386), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n402), .B(new_n381), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n376), .B1(new_n397), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n397), .A2(new_n405), .A3(new_n376), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT93), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n405), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT93), .ZN(new_n411));
  INV_X1    g225(.A(new_n376), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n293), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G478), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(KEYINPUT15), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n414), .B(new_n416), .Z(new_n417));
  NAND2_X1  g231(.A1(new_n360), .A2(new_n363), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT90), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n360), .A2(new_n304), .A3(new_n363), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT20), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G952), .ZN(new_n422));
  AOI211_X1 g236(.A(G953), .B(new_n422), .C1(G234), .C2(G237), .ZN(new_n423));
  INV_X1    g237(.A(G898), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n322), .B1(KEYINPUT21), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(KEYINPUT21), .B2(new_n424), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n293), .B1(G234), .B2(G237), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n374), .A2(new_n417), .A3(new_n421), .A4(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G214), .B1(G237), .B2(G902), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n268), .A2(new_n271), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n199), .A2(new_n201), .A3(new_n269), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G125), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(G125), .B2(new_n233), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT83), .B(G224), .Z(new_n438));
  OAI21_X1  g252(.A(KEYINPUT7), .B1(new_n438), .B2(G953), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G119), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G116), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n383), .A2(G119), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT2), .B(G113), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n446), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n266), .A2(new_n450), .A3(new_n274), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT5), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G113), .B1(new_n442), .B2(KEYINPUT5), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n453), .A2(new_n455), .B1(new_n447), .B2(new_n445), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n227), .A2(KEYINPUT81), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n448), .B1(new_n452), .B2(new_n454), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n252), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n451), .A2(new_n457), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n439), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n436), .B(new_n463), .C1(G125), .C2(new_n233), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n440), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n452), .B1(new_n455), .B2(KEYINPUT85), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(KEYINPUT85), .B2(new_n455), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n448), .A3(new_n227), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n459), .A2(new_n252), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(KEYINPUT86), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(KEYINPUT86), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n461), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(G902), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n451), .A2(new_n457), .A3(new_n460), .ZN(new_n477));
  INV_X1    g291(.A(new_n461), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT82), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n462), .A3(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n477), .B(new_n478), .C1(new_n480), .C2(new_n481), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n438), .A2(G953), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n437), .B(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n476), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n476), .B2(new_n487), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n432), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n431), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n302), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n375), .B1(G234), .B2(new_n293), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT73), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT22), .B(G137), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G110), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n506));
  OAI211_X1 g320(.A(G119), .B(new_n202), .C1(new_n506), .C2(KEYINPUT23), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n441), .B2(G128), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT68), .B1(new_n441), .B2(G128), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n505), .B(new_n507), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(G119), .B(G128), .Z(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT24), .B(G110), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n506), .B1(G119), .B2(new_n202), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(KEYINPUT70), .A3(new_n505), .A4(new_n507), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n348), .A3(new_n335), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n313), .A2(G146), .B1(new_n332), .B2(new_n334), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n521), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n441), .A2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n508), .A2(KEYINPUT68), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n517), .A2(new_n518), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n530), .A2(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n348), .B2(new_n355), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n504), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n504), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n532), .B(new_n535), .C1(new_n523), .C2(new_n526), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n293), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT25), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n524), .A2(new_n525), .A3(new_n521), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n525), .B1(new_n524), .B2(new_n521), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n533), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n535), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n527), .A2(new_n533), .A3(new_n504), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT25), .A3(new_n293), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n500), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n499), .A2(G902), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT75), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT25), .B1(new_n545), .B2(new_n293), .ZN(new_n553));
  AOI211_X1 g367(.A(new_n538), .B(G902), .C1(new_n543), .C2(new_n544), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n499), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT75), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n550), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G472), .ZN(new_n559));
  INV_X1    g373(.A(new_n238), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n236), .A2(G137), .ZN(new_n561));
  OAI21_X1  g375(.A(G131), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n244), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n233), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n450), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n245), .A2(new_n433), .A3(new_n434), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT65), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(KEYINPUT65), .ZN(new_n572));
  INV_X1    g386(.A(new_n567), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT1), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n205), .B2(G143), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n268), .B1(new_n575), .B2(new_n202), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n563), .B1(new_n576), .B2(new_n204), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n565), .A2(KEYINPUT65), .A3(new_n569), .A4(new_n567), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n568), .B1(new_n580), .B2(new_n450), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT26), .B(G101), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n325), .A2(G210), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT67), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n245), .A2(new_n272), .B1(new_n233), .B2(new_n564), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT28), .B1(new_n588), .B2(new_n566), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n450), .B1(new_n573), .B2(new_n577), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n589), .B1(new_n592), .B2(KEYINPUT28), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT29), .B1(new_n593), .B2(new_n586), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT67), .ZN(new_n595));
  INV_X1    g409(.A(new_n586), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n566), .B1(new_n578), .B2(new_n579), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n568), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n587), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT28), .B1(new_n568), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n589), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n596), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n604), .B2(KEYINPUT29), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n559), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT31), .ZN(new_n607));
  NOR4_X1   g421(.A1(new_n597), .A2(new_n607), .A3(new_n568), .A4(new_n596), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT31), .B1(new_n603), .B2(new_n596), .ZN(new_n609));
  INV_X1    g423(.A(new_n572), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n570), .B(new_n610), .C1(new_n565), .C2(new_n567), .ZN(new_n611));
  AND4_X1   g425(.A1(KEYINPUT65), .A2(new_n565), .A3(new_n569), .A4(new_n567), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n450), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n591), .A3(new_n586), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n608), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT32), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n559), .A4(new_n293), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT28), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n590), .B2(new_n591), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n596), .B1(new_n619), .B2(new_n589), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n614), .A2(new_n607), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n581), .A2(KEYINPUT31), .A3(new_n586), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(new_n559), .A3(new_n293), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT32), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n606), .B1(new_n617), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n558), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n302), .A2(new_n495), .A3(KEYINPUT94), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n498), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  NAND2_X1  g443(.A1(new_n291), .A2(new_n301), .ZN(new_n630));
  INV_X1    g444(.A(new_n189), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n621), .A2(new_n293), .A3(new_n622), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n623), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n632), .A2(new_n558), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n409), .A2(new_n413), .A3(new_n637), .ZN(new_n638));
  OR3_X1    g452(.A1(new_n410), .A2(KEYINPUT96), .A3(new_n412), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n408), .B1(new_n406), .B2(KEYINPUT96), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT33), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n638), .A2(new_n641), .A3(G478), .A4(new_n293), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n414), .A2(new_n415), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT97), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n645), .A2(new_n647), .B1(new_n374), .B2(new_n421), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n476), .A2(new_n487), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n488), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n476), .A2(new_n487), .A3(new_n489), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n432), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n649), .A2(new_n429), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n636), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  XNOR2_X1  g471(.A(new_n414), .B(new_n416), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n374), .A2(new_n421), .A3(new_n658), .A4(new_n430), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT98), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n651), .A2(new_n432), .A3(new_n652), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n659), .A2(KEYINPUT98), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n636), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NOR2_X1   g481(.A1(new_n504), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n542), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n549), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n555), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n635), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n498), .A2(new_n627), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  INV_X1    g491(.A(new_n606), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n623), .A2(KEYINPUT32), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n623), .A2(KEYINPUT32), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n661), .A3(new_n671), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n374), .A2(new_n421), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT99), .ZN(new_n684));
  INV_X1    g498(.A(new_n428), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n322), .A2(G900), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n423), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n428), .A2(KEYINPUT99), .A3(new_n686), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n683), .A2(new_n417), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n302), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n677), .B1(new_n682), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n625), .A2(new_n653), .A3(new_n672), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n302), .A2(new_n693), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT100), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT101), .B(G128), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G30));
  NOR2_X1   g515(.A1(new_n492), .A2(new_n493), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n432), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n417), .B1(new_n374), .B2(new_n421), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n617), .A2(new_n624), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n581), .A2(new_n596), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n293), .B1(new_n592), .B2(new_n586), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n671), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n691), .B(KEYINPUT39), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT40), .B1(new_n302), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n302), .A2(KEYINPUT40), .A3(new_n714), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n708), .B(new_n713), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G143), .ZN(G45));
  NAND2_X1  g532(.A1(new_n647), .A2(new_n645), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n683), .A3(new_n691), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n632), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n696), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  OR2_X1    g537(.A1(new_n300), .A2(new_n292), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n297), .A2(new_n299), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n292), .A3(new_n293), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n631), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n654), .A2(new_n626), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n664), .A2(new_n626), .A3(new_n728), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NOR2_X1   g547(.A1(new_n727), .A2(new_n431), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n696), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  NOR2_X1   g550(.A1(new_n707), .A2(new_n653), .ZN(new_n737));
  NOR2_X1   g551(.A1(G472), .A2(G902), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT103), .ZN(new_n739));
  AOI22_X1  g553(.A1(G472), .A2(new_n633), .B1(new_n615), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n547), .A2(new_n551), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(new_n728), .A3(new_n742), .A4(new_n430), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n671), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n720), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n661), .A3(new_n728), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  INV_X1    g562(.A(new_n741), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n625), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n720), .ZN(new_n751));
  INV_X1    g565(.A(new_n294), .ZN(new_n752));
  OAI211_X1 g566(.A(G469), .B(new_n284), .C1(new_n289), .C2(new_n194), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n726), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n492), .A2(new_n493), .A3(new_n705), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n754), .A2(new_n755), .A3(new_n631), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n750), .A2(KEYINPUT42), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n547), .A2(KEYINPUT75), .A3(new_n551), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n556), .B1(new_n555), .B2(new_n550), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n760), .A3(new_n681), .A4(new_n751), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n761), .A2(KEYINPUT104), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT104), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  NAND4_X1  g580(.A1(new_n756), .A2(new_n760), .A3(new_n681), .A4(new_n693), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  AND2_X1   g582(.A1(new_n374), .A2(new_n421), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n719), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT43), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n635), .A2(new_n671), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n755), .B1(new_n774), .B2(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT44), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n279), .A2(new_n780), .A3(new_n285), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT105), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n286), .A2(new_n290), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n292), .B1(new_n783), .B2(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(KEYINPUT106), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n752), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n790), .A2(new_n791), .B1(new_n292), .B2(new_n300), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n752), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n189), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n779), .A2(new_n794), .A3(new_n714), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  NOR2_X1   g610(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n794), .B1(new_n799), .B2(new_n797), .ZN(new_n800));
  INV_X1    g614(.A(new_n493), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n476), .A2(new_n487), .A3(new_n491), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n432), .A3(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n760), .A2(new_n681), .A3(new_n720), .A4(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n798), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  AND2_X1   g620(.A1(new_n772), .A2(new_n423), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n727), .A2(new_n803), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n750), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT48), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n809), .A2(KEYINPUT114), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n709), .A2(new_n712), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n808), .A2(new_n812), .A3(new_n760), .A4(new_n423), .ZN(new_n813));
  OAI211_X1 g627(.A(G952), .B(new_n322), .C1(new_n813), .C2(new_n649), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n807), .A2(new_n728), .A3(new_n742), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n817), .A2(KEYINPUT113), .A3(new_n661), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT113), .B1(new_n817), .B2(new_n661), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n811), .B(new_n816), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n813), .A2(new_n683), .A3(new_n719), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n807), .A2(new_n808), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n745), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n705), .A3(new_n704), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n724), .A2(new_n726), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n631), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n798), .B2(new_n800), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n807), .A2(new_n742), .A3(new_n755), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n820), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n828), .B(KEYINPUT51), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n661), .A2(new_n691), .A3(new_n706), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n754), .A2(new_n631), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n721), .A2(new_n696), .B1(new_n840), .B2(new_n713), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n682), .A2(new_n694), .A3(new_n677), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT100), .B1(new_n696), .B2(new_n697), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n747), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n648), .B1(new_n658), .B2(new_n769), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n494), .A2(new_n429), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n636), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n628), .A2(new_n674), .A3(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n803), .A2(new_n683), .A3(new_n658), .A4(new_n692), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n681), .A3(new_n302), .A4(new_n671), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT110), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n746), .B2(new_n756), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n648), .A2(new_n740), .A3(new_n671), .A4(new_n691), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n754), .A2(new_n755), .A3(new_n631), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT110), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n767), .B(new_n852), .C1(new_n854), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n699), .A2(new_n860), .A3(new_n747), .A4(new_n841), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n729), .A2(new_n732), .A3(new_n735), .A4(new_n743), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n765), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n765), .B2(new_n864), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n845), .A2(new_n861), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n628), .A2(new_n674), .A3(new_n849), .ZN(new_n871));
  INV_X1    g685(.A(new_n858), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n765), .A2(new_n864), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(KEYINPUT111), .B(new_n869), .C1(new_n870), .C2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n732), .A2(new_n729), .A3(new_n735), .A4(new_n743), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n761), .A2(new_n762), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT104), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n761), .A2(KEYINPUT104), .A3(new_n762), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n876), .B1(new_n881), .B2(new_n757), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n861), .A3(new_n845), .A4(new_n859), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT111), .B1(new_n883), .B2(new_n869), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n867), .B(new_n868), .C1(new_n875), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n869), .B1(new_n870), .B2(new_n873), .ZN(new_n886));
  INV_X1    g700(.A(new_n882), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(new_n862), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n837), .A2(new_n890), .B1(G952), .B2(G953), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n829), .B(KEYINPUT49), .Z(new_n892));
  NOR4_X1   g706(.A1(new_n770), .A2(new_n749), .A3(new_n189), .A4(new_n705), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n812), .A3(new_n704), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(G75));
  NOR3_X1   g709(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT111), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(new_n874), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n293), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(KEYINPUT115), .A3(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n483), .A2(new_n484), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n486), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT115), .B1(new_n900), .B2(G210), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n909), .A2(new_n905), .B1(G952), .B2(new_n322), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(G51));
  NOR2_X1   g725(.A1(new_n322), .A2(G952), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n867), .B1(new_n875), .B2(new_n884), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(G902), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n789), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n725), .B(KEYINPUT116), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n885), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n294), .B(KEYINPUT57), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n915), .B1(new_n920), .B2(KEYINPUT117), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n922));
  INV_X1    g736(.A(new_n919), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n917), .B2(new_n885), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n912), .B1(new_n921), .B2(new_n925), .ZN(G54));
  NAND2_X1  g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT118), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n899), .A2(new_n293), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT119), .B1(new_n929), .B2(new_n360), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n912), .B1(new_n929), .B2(new_n360), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  INV_X1    g746(.A(new_n360), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n932), .B(new_n933), .C1(new_n914), .C2(new_n928), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n930), .A2(new_n931), .A3(new_n937), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G60));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n890), .A2(new_n942), .B1(new_n641), .B2(new_n638), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n638), .A2(new_n641), .A3(new_n942), .ZN(new_n944));
  AOI211_X1 g758(.A(new_n912), .B(new_n943), .C1(new_n918), .C2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n545), .B1(new_n913), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n912), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n913), .A2(new_n669), .A3(new_n948), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n953), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n954), .A2(new_n950), .A3(new_n955), .ZN(new_n956));
  XOR2_X1   g770(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(G66));
  AOI21_X1  g772(.A(new_n427), .B1(G953), .B2(new_n438), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n850), .A2(new_n876), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n903), .B1(G898), .B2(new_n322), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT123), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n961), .B(new_n964), .ZN(G69));
  NAND4_X1  g779(.A1(new_n794), .A2(new_n714), .A3(new_n737), .A4(new_n750), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n765), .A2(new_n767), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n699), .A2(new_n722), .A3(new_n747), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n795), .A2(new_n805), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n322), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n580), .B(new_n319), .Z(new_n972));
  XNOR2_X1  g786(.A(new_n686), .B(KEYINPUT127), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n699), .A2(new_n717), .A3(new_n722), .A4(new_n747), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n302), .A2(new_n714), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n978), .A2(new_n846), .A3(new_n803), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n626), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n795), .A2(new_n805), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT125), .Z(new_n983));
  OAI211_X1 g797(.A(new_n322), .B(new_n972), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT126), .B1(new_n975), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n686), .B1(new_n191), .B2(G953), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  AOI211_X1 g802(.A(KEYINPUT126), .B(new_n986), .C1(new_n975), .C2(new_n984), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  INV_X1    g806(.A(new_n960), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n970), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n581), .A3(new_n596), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n587), .A2(new_n614), .A3(new_n598), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n992), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n912), .B1(new_n888), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n981), .A2(new_n983), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n992), .B1(new_n1000), .B2(new_n993), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n999), .B1(new_n710), .B2(new_n1001), .ZN(G57));
endmodule


