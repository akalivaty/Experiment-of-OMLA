//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OR3_X1    g0010(.A1(new_n210), .A2(KEYINPUT64), .A3(G13), .ZN(new_n211));
  OAI21_X1  g0011(.A(KEYINPUT64), .B1(new_n210), .B2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n206), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n208), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n217), .A2(KEYINPUT0), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(KEYINPUT0), .B2(new_n217), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n216), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G97), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n215), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n210), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n223), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  NAND2_X1  g0044(.A1(G68), .A2(G77), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n203), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  OAI21_X1  g0053(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n257), .A3(G274), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n254), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G222), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G223), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n257), .B1(new_n271), .B2(new_n202), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n261), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G200), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(G190), .B2(new_n273), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n208), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT68), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT8), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n280), .A2(KEYINPUT67), .A3(G58), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G50), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n229), .A3(new_n201), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n286), .A2(G20), .B1(G150), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n218), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n289), .A2(new_n292), .B1(G50), .B2(new_n293), .ZN(new_n294));
  OR3_X1    g0094(.A1(new_n208), .A2(KEYINPUT69), .A3(G1), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT69), .B1(new_n208), .B2(G1), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n285), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n293), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n291), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT9), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n294), .A2(KEYINPUT9), .A3(new_n303), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n276), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT73), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n306), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n304), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n313), .A2(new_n308), .A3(KEYINPUT10), .A4(new_n276), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n294), .A2(new_n303), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT71), .A2(G179), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT71), .A2(G179), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n273), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G169), .B2(new_n273), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G20), .A2(G77), .ZN(new_n323));
  INV_X1    g0123(.A(new_n287), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n323), .B1(new_n282), .B2(new_n324), .C1(new_n277), .C2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n291), .B1(new_n202), .B2(new_n300), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n295), .A2(new_n296), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n301), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G77), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n262), .A2(G232), .A3(new_n264), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n226), .B2(new_n262), .ZN(new_n335));
  INV_X1    g0135(.A(G238), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n271), .A2(new_n336), .A3(new_n264), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n333), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G274), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n333), .A2(new_n339), .A3(new_n254), .ZN(new_n340));
  INV_X1    g0140(.A(new_n259), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(G244), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n332), .B1(new_n344), .B2(G169), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n319), .B2(new_n344), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n332), .B1(G200), .B2(new_n343), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(KEYINPUT72), .B1(G190), .B2(new_n344), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n331), .B(new_n327), .C1(new_n344), .C2(new_n274), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT72), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n346), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n315), .A2(new_n322), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n279), .A2(G77), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n354), .B1(new_n208), .B2(G68), .C1(new_n285), .C2(new_n324), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n300), .A2(new_n201), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT12), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n330), .A2(G68), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT11), .B1(new_n355), .B2(new_n291), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n260), .A2(new_n264), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n230), .A2(G1698), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n262), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G97), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n257), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n258), .B1(new_n259), .B2(new_n336), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT13), .B1(new_n367), .B2(new_n369), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n372), .A2(G190), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT74), .A4(new_n371), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n376), .A2(G200), .A3(new_n377), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n362), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(G169), .A3(new_n377), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n372), .A2(new_n373), .A3(G179), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n376), .A2(new_n385), .A3(G169), .A4(new_n377), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n386), .A2(KEYINPUT75), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(KEYINPUT75), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n381), .B(new_n384), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n379), .B1(new_n389), .B2(new_n362), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n262), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n201), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n229), .A2(new_n201), .ZN(new_n397));
  NOR2_X1   g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n287), .A2(G159), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n392), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT78), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT77), .B1(new_n267), .B2(G33), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT77), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(new_n269), .A3(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n406), .A3(new_n268), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n208), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n393), .A3(new_n208), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(G68), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n401), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(KEYINPUT16), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT78), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n392), .C1(new_n396), .C2(new_n401), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n403), .A2(new_n413), .A3(new_n291), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n329), .A2(new_n283), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n300), .B2(new_n283), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n340), .B1(G232), .B2(new_n341), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT79), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n260), .A2(G1698), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(G223), .B2(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n423), .B1(new_n407), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n333), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n319), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G169), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n419), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT18), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n419), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n274), .B1(new_n420), .B2(new_n427), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(G190), .B2(new_n428), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n416), .A2(new_n438), .A3(new_n418), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n416), .A2(new_n438), .A3(KEYINPUT17), .A4(new_n418), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n434), .A2(new_n436), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n353), .A2(new_n391), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT90), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G116), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G20), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT23), .B1(new_n226), .B2(G20), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n404), .A2(new_n406), .A3(new_n208), .A4(new_n268), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT22), .A2(G87), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n208), .A2(G87), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n271), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT89), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(KEYINPUT89), .C1(new_n453), .C2(new_n454), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n452), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT24), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n458), .B1(new_n453), .B2(new_n454), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT89), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n460), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n452), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n292), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT25), .B1(new_n300), .B2(new_n226), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n207), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n293), .A2(new_n474), .A3(new_n218), .A4(new_n290), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n472), .A2(new_n473), .B1(G107), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n446), .B1(new_n470), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n468), .B1(new_n467), .B2(new_n452), .ZN(new_n480));
  INV_X1    g0280(.A(new_n452), .ZN(new_n481));
  AOI211_X1 g0281(.A(KEYINPUT24), .B(new_n481), .C1(new_n466), .C2(new_n460), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n291), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(KEYINPUT90), .A3(new_n477), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n215), .A2(G1698), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(G250), .B2(G1698), .ZN(new_n486));
  INV_X1    g0286(.A(G294), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n407), .A2(new_n486), .B1(new_n269), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT5), .B(G41), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n333), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n488), .A2(new_n333), .B1(new_n492), .B2(G264), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n491), .A2(new_n257), .A3(G274), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G179), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(G169), .B2(new_n495), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n479), .A2(new_n484), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n208), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT85), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(KEYINPUT85), .A3(new_n208), .ZN(new_n505));
  INV_X1    g0305(.A(G87), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n231), .A3(new_n226), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n277), .B2(new_n231), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n508), .B(new_n510), .C1(new_n201), .C2(new_n453), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n292), .B1(new_n511), .B2(KEYINPUT86), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n404), .A2(new_n406), .A3(new_n268), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n208), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT86), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n508), .A4(new_n510), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n512), .A2(new_n516), .B1(new_n300), .B2(new_n325), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n225), .A2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G238), .B2(G1698), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n447), .B1(new_n407), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n333), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n206), .B1(new_n489), .B2(G1), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n207), .A2(new_n339), .A3(G45), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n257), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n518), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n525), .ZN(new_n527));
  AOI211_X1 g0327(.A(KEYINPUT84), .B(new_n527), .C1(new_n521), .C2(new_n333), .ZN(new_n528));
  OAI21_X1  g0328(.A(G200), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n476), .A2(G87), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G238), .A2(G1698), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n225), .B2(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(new_n268), .A3(new_n404), .A4(new_n406), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n257), .B1(new_n533), .B2(new_n447), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT84), .B1(new_n534), .B2(new_n527), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n522), .A2(new_n518), .A3(new_n525), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(G190), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n517), .A2(new_n529), .A3(new_n530), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n510), .B1(new_n453), .B2(new_n201), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT86), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(new_n516), .A3(new_n291), .ZN(new_n542));
  INV_X1    g0342(.A(new_n325), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n476), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n325), .A2(new_n300), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n431), .B1(new_n526), .B2(new_n528), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n535), .A2(new_n536), .A3(new_n319), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G257), .A2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n216), .B2(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n552), .A2(new_n268), .A3(new_n404), .A4(new_n406), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n271), .A2(G303), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n333), .ZN(new_n556));
  AND2_X1   g0356(.A1(KEYINPUT5), .A2(G41), .ZN(new_n557));
  NOR2_X1   g0357(.A1(KEYINPUT5), .A2(G41), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n490), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(G270), .A3(new_n257), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n494), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n208), .A2(G116), .B1(KEYINPUT87), .B2(KEYINPUT20), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n292), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT80), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT80), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(G33), .A3(G283), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n208), .B1(new_n231), .B2(G33), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n565), .B(new_n566), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G20), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n291), .B(new_n576), .C1(KEYINPUT87), .C2(KEYINPUT20), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n568), .B2(new_n570), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT87), .B(KEYINPUT20), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n293), .A2(new_n575), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n476), .B2(new_n575), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n563), .A2(new_n582), .A3(G169), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n257), .B1(new_n553), .B2(new_n554), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n585), .A2(new_n496), .A3(new_n561), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n583), .A2(new_n584), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT88), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n563), .A2(new_n582), .A3(KEYINPUT21), .A4(G169), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n556), .A2(new_n562), .A3(G190), .ZN(new_n591));
  OAI21_X1  g0391(.A(G200), .B1(new_n585), .B2(new_n561), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(G169), .B1(new_n585), .B2(new_n561), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n584), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n586), .A2(new_n582), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n593), .A3(new_n589), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT88), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n550), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n494), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n559), .A2(G257), .A3(new_n257), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n559), .A2(KEYINPUT81), .A3(G257), .A4(new_n257), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n225), .A2(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n404), .A2(new_n406), .A3(new_n268), .A4(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT4), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n268), .A2(new_n270), .A3(G250), .A4(G1698), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(KEYINPUT4), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n571), .C1(new_n271), .C2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n333), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n606), .A2(new_n614), .A3(new_n319), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT83), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n606), .A2(new_n614), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n431), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT6), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n619), .A2(new_n231), .A3(G107), .ZN(new_n620));
  XNOR2_X1  g0420(.A(G97), .B(G107), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n622), .A2(new_n208), .B1(new_n202), .B2(new_n324), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n226), .B1(new_n394), .B2(new_n395), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n291), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n293), .A2(G97), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n476), .B2(G97), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT83), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n606), .A2(new_n614), .A3(new_n629), .A4(new_n319), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n616), .A2(new_n618), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n625), .A2(new_n627), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n617), .A2(G200), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n606), .A2(new_n614), .A3(G190), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT82), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n635), .A2(KEYINPUT82), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G190), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n495), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(G200), .B2(new_n495), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n483), .A3(new_n477), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n500), .A2(new_n600), .A3(new_n638), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n445), .A2(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n522), .A2(new_n525), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n517), .A2(new_n530), .A3(new_n537), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n431), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n546), .A2(new_n548), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n463), .A2(new_n469), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n478), .B1(new_n651), .B2(new_n291), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n652), .B2(new_n641), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n587), .A2(new_n589), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n652), .B2(new_n498), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n653), .A2(new_n638), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n647), .A2(new_n649), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n616), .A2(new_n618), .A3(KEYINPUT91), .A4(new_n630), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n616), .A2(new_n630), .A3(new_n618), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT91), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n632), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n550), .B2(new_n631), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n649), .A3(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n444), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n322), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n419), .A2(new_n435), .A3(new_n432), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n435), .B1(new_n419), .B2(new_n432), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n379), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n672), .A2(new_n346), .B1(new_n389), .B2(new_n362), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n441), .A2(new_n442), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n671), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n668), .B1(new_n676), .B2(new_n315), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n594), .A2(new_n599), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n679), .B1(new_n590), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n654), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n582), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n479), .A2(new_n484), .A3(new_n685), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n500), .A2(new_n694), .A3(new_n642), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n500), .B2(new_n686), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n654), .A2(new_n685), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n500), .A2(new_n642), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n499), .B1(new_n470), .B2(new_n478), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n685), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT92), .ZN(G399));
  NOR2_X1   g0504(.A1(new_n214), .A2(G41), .ZN(new_n705));
  NOR4_X1   g0505(.A1(new_n705), .A2(new_n207), .A3(G116), .A4(new_n507), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n221), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  INV_X1    g0508(.A(KEYINPUT98), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n660), .A2(new_n661), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n628), .A3(new_n659), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT26), .B1(new_n711), .B2(new_n650), .ZN(new_n712));
  INV_X1    g0512(.A(new_n631), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n658), .A3(new_n549), .A4(new_n538), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(new_n649), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT97), .ZN(new_n716));
  INV_X1    g0516(.A(new_n642), .ZN(new_n717));
  NOR4_X1   g0517(.A1(new_n717), .A2(new_n636), .A3(new_n637), .A4(new_n650), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n500), .A2(new_n654), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n715), .A2(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n712), .A2(KEYINPUT97), .A3(new_n649), .A4(new_n714), .ZN(new_n721));
  AOI211_X1 g0521(.A(new_n709), .B(new_n685), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n715), .A2(new_n716), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n719), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT98), .B1(new_n725), .B2(new_n686), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT29), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n666), .A2(new_n686), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n617), .A2(new_n495), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n429), .B1(new_n556), .B2(new_n562), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n534), .A2(KEYINPUT93), .A3(new_n527), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n522), .B2(new_n525), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT93), .B1(new_n534), .B2(new_n527), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n522), .A2(new_n737), .A3(new_n525), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n735), .B1(new_n743), .B2(new_n734), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n733), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n586), .A2(new_n493), .A3(new_n614), .A4(new_n606), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n535), .A2(new_n536), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT95), .ZN(new_n750));
  OR3_X1    g0550(.A1(new_n747), .A2(new_n746), .A3(new_n748), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT95), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n752), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n745), .A2(new_n750), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n685), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n745), .A2(new_n751), .A3(new_n749), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n757), .B(new_n759), .C1(new_n643), .C2(new_n685), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G330), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n732), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n708), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT101), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n431), .A2(KEYINPUT102), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n208), .B1(KEYINPUT102), .B2(new_n431), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n218), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n213), .A2(new_n407), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n249), .A2(G45), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT100), .Z(new_n775));
  AOI211_X1 g0575(.A(new_n773), .B(new_n775), .C1(new_n489), .C2(new_n221), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n213), .A2(new_n262), .ZN(new_n777));
  INV_X1    g0577(.A(G355), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n778), .B1(G116), .B2(new_n213), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n772), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G13), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n207), .B1(new_n782), .B2(G45), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n705), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n208), .A2(new_n274), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n429), .A2(G190), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT104), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(KEYINPUT104), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT103), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n208), .A2(new_n639), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n429), .A2(new_n274), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n208), .A2(G190), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n429), .A2(new_n274), .A3(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n229), .A2(new_n796), .B1(new_n798), .B2(new_n202), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n793), .A2(G50), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n795), .A2(new_n496), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G179), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G190), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n262), .B1(new_n801), .B2(new_n506), .C1(new_n805), .C2(new_n231), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n797), .A2(new_n496), .A3(G200), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT106), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT106), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n226), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n429), .A2(new_n639), .A3(new_n787), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n806), .B(new_n811), .C1(G68), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n797), .A2(new_n802), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G159), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT105), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT32), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n799), .A2(new_n794), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n800), .A2(new_n814), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n810), .ZN(new_n822));
  INV_X1    g0622(.A(new_n798), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n822), .A2(G283), .B1(new_n823), .B2(G311), .ZN(new_n824));
  INV_X1    g0624(.A(G329), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n271), .B1(new_n815), .B2(new_n825), .C1(new_n801), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G294), .B2(new_n804), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT107), .B(G326), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n824), .B(new_n828), .C1(new_n792), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G322), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT33), .B(G317), .Z(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n796), .B1(new_n812), .B2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT108), .Z(new_n834));
  OAI21_X1  g0634(.A(new_n821), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n786), .B1(new_n835), .B2(new_n771), .ZN(new_n836));
  INV_X1    g0636(.A(new_n767), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n780), .B(new_n836), .C1(new_n690), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n690), .A2(G330), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n786), .B1(new_n691), .B2(new_n692), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n346), .A2(new_n686), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n686), .B1(new_n327), .B2(new_n331), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n348), .B2(new_n351), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n346), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n728), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n686), .B(new_n848), .C1(new_n656), .C2(new_n665), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n762), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT109), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n847), .A2(new_n849), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n786), .C1(new_n762), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n766), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n771), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n786), .B1(new_n202), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n771), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n822), .A2(G87), .ZN(new_n858));
  INV_X1    g0658(.A(new_n796), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G283), .A2(new_n813), .B1(new_n859), .B2(G294), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n860), .C1(new_n575), .C2(new_n798), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n792), .A2(new_n826), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n805), .A2(new_n231), .ZN(new_n863));
  INV_X1    g0663(.A(G311), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n271), .B1(new_n815), .B2(new_n864), .C1(new_n801), .C2(new_n226), .ZN(new_n865));
  NOR4_X1   g0665(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G143), .A2(new_n859), .B1(new_n813), .B2(G150), .ZN(new_n867));
  INV_X1    g0667(.A(G159), .ZN(new_n868));
  INV_X1    g0668(.A(G137), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n868), .B2(new_n798), .C1(new_n792), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT34), .ZN(new_n871));
  INV_X1    g0671(.A(G132), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n513), .B1(new_n872), .B2(new_n815), .C1(new_n285), .C2(new_n801), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n810), .A2(new_n201), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n873), .B(new_n874), .C1(G58), .C2(new_n804), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n866), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n856), .B1(new_n857), .B2(new_n876), .C1(new_n848), .C2(new_n766), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n853), .A2(new_n877), .ZN(G384));
  NOR2_X1   g0678(.A1(new_n782), .A2(new_n207), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n727), .A2(new_n444), .A3(new_n730), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n677), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT112), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n419), .A2(new_n432), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n419), .B2(new_n432), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n683), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n419), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(KEYINPUT113), .B(KEYINPUT37), .Z(new_n890));
  AND3_X1   g0690(.A1(new_n889), .A2(new_n439), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n413), .A2(new_n291), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT16), .B1(new_n411), .B2(new_n412), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n418), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n432), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n888), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(new_n439), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n887), .A2(new_n891), .B1(KEYINPUT37), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n671), .B2(new_n674), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n882), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n433), .A2(KEYINPUT112), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n439), .A2(new_n890), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(new_n889), .A4(new_n884), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n896), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n443), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT75), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n386), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n384), .A2(new_n381), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n362), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n362), .A2(new_n685), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n672), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n362), .B(new_n685), .C1(new_n389), .C2(new_n379), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n849), .A2(KEYINPUT111), .A3(new_n843), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT111), .B1(new_n849), .B2(new_n843), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n909), .B(new_n917), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n671), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n683), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n433), .A2(new_n889), .A3(new_n439), .ZN(new_n923));
  INV_X1    g0723(.A(new_n890), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n903), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n889), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n443), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n882), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n908), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n913), .A2(new_n685), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n920), .A2(new_n922), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n881), .B(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n757), .B(new_n939), .C1(new_n643), .C2(new_n685), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n846), .B1(new_n915), .B2(new_n916), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n905), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n926), .B2(new_n928), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT40), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n909), .A2(new_n946), .A3(new_n940), .A4(new_n941), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n940), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n445), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n948), .A2(new_n950), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n952), .A2(new_n953), .A3(new_n692), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n879), .B1(new_n938), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n938), .B2(new_n955), .ZN(new_n957));
  INV_X1    g0757(.A(new_n622), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(G116), .A3(new_n219), .A4(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n201), .A2(G50), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT110), .Z(new_n964));
  NOR3_X1   g0764(.A1(new_n397), .A2(new_n220), .A3(new_n202), .ZN(new_n965));
  OAI211_X1 g0765(.A(G1), .B(new_n781), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n957), .A2(new_n962), .A3(new_n966), .ZN(G367));
  NOR2_X1   g0767(.A1(new_n239), .A2(new_n773), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n772), .B1(new_n213), .B2(new_n325), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n785), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n822), .A2(G97), .B1(G294), .B2(new_n813), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n826), .B2(new_n796), .ZN(new_n972));
  INV_X1    g0772(.A(new_n801), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n801), .B2(new_n575), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(new_n226), .C2(new_n805), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  INV_X1    g0778(.A(G283), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n407), .B1(new_n978), .B2(new_n815), .C1(new_n798), .C2(new_n979), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n972), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n793), .A2(G311), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n793), .A2(G143), .ZN(new_n983));
  INV_X1    g0783(.A(G150), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n810), .A2(new_n202), .B1(new_n984), .B2(new_n796), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n805), .A2(new_n201), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n262), .B1(new_n815), .B2(new_n869), .C1(new_n801), .C2(new_n229), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n285), .A2(new_n798), .B1(new_n812), .B2(new_n868), .ZN(new_n988));
  NOR4_X1   g0788(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n981), .A2(new_n982), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT47), .Z(new_n991));
  AOI21_X1  g0791(.A(new_n970), .B1(new_n991), .B2(new_n771), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n517), .A2(new_n530), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n685), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n657), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n649), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n992), .B1(new_n837), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n700), .B1(new_n696), .B2(new_n699), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n693), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n731), .A2(new_n761), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n711), .A2(new_n686), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n628), .A2(new_n685), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1002), .B1(new_n638), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n702), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT44), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n702), .A2(new_n1004), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n698), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n697), .A3(new_n1008), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n763), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n705), .B(KEYINPUT41), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n784), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n631), .B1(new_n1004), .B2(new_n500), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n686), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT42), .B1(new_n1004), .B2(new_n700), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT115), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1004), .A2(KEYINPUT42), .A3(new_n700), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(KEYINPUT115), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(KEYINPUT114), .A2(KEYINPUT43), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(KEYINPUT114), .A2(KEYINPUT43), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n997), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT43), .B2(new_n997), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1022), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n697), .A2(new_n1004), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1031), .B(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n998), .B1(new_n1016), .B2(new_n1034), .ZN(G387));
  OR2_X1    g0835(.A1(new_n696), .A2(new_n837), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n243), .A2(new_n489), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n507), .A2(G116), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1037), .A2(new_n773), .B1(new_n1038), .B2(new_n777), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n282), .A2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1041), .A2(new_n489), .A3(new_n245), .A4(new_n1038), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1039), .A2(new_n1042), .B1(new_n226), .B2(new_n214), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n772), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n785), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n793), .A2(G159), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n973), .A2(G77), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n984), .B2(new_n815), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n805), .A2(new_n325), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n407), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n822), .A2(G97), .B1(G50), .B2(new_n859), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G68), .A2(new_n823), .B1(new_n813), .B2(new_n283), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1046), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n805), .A2(new_n979), .B1(new_n801), .B2(new_n487), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G303), .A2(new_n823), .B1(new_n813), .B2(G311), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n978), .B2(new_n796), .C1(new_n792), .C2(new_n831), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT48), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n407), .B1(new_n829), .B2(new_n815), .C1(new_n810), .C2(new_n575), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1053), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1045), .B1(new_n1063), .B2(new_n771), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1000), .A2(new_n784), .B1(new_n1036), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n763), .A2(new_n1000), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1001), .A2(new_n705), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(G393));
  INV_X1    g0868(.A(new_n1012), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n784), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1004), .A2(new_n767), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n772), .B1(new_n231), .B2(new_n213), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n213), .A2(new_n252), .A3(new_n407), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n785), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n858), .B1(new_n285), .B2(new_n812), .C1(new_n282), .C2(new_n798), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n805), .A2(new_n202), .ZN(new_n1076));
  INV_X1    g0876(.A(G143), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n801), .A2(new_n201), .B1(new_n815), .B2(new_n1077), .ZN(new_n1078));
  OR4_X1    g0878(.A1(new_n407), .A2(new_n1075), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n792), .A2(new_n984), .B1(new_n868), .B2(new_n796), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  AOI22_X1  g0881(.A1(new_n793), .A2(G317), .B1(G311), .B2(new_n859), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n271), .B1(new_n815), .B2(new_n831), .C1(new_n801), .C2(new_n979), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G116), .B2(new_n804), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n813), .A2(G303), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n811), .B1(G294), .B2(new_n823), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1079), .A2(new_n1081), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1074), .B1(new_n1091), .B2(new_n771), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1071), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1070), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n705), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1001), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1069), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1012), .A2(new_n1001), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n940), .A2(G330), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n444), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n880), .A2(new_n677), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n725), .A2(new_n686), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n709), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n725), .A2(KEYINPUT98), .A3(new_n686), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n1108), .A3(new_n843), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n845), .A2(new_n346), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n760), .A2(G330), .A3(new_n848), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n917), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1101), .B2(new_n846), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1102), .A2(new_n941), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n919), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n849), .A2(KEYINPUT111), .A3(new_n843), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1119), .A2(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1105), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1115), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT38), .B1(new_n905), .B2(new_n907), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n942), .A2(new_n1128), .A3(new_n932), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT39), .B1(new_n930), .B2(new_n908), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n934), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1109), .A2(new_n1111), .A3(new_n917), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n934), .B1(new_n930), .B2(new_n908), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1127), .B(new_n1134), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1134), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1119), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1126), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1119), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1136), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n722), .A2(new_n726), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1110), .B1(new_n1144), .B2(new_n843), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n917), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1142), .B1(new_n1146), .B2(new_n1134), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1138), .A2(new_n1139), .A3(new_n1115), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1123), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1104), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1141), .A2(new_n1151), .A3(new_n705), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n855), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n785), .B1(new_n283), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT118), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1131), .A2(new_n766), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n271), .B1(new_n801), .B2(new_n506), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n823), .A2(G97), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1076), .B(new_n874), .C1(G294), .C2(new_n816), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n226), .B2(new_n812), .C1(new_n575), .C2(new_n796), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G283), .C2(new_n793), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n801), .A2(new_n984), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n271), .B1(new_n816), .B2(G125), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n868), .C2(new_n805), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G132), .A2(new_n859), .B1(new_n813), .B2(G137), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT54), .B(G143), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1169), .B1(new_n285), .B2(new_n810), .C1(new_n798), .C2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1168), .B(new_n1171), .C1(G128), .C2(new_n793), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1163), .A2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1155), .B(new_n1156), .C1(new_n771), .C2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n784), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1152), .A2(new_n1176), .ZN(G378));
  NAND3_X1  g0977(.A1(new_n311), .A2(new_n314), .A3(new_n322), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n316), .A2(new_n683), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n311), .A2(new_n314), .A3(new_n322), .A4(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n854), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n793), .A2(G116), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1047), .B1(new_n979), .B2(new_n815), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n513), .A2(G41), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1189), .A2(new_n986), .A3(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G97), .A2(new_n813), .B1(new_n859), .B2(G107), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n822), .A2(G58), .B1(new_n823), .B2(new_n543), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1188), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  INV_X1    g0995(.A(G41), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G50), .B1(new_n269), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1194), .A2(new_n1195), .B1(new_n1190), .B2(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G33), .B(G41), .C1(new_n816), .C2(G124), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n859), .B1(new_n823), .B2(G137), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1170), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n973), .A2(new_n1201), .B1(new_n804), .B2(G150), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(new_n872), .C2(new_n812), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G125), .B2(new_n793), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT59), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1199), .B1(new_n868), .B2(new_n810), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1204), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1198), .B1(new_n1195), .B2(new_n1194), .C1(new_n1206), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n771), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n855), .A2(new_n285), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1187), .A2(new_n785), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1186), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n948), .B2(G330), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n692), .B(new_n1186), .C1(new_n945), .C2(new_n947), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n937), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n940), .A2(new_n941), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT40), .B1(new_n900), .B2(new_n908), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(KEYINPUT40), .A2(new_n944), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1186), .B1(new_n1220), .B2(new_n692), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n946), .B1(new_n1218), .B2(new_n931), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n946), .B1(new_n942), .B2(new_n1128), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n940), .A2(new_n941), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G330), .B(new_n1214), .C1(new_n1222), .C2(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1131), .A2(new_n934), .B1(new_n921), .B2(new_n683), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1221), .A2(new_n920), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1217), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1213), .B1(new_n1229), .B2(new_n784), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1104), .B1(new_n1175), .B2(new_n1150), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(KEYINPUT57), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n705), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1148), .B1(new_n1234), .B2(new_n1119), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1105), .B1(new_n1235), .B2(new_n1126), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1229), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1230), .B1(new_n1233), .B2(new_n1237), .ZN(G375));
  NAND2_X1  g1038(.A1(new_n1104), .A2(new_n1149), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1126), .A2(new_n1015), .A3(new_n1239), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n783), .B(KEYINPUT121), .Z(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1114), .A2(new_n854), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n785), .B1(G68), .B2(new_n1153), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n793), .A2(G294), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n271), .B1(new_n815), .B2(new_n826), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1246), .B(new_n1049), .C1(G97), .C2(new_n973), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n822), .A2(G77), .B1(G116), .B2(new_n813), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G107), .A2(new_n823), .B1(new_n859), .B2(G283), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n792), .A2(new_n872), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT122), .ZN(new_n1252));
  INV_X1    g1052(.A(G128), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n801), .A2(new_n868), .B1(new_n815), .B2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n407), .B(new_n1254), .C1(G50), .C2(new_n804), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n822), .A2(G58), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G137), .A2(new_n859), .B1(new_n823), .B2(G150), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n813), .A2(new_n1201), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1250), .B1(new_n1252), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1244), .B1(new_n1260), .B2(new_n771), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1125), .A2(new_n1242), .B1(new_n1243), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1240), .A2(new_n1262), .ZN(G381));
  INV_X1    g1063(.A(G375), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT123), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1152), .A2(new_n1176), .A3(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1099), .B(new_n998), .C1(new_n1016), .C2(new_n1034), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1264), .A2(new_n1268), .A3(new_n1270), .A4(new_n1271), .ZN(G407));
  NAND2_X1  g1072(.A1(new_n684), .A2(G213), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT124), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1264), .A2(new_n1268), .A3(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(G407), .A2(G213), .A3(new_n1275), .ZN(G409));
  XNOR2_X1  g1076(.A(G393), .B(G396), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G390), .A2(G387), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n1269), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1269), .A3(new_n1277), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1280), .A2(KEYINPUT127), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT127), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1236), .A2(new_n1015), .A3(new_n1229), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1215), .A2(new_n1216), .A3(new_n937), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1221), .A2(new_n1226), .B1(new_n1227), .B2(new_n920), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1242), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT125), .B1(new_n1288), .B2(new_n1212), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1241), .B1(new_n1217), .B2(new_n1228), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1213), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1285), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1265), .A2(new_n1267), .A3(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1230), .C1(new_n1233), .C2(new_n1237), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1239), .A2(KEYINPUT60), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT60), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1104), .A2(new_n1149), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n705), .B1(new_n1104), .B2(new_n1149), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(G384), .A3(new_n1262), .ZN(new_n1305));
  INV_X1    g1105(.A(G384), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1262), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1305), .A2(new_n1309), .A3(KEYINPUT126), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1297), .A2(new_n1273), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1274), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1315), .A2(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1305), .A2(new_n1309), .A3(KEYINPUT126), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT126), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1321), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1310), .A2(G2897), .A3(new_n1274), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1320), .B1(new_n1326), .B2(new_n1317), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1284), .B1(new_n1319), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1315), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1297), .A2(new_n1273), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1317), .A2(KEYINPUT63), .A3(new_n1314), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1280), .A2(new_n1320), .A3(new_n1281), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1330), .A2(new_n1332), .A3(new_n1333), .A4(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1328), .A2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(new_n1268), .A2(G375), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1296), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1314), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1310), .A3(new_n1296), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1284), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1339), .B(new_n1340), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(G402));
endmodule


