

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XOR2_X1 U324 ( .A(n431), .B(n430), .Z(n292) );
  XNOR2_X1 U325 ( .A(n476), .B(KEYINPUT48), .ZN(n477) );
  XNOR2_X1 U326 ( .A(n478), .B(n477), .ZN(n536) );
  XNOR2_X1 U327 ( .A(n298), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U328 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n480) );
  XNOR2_X1 U329 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U330 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U331 ( .A(n419), .B(KEYINPUT37), .ZN(n420) );
  NAND2_X1 U332 ( .A1(n397), .A2(n396), .ZN(n494) );
  XNOR2_X1 U333 ( .A(n421), .B(n420), .ZN(n522) );
  XNOR2_X1 U334 ( .A(KEYINPUT123), .B(n487), .ZN(n571) );
  INV_X1 U335 ( .A(KEYINPUT40), .ZN(n457) );
  XNOR2_X1 U336 ( .A(n488), .B(G176GAT), .ZN(n489) );
  XNOR2_X1 U337 ( .A(n457), .B(G43GAT), .ZN(n458) );
  XNOR2_X1 U338 ( .A(n490), .B(n489), .ZN(G1349GAT) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(G1330GAT) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(G134GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n293), .B(G99GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n294), .B(G120GAT), .ZN(n387) );
  XOR2_X1 U344 ( .A(n295), .B(n387), .Z(n302) );
  XOR2_X1 U345 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n297) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n341) );
  XOR2_X1 U348 ( .A(n341), .B(G15GAT), .Z(n300) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n311) );
  XOR2_X1 U351 ( .A(G183GAT), .B(G127GAT), .Z(n304) );
  XNOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n309) );
  INV_X1 U354 ( .A(G71GAT), .ZN(n305) );
  XOR2_X1 U355 ( .A(G71GAT), .B(G176GAT), .Z(n307) );
  XNOR2_X1 U356 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U358 ( .A(n309), .B(n308), .Z(n310) );
  XOR2_X1 U359 ( .A(n311), .B(n310), .Z(n312) );
  XOR2_X1 U360 ( .A(KEYINPUT36), .B(KEYINPUT101), .Z(n329) );
  XOR2_X1 U361 ( .A(G36GAT), .B(G190GAT), .Z(n332) );
  XOR2_X1 U362 ( .A(G99GAT), .B(G85GAT), .Z(n424) );
  XOR2_X1 U363 ( .A(n332), .B(n424), .Z(n314) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G218GAT), .Z(n352) );
  XOR2_X1 U365 ( .A(G29GAT), .B(G134GAT), .Z(n386) );
  XNOR2_X1 U366 ( .A(n352), .B(n386), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n320) );
  XOR2_X1 U368 ( .A(G43GAT), .B(KEYINPUT8), .Z(n316) );
  XNOR2_X1 U369 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n446) );
  XOR2_X1 U371 ( .A(G92GAT), .B(n446), .Z(n318) );
  NAND2_X1 U372 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U375 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n322) );
  XNOR2_X1 U376 ( .A(KEYINPUT10), .B(KEYINPUT78), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U378 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n324) );
  XNOR2_X1 U379 ( .A(G162GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U381 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n464) );
  XNOR2_X1 U383 ( .A(n329), .B(n464), .ZN(n589) );
  XOR2_X1 U384 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n331) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U387 ( .A(n333), .B(n332), .Z(n335) );
  XOR2_X1 U388 ( .A(G197GAT), .B(KEYINPUT21), .Z(n351) );
  XNOR2_X1 U389 ( .A(G218GAT), .B(n351), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U391 ( .A(G8GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n336), .B(G211GAT), .ZN(n404) );
  XOR2_X1 U393 ( .A(n337), .B(n404), .Z(n343) );
  XOR2_X1 U394 ( .A(G92GAT), .B(G64GAT), .Z(n339) );
  XNOR2_X1 U395 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U397 ( .A(G176GAT), .B(n340), .Z(n435) );
  XNOR2_X1 U398 ( .A(n341), .B(n435), .ZN(n342) );
  XOR2_X1 U399 ( .A(n343), .B(n342), .Z(n527) );
  XNOR2_X1 U400 ( .A(n527), .B(KEYINPUT27), .ZN(n394) );
  INV_X1 U401 ( .A(n312), .ZN(n539) );
  XOR2_X1 U402 ( .A(KEYINPUT86), .B(KEYINPUT3), .Z(n345) );
  XNOR2_X1 U403 ( .A(G162GAT), .B(KEYINPUT87), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U405 ( .A(n346), .B(KEYINPUT2), .Z(n348) );
  XNOR2_X1 U406 ( .A(G141GAT), .B(G155GAT), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n391) );
  XOR2_X1 U408 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n350) );
  XNOR2_X1 U409 ( .A(G22GAT), .B(G204GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n356) );
  XOR2_X1 U411 ( .A(G211GAT), .B(KEYINPUT88), .Z(n354) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U415 ( .A1(G228GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U417 ( .A(n359), .B(KEYINPUT22), .Z(n363) );
  XOR2_X1 U418 ( .A(G78GAT), .B(G148GAT), .Z(n361) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n427) );
  XNOR2_X1 U421 ( .A(n427), .B(KEYINPUT85), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n391), .B(n364), .ZN(n484) );
  NOR2_X1 U424 ( .A1(n539), .A2(n484), .ZN(n366) );
  XNOR2_X1 U425 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n365) );
  XOR2_X1 U426 ( .A(n366), .B(n365), .Z(n552) );
  NOR2_X1 U427 ( .A1(n394), .A2(n552), .ZN(n367) );
  XNOR2_X1 U428 ( .A(KEYINPUT97), .B(n367), .ZN(n373) );
  XNOR2_X1 U429 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n371) );
  INV_X1 U430 ( .A(n527), .ZN(n479) );
  NAND2_X1 U431 ( .A1(n479), .A2(n539), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n368), .B(KEYINPUT98), .ZN(n369) );
  NAND2_X1 U433 ( .A1(n369), .A2(n484), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  NAND2_X1 U435 ( .A1(n373), .A2(n372), .ZN(n392) );
  XOR2_X1 U436 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n375) );
  XNOR2_X1 U437 ( .A(G148GAT), .B(G85GAT), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U439 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n377) );
  XNOR2_X1 U440 ( .A(KEYINPUT90), .B(G57GAT), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U442 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U443 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n381) );
  NAND2_X1 U444 ( .A1(G225GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U446 ( .A(KEYINPUT92), .B(n382), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U448 ( .A(G1GAT), .B(G127GAT), .Z(n403) );
  XOR2_X1 U449 ( .A(n385), .B(n403), .Z(n389) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U452 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U453 ( .A1(n392), .A2(n393), .ZN(n397) );
  XOR2_X1 U454 ( .A(KEYINPUT93), .B(n393), .Z(n524) );
  NOR2_X1 U455 ( .A1(n524), .A2(n394), .ZN(n537) );
  XNOR2_X1 U456 ( .A(KEYINPUT28), .B(n484), .ZN(n533) );
  INV_X1 U457 ( .A(n533), .ZN(n541) );
  NOR2_X1 U458 ( .A1(n539), .A2(n541), .ZN(n395) );
  NAND2_X1 U459 ( .A1(n537), .A2(n395), .ZN(n396) );
  XNOR2_X1 U460 ( .A(G22GAT), .B(G15GAT), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n398), .B(KEYINPUT71), .ZN(n445) );
  INV_X1 U462 ( .A(G57GAT), .ZN(n399) );
  NAND2_X1 U463 ( .A1(G71GAT), .A2(n399), .ZN(n401) );
  NAND2_X1 U464 ( .A1(n305), .A2(G57GAT), .ZN(n400) );
  NAND2_X1 U465 ( .A1(n401), .A2(n400), .ZN(n402) );
  XOR2_X1 U466 ( .A(KEYINPUT13), .B(n402), .Z(n422) );
  XNOR2_X1 U467 ( .A(n445), .B(n422), .ZN(n417) );
  XOR2_X1 U468 ( .A(n404), .B(n403), .Z(n406) );
  XNOR2_X1 U469 ( .A(G155GAT), .B(G78GAT), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U471 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n408) );
  NAND2_X1 U472 ( .A1(G231GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U474 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U475 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n412) );
  XNOR2_X1 U476 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n413), .B(KEYINPUT14), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n491) );
  NAND2_X1 U481 ( .A1(n494), .A2(n491), .ZN(n418) );
  NOR2_X1 U482 ( .A1(n589), .A2(n418), .ZN(n421) );
  INV_X1 U483 ( .A(KEYINPUT102), .ZN(n419) );
  INV_X1 U484 ( .A(KEYINPUT31), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n426) );
  XNOR2_X1 U486 ( .A(G120GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n427), .B(KEYINPUT76), .ZN(n429) );
  AND2_X1 U489 ( .A1(G230GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U491 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n433) );
  XNOR2_X1 U492 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n292), .B(n436), .ZN(n460) );
  XOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n438) );
  XNOR2_X1 U497 ( .A(G113GAT), .B(G1GAT), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n454) );
  XOR2_X1 U499 ( .A(G141GAT), .B(G197GAT), .Z(n440) );
  XNOR2_X1 U500 ( .A(G169GAT), .B(G50GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U502 ( .A(G36GAT), .B(G29GAT), .Z(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n450) );
  XNOR2_X1 U504 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n443), .B(G8GAT), .ZN(n444) );
  XOR2_X1 U506 ( .A(n444), .B(KEYINPUT69), .Z(n448) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n452) );
  NAND2_X1 U510 ( .A1(G229GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n579) );
  NOR2_X1 U513 ( .A1(n460), .A2(n579), .ZN(n495) );
  NAND2_X1 U514 ( .A1(n522), .A2(n495), .ZN(n455) );
  XOR2_X1 U515 ( .A(KEYINPUT103), .B(n455), .Z(n456) );
  XNOR2_X1 U516 ( .A(KEYINPUT38), .B(n456), .ZN(n508) );
  NOR2_X1 U517 ( .A1(n312), .A2(n508), .ZN(n459) );
  INV_X1 U518 ( .A(n524), .ZN(n483) );
  XOR2_X1 U519 ( .A(KEYINPUT112), .B(n491), .Z(n568) );
  INV_X1 U520 ( .A(n579), .ZN(n565) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT64), .ZN(n462) );
  INV_X1 U522 ( .A(KEYINPUT41), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n462), .B(n461), .ZN(n557) );
  NAND2_X1 U524 ( .A1(n565), .A2(n557), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT46), .B(n463), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n568), .A2(n466), .ZN(n467) );
  XNOR2_X1 U528 ( .A(KEYINPUT47), .B(n467), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n491), .A2(n589), .ZN(n469) );
  XNOR2_X1 U530 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U532 ( .A(KEYINPUT65), .B(n470), .Z(n471) );
  NOR2_X1 U533 ( .A1(n460), .A2(n471), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n472), .B(KEYINPUT114), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n473), .A2(n579), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n478) );
  INV_X1 U537 ( .A(KEYINPUT115), .ZN(n476) );
  NAND2_X1 U538 ( .A1(n479), .A2(n536), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n483), .A2(n482), .ZN(n578) );
  NAND2_X1 U540 ( .A1(n578), .A2(n484), .ZN(n485) );
  XNOR2_X1 U541 ( .A(n485), .B(KEYINPUT55), .ZN(n486) );
  NAND2_X1 U542 ( .A1(n486), .A2(n539), .ZN(n487) );
  NAND2_X1 U543 ( .A1(n571), .A2(n557), .ZN(n490) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n488) );
  INV_X1 U545 ( .A(n491), .ZN(n586) );
  NAND2_X1 U546 ( .A1(n464), .A2(n586), .ZN(n492) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n492), .Z(n493) );
  AND2_X1 U548 ( .A1(n494), .A2(n493), .ZN(n513) );
  NAND2_X1 U549 ( .A1(n495), .A2(n513), .ZN(n502) );
  NOR2_X1 U550 ( .A1(n524), .A2(n502), .ZN(n496) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(n496), .Z(n497) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n497), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n527), .A2(n502), .ZN(n498) );
  XOR2_X1 U554 ( .A(KEYINPUT100), .B(n498), .Z(n499) );
  XNOR2_X1 U555 ( .A(G8GAT), .B(n499), .ZN(G1325GAT) );
  NOR2_X1 U556 ( .A1(n312), .A2(n502), .ZN(n501) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n501), .B(n500), .ZN(G1326GAT) );
  NOR2_X1 U559 ( .A1(n533), .A2(n502), .ZN(n503) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n503), .Z(G1327GAT) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n506) );
  NOR2_X1 U562 ( .A1(n508), .A2(n524), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT104), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n508), .A2(n527), .ZN(n507) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n507), .Z(G1329GAT) );
  XNOR2_X1 U567 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n510) );
  NOR2_X1 U568 ( .A1(n533), .A2(n508), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  NAND2_X1 U571 ( .A1(n557), .A2(n579), .ZN(n512) );
  XNOR2_X1 U572 ( .A(n512), .B(KEYINPUT107), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n523), .A2(n513), .ZN(n518) );
  NOR2_X1 U574 ( .A1(n524), .A2(n518), .ZN(n514) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n514), .Z(n515) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n515), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n527), .A2(n518), .ZN(n516) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n516), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n312), .A2(n518), .ZN(n517) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n533), .A2(n518), .ZN(n520) );
  XNOR2_X1 U582 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n522), .ZN(n532) );
  NOR2_X1 U586 ( .A1(n524), .A2(n532), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n527), .A2(n532), .ZN(n528) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n528), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n312), .A2(n532), .ZN(n529) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n531) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n535) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U597 ( .A(n535), .B(n534), .Z(G1339GAT) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(n538), .Z(n553) );
  NAND2_X1 U600 ( .A1(n539), .A2(n553), .ZN(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n548), .A2(n565), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U605 ( .A1(n548), .A2(n557), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n546) );
  NAND2_X1 U608 ( .A1(n548), .A2(n568), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n550) );
  INV_X1 U612 ( .A(n464), .ZN(n572) );
  NAND2_X1 U613 ( .A1(n548), .A2(n572), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT120), .ZN(n556) );
  INV_X1 U617 ( .A(n552), .ZN(n577) );
  NAND2_X1 U618 ( .A1(n577), .A2(n553), .ZN(n554) );
  XNOR2_X1 U619 ( .A(KEYINPUT119), .B(n554), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n565), .A2(n562), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U623 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n586), .A2(n562), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U628 ( .A(G162GAT), .B(KEYINPUT121), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n572), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n565), .A2(n571), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT125), .Z(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT58), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n588) );
  NOR2_X1 U644 ( .A1(n579), .A2(n588), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U647 ( .A(n588), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n585), .A2(n460), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

