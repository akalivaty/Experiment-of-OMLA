//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(G127gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n204), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n202), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n203), .A2(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT68), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT27), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G183gat), .ZN(new_n222));
  AND4_X1   g021(.A1(KEYINPUT68), .A2(new_n220), .A3(new_n222), .A4(new_n217), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n215), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n222), .A3(new_n217), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n216), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n214), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(G169gat), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT26), .B1(new_n231), .B2(new_n232), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n224), .A2(new_n229), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n242), .A2(G169gat), .A3(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n236), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n242), .B1(G169gat), .B2(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n217), .ZN(new_n247));
  NAND3_X1  g046(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n247), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n250), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n245), .B(new_n246), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n243), .A2(KEYINPUT66), .A3(new_n244), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT23), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(new_n236), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n246), .A2(KEYINPUT25), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n247), .A2(new_n248), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT24), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n230), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n260), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n241), .A2(new_n254), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n213), .B1(new_n239), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G227gat), .ZN(new_n268));
  INV_X1    g067(.A(G233gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT66), .B1(new_n243), .B2(new_n244), .ZN(new_n271));
  INV_X1    g070(.A(new_n260), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(new_n247), .A3(new_n248), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n256), .A3(new_n236), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n246), .A3(new_n236), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n250), .B1(new_n230), .B2(new_n263), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n278), .B2(new_n252), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n275), .B1(new_n279), .B2(new_n240), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n224), .A2(new_n229), .A3(new_n238), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n208), .A2(new_n207), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n282), .B(new_n205), .C1(KEYINPUT1), .C2(new_n202), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n212), .A2(new_n208), .A3(new_n210), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n267), .A2(new_n270), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G71gat), .B(G99gat), .Z(new_n291));
  XNOR2_X1  g090(.A(G15gat), .B(G43gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT33), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT34), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n267), .A2(new_n286), .ZN(new_n301));
  INV_X1    g100(.A(new_n270), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g102(.A(KEYINPUT34), .B(new_n270), .C1(new_n267), .C2(new_n286), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n294), .A3(new_n298), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT36), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(KEYINPUT36), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G141gat), .ZN(new_n318));
  INV_X1    g117(.A(G148gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT2), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(KEYINPUT76), .A3(new_n321), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n317), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT77), .B1(new_n314), .B2(new_n315), .ZN(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(KEYINPUT2), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n327), .A2(new_n333), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT3), .B1(new_n326), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n323), .B1(new_n334), .B2(new_n335), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n325), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n316), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n338), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n346), .A3(new_n285), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n338), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n349), .A2(new_n285), .A3(KEYINPUT4), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n351));
  AND3_X1   g150(.A1(new_n327), .A2(new_n336), .A3(new_n337), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n352), .A2(new_n333), .B1(new_n343), .B2(new_n316), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n353), .B2(new_n213), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n347), .B(new_n348), .C1(new_n350), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n213), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n285), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n348), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n349), .B2(new_n285), .ZN(new_n363));
  INV_X1    g162(.A(new_n351), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n353), .A2(new_n213), .A3(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n363), .A2(new_n356), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n213), .B1(KEYINPUT3), .B2(new_n349), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n360), .B1(new_n367), .B2(new_n346), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n355), .A2(new_n361), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT80), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT6), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n361), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n366), .A2(new_n368), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G211gat), .A2(G218gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT22), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(G197gat), .A2(G204gat), .ZN(new_n388));
  AND2_X1   g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G211gat), .B(G218gat), .Z(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G197gat), .B(G204gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n387), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(KEYINPUT72), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT72), .B1(new_n392), .B2(new_n395), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT73), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n280), .A2(new_n281), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n401), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n280), .B2(new_n281), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n399), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n401), .ZN(new_n408));
  INV_X1    g207(.A(new_n398), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n396), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT29), .B1(new_n280), .B2(new_n281), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n408), .B(new_n410), .C1(new_n401), .C2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G64gat), .B(G92gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  NAND3_X1  g214(.A1(new_n407), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT75), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n407), .A2(KEYINPUT75), .A3(new_n412), .A4(new_n415), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n407), .B2(new_n412), .ZN(new_n422));
  INV_X1    g221(.A(new_n416), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n384), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT31), .B(G50gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n403), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n353), .B2(new_n345), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n434), .B2(new_n410), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n392), .A2(new_n395), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT3), .B1(new_n438), .B2(KEYINPUT83), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n392), .B2(new_n395), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n353), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT84), .B1(new_n435), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n346), .A2(new_n403), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n431), .B1(new_n445), .B2(new_n399), .ZN(new_n446));
  INV_X1    g245(.A(new_n442), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n345), .B1(new_n440), .B2(new_n441), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n349), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G22gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n434), .B2(new_n410), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n445), .A2(new_n399), .A3(KEYINPUT82), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n403), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n345), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n349), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n431), .B(KEYINPUT81), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n452), .A2(new_n453), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n453), .B1(new_n452), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n430), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n450), .B1(new_n446), .B2(new_n449), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n461), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n445), .A2(new_n399), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n470), .A2(new_n454), .B1(new_n349), .B2(new_n458), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n471), .B2(new_n456), .ZN(new_n472));
  OAI21_X1  g271(.A(G22gat), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n453), .A3(new_n462), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n429), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n313), .B1(new_n426), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n415), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n407), .A2(new_n412), .ZN(new_n481));
  INV_X1    g280(.A(new_n415), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n410), .B1(new_n404), .B2(new_n406), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n408), .B(new_n399), .C1(new_n401), .C2(new_n411), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT37), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n418), .B(new_n420), .C1(new_n483), .C2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n384), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n479), .B1(new_n407), .B2(new_n412), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT38), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n490), .A2(new_n492), .B1(new_n475), .B2(new_n465), .ZN(new_n493));
  INV_X1    g292(.A(new_n381), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n363), .A2(new_n365), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n340), .A2(new_n346), .A3(new_n285), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n360), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(KEYINPUT39), .C1(new_n360), .C2(new_n359), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(new_n360), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n500), .A2(new_n501), .A3(new_n375), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n500), .B2(new_n375), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n421), .A2(new_n424), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT40), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT86), .B1(new_n493), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n489), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n382), .A2(new_n383), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n492), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(new_n509), .A3(KEYINPUT86), .A4(new_n476), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n478), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n305), .A2(new_n294), .A3(new_n298), .ZN(new_n517));
  INV_X1    g316(.A(new_n303), .ZN(new_n518));
  INV_X1    g317(.A(new_n304), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n294), .A2(new_n298), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n463), .A2(new_n464), .A3(new_n430), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n429), .B1(new_n473), .B2(new_n474), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT35), .B1(new_n524), .B2(new_n425), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT88), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n421), .A2(new_n424), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n476), .A2(new_n527), .A3(new_n384), .A4(new_n521), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT35), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT87), .B1(new_n528), .B2(KEYINPUT35), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n309), .B1(new_n475), .B2(new_n465), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT87), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n426), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n526), .A2(new_n530), .A3(new_n531), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(G1gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT16), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(G1gat), .B2(new_n538), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G8gat), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n541), .B(new_n544), .C1(G1gat), .C2(new_n538), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G43gat), .B(G50gat), .Z(new_n547));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT14), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G43gat), .B(G50gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  NAND2_X1  g356(.A1(G29gat), .A2(G36gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT90), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n549), .A2(new_n555), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(new_n554), .A3(new_n558), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT15), .A3(new_n556), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n546), .B1(new_n563), .B2(KEYINPUT17), .ZN(new_n564));
  AOI211_X1 g363(.A(KEYINPUT91), .B(KEYINPUT17), .C1(new_n560), .C2(new_n562), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n562), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n564), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT92), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n563), .B(new_n546), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n571), .B(KEYINPUT13), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n572), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT91), .B1(new_n563), .B2(KEYINPUT17), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n566), .A3(new_n568), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n581), .B1(new_n584), .B2(new_n564), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n585), .A2(KEYINPUT93), .A3(KEYINPUT18), .A4(new_n571), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n570), .A2(KEYINPUT18), .A3(new_n571), .A4(new_n572), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n573), .A2(KEYINPUT92), .A3(new_n574), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n580), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G113gat), .B(G141gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G169gat), .B(G197gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(KEYINPUT12), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(KEYINPUT12), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n599), .B(new_n598), .C1(new_n576), .C2(new_n578), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n574), .B2(new_n573), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n592), .A2(new_n600), .B1(new_n590), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT95), .B1(new_n612), .B2(new_n607), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(KEYINPUT95), .A3(new_n607), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n610), .B(new_n606), .C1(new_n617), .C2(new_n613), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n618), .A3(KEYINPUT96), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n611), .A2(new_n620), .A3(new_n614), .A4(new_n615), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n567), .ZN(new_n623));
  INV_X1    g422(.A(G232gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n269), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n567), .A2(new_n568), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n569), .A2(new_n565), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT97), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n622), .A2(new_n629), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n584), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n628), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT97), .B1(new_n630), .B2(new_n631), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n584), .A2(new_n633), .A3(new_n634), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n627), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n638), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n638), .A2(new_n643), .A3(KEYINPUT99), .A4(new_n647), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n638), .A2(KEYINPUT98), .A3(new_n643), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n641), .A2(new_n653), .A3(new_n642), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n646), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(G57gat), .A2(G64gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(G57gat), .A2(G64gat), .ZN(new_n658));
  AND2_X1   g457(.A1(G71gat), .A2(G78gat), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n657), .B(new_n658), .C1(new_n659), .C2(KEYINPUT9), .ZN(new_n660));
  AOI22_X1  g459(.A1(KEYINPUT94), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(G71gat), .B2(G78gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(KEYINPUT21), .ZN(new_n664));
  NAND2_X1  g463(.A1(G231gat), .A2(G233gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n204), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n546), .B1(KEYINPUT21), .B2(new_n663), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n666), .B(G127gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n328), .ZN(new_n674));
  XOR2_X1   g473(.A(G183gat), .B(G211gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n669), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n669), .B2(new_n672), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n656), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT10), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n616), .A3(new_n618), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n681), .B(new_n682), .C1(new_n622), .C2(new_n663), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n622), .A2(KEYINPUT10), .A3(new_n663), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n622), .B2(new_n663), .ZN(new_n688));
  INV_X1    g487(.A(new_n686), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(G120gat), .B(G148gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT100), .ZN(new_n692));
  XNOR2_X1  g491(.A(G176gat), .B(G204gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n687), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n689), .B1(new_n683), .B2(new_n684), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(KEYINPUT101), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n698));
  AOI211_X1 g497(.A(new_n698), .B(new_n689), .C1(new_n683), .C2(new_n684), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n690), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n694), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n695), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND4_X1   g501(.A1(new_n537), .A2(new_n604), .A3(new_n680), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n512), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n507), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G8gat), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT16), .B(G8gat), .Z(new_n709));
  NAND3_X1  g508(.A1(new_n703), .A2(new_n507), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n710), .A2(KEYINPUT102), .A3(new_n708), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT102), .B1(new_n710), .B2(new_n708), .ZN(new_n712));
  OAI221_X1 g511(.A(new_n707), .B1(new_n708), .B2(new_n710), .C1(new_n711), .C2(new_n712), .ZN(G1325gat));
  INV_X1    g512(.A(G15gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n703), .A2(new_n714), .A3(new_n521), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n311), .A2(new_n312), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n703), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n717), .B2(new_n714), .ZN(G1326gat));
  INV_X1    g517(.A(new_n476), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT43), .B(G22gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  INV_X1    g521(.A(KEYINPUT86), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n418), .A2(new_n420), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n486), .B(new_n487), .C1(new_n422), .C2(new_n480), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n724), .A2(new_n383), .A3(new_n382), .A4(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n492), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n476), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n477), .B1(new_n730), .B2(new_n514), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n526), .A2(new_n530), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n531), .A2(new_n535), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n656), .ZN(new_n735));
  INV_X1    g534(.A(new_n679), .ZN(new_n736));
  INV_X1    g535(.A(new_n695), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n687), .A2(new_n698), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n696), .A2(KEYINPUT101), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n738), .A2(new_n739), .B1(new_n689), .B2(new_n688), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(new_n694), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n604), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n734), .A2(new_n735), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n550), .A3(new_n512), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT44), .B1(new_n537), .B2(new_n656), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n748), .B(new_n735), .C1(new_n516), .C2(new_n536), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n743), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n384), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n753), .ZN(G1328gat));
  NAND3_X1  g553(.A1(new_n744), .A2(new_n551), .A3(new_n507), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT46), .Z(new_n756));
  OAI21_X1  g555(.A(G36gat), .B1(new_n752), .B2(new_n527), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(G43gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n748), .B1(new_n734), .B2(new_n735), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n537), .A2(KEYINPUT44), .A3(new_n656), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n760), .A2(new_n716), .A3(new_n761), .A4(new_n751), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(KEYINPUT104), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT104), .B2(new_n762), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n744), .A2(new_n759), .A3(new_n521), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(G43gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n765), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT103), .B(KEYINPUT47), .Z(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(G1330gat));
  NOR2_X1   g570(.A1(new_n476), .A2(G50gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n744), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n750), .A2(new_n719), .A3(new_n751), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(G50gat), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n774), .A2(new_n775), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1331gat));
  AND4_X1   g580(.A1(new_n537), .A2(new_n603), .A3(new_n680), .A4(new_n741), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n512), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n507), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT49), .B(G64gat), .Z(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(G1333gat));
  XNOR2_X1  g587(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(G71gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n782), .A2(new_n791), .A3(new_n521), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n782), .B2(new_n716), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n782), .A2(new_n716), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G71gat), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT107), .B1(new_n798), .B2(new_n792), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n790), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n795), .B1(new_n793), .B2(new_n794), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(KEYINPUT107), .A3(new_n792), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n789), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1334gat));
  NAND2_X1  g603(.A1(new_n782), .A2(new_n719), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G78gat), .ZN(G1335gat));
  AND3_X1   g605(.A1(new_n679), .A2(KEYINPUT108), .A3(new_n603), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT108), .B1(new_n679), .B2(new_n603), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n702), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n750), .A2(new_n512), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G85gat), .ZN(new_n812));
  AOI211_X1 g611(.A(new_n735), .B(new_n809), .C1(new_n516), .C2(new_n536), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT51), .ZN(new_n814));
  INV_X1    g613(.A(new_n809), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n537), .A2(new_n656), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n819), .A2(new_n608), .A3(new_n512), .A4(new_n741), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n812), .A2(new_n820), .A3(KEYINPUT109), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1336gat));
  NAND4_X1  g624(.A1(new_n760), .A2(new_n507), .A3(new_n761), .A4(new_n810), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G92gat), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n817), .B1(new_n813), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n741), .A2(new_n609), .A3(new_n507), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT110), .Z(new_n831));
  NAND3_X1  g630(.A1(new_n816), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(new_n819), .B2(new_n831), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n836), .A2(new_n837), .A3(new_n827), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n836), .B2(new_n827), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(G1337gat));
  INV_X1    g639(.A(G99gat), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n819), .A2(new_n841), .A3(new_n521), .A4(new_n741), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n750), .A2(new_n716), .A3(new_n810), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n841), .ZN(G1338gat));
  NOR3_X1   g643(.A1(new_n476), .A2(G106gat), .A3(new_n702), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n819), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n760), .A2(new_n719), .A3(new_n761), .A4(new_n810), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G106gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(KEYINPUT114), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n847), .A2(G106gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n829), .A2(new_n832), .A3(new_n845), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(KEYINPUT53), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n857));
  AOI211_X1 g656(.A(KEYINPUT113), .B(new_n857), .C1(new_n853), .C2(new_n854), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n856), .B2(new_n858), .ZN(G1339gat));
  NAND2_X1  g658(.A1(new_n590), .A2(new_n602), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n576), .A2(new_n578), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n585), .B2(new_n571), .ZN(new_n862));
  INV_X1    g661(.A(new_n597), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT115), .B1(new_n865), .B2(new_n702), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n590), .A2(new_n602), .B1(new_n862), .B2(new_n863), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n741), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n697), .A2(new_n699), .A3(KEYINPUT54), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n683), .A2(new_n689), .A3(new_n684), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n687), .A2(KEYINPUT54), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n701), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n870), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n738), .A2(new_n876), .A3(new_n739), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n877), .A2(KEYINPUT55), .A3(new_n701), .A4(new_n873), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n737), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n866), .B(new_n869), .C1(new_n879), .C2(new_n603), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n735), .ZN(new_n881));
  INV_X1    g680(.A(new_n879), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n656), .A2(new_n882), .A3(new_n868), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n736), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR4_X1   g683(.A1(new_n656), .A2(new_n604), .A3(new_n679), .A4(new_n741), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n524), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n507), .A2(new_n384), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n604), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n741), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g693(.A1(new_n889), .A2(new_n679), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(new_n204), .ZN(G1342gat));
  NOR2_X1   g695(.A1(new_n735), .A2(new_n507), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n898), .B2(new_n384), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n898), .A2(G134gat), .A3(new_n384), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n901), .A2(KEYINPUT116), .A3(new_n900), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT116), .B1(new_n901), .B2(new_n900), .ZN(new_n903));
  OAI221_X1 g702(.A(new_n899), .B1(new_n900), .B2(new_n901), .C1(new_n902), .C2(new_n903), .ZN(G1343gat));
  OAI21_X1  g703(.A(new_n719), .B1(new_n884), .B2(new_n885), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n476), .A2(new_n906), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n879), .A2(new_n603), .B1(new_n702), .B2(new_n865), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n735), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n736), .B1(new_n910), .B2(new_n883), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n911), .B2(new_n885), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT117), .B(new_n908), .C1(new_n911), .C2(new_n885), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n313), .A2(new_n888), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G141gat), .B1(new_n918), .B2(new_n603), .ZN(new_n919));
  INV_X1    g718(.A(new_n905), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n917), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n318), .A3(new_n604), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT58), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT58), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n926), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1344gat));
  OAI21_X1  g727(.A(new_n908), .B1(new_n884), .B2(new_n885), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n885), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n476), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n929), .B1(new_n931), .B2(KEYINPUT57), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n741), .B1(new_n917), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n934), .B1(new_n933), .B2(new_n917), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT59), .B1(new_n936), .B2(new_n319), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n741), .A3(new_n917), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n319), .A2(KEYINPUT59), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(KEYINPUT118), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT118), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n922), .A2(new_n319), .A3(new_n741), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1345gat));
  OAI21_X1  g743(.A(G155gat), .B1(new_n918), .B2(new_n679), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n922), .A2(new_n328), .A3(new_n736), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(KEYINPUT120), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1346gat));
  OAI21_X1  g750(.A(G162gat), .B1(new_n918), .B2(new_n735), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n716), .A2(G162gat), .A3(new_n384), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n920), .A2(new_n897), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n952), .A2(KEYINPUT121), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1347gat));
  NAND2_X1  g758(.A1(new_n507), .A2(new_n384), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n886), .A2(new_n524), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n604), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(G169gat), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT122), .ZN(G1348gat));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n741), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g765(.A1(new_n961), .A2(new_n736), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(new_n219), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n968), .B1(new_n216), .B2(new_n967), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n969), .B(new_n971), .ZN(G1350gat));
  NOR2_X1   g771(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n973), .B1(new_n961), .B2(new_n656), .ZN(new_n974));
  NAND2_X1  g773(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n974), .B(new_n975), .Z(G1351gat));
  NOR2_X1   g775(.A1(new_n716), .A2(new_n960), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n932), .B2(KEYINPUT124), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n980), .B(new_n929), .C1(new_n931), .C2(KEYINPUT57), .ZN(new_n981));
  AND4_X1   g780(.A1(G197gat), .A2(new_n979), .A3(new_n604), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n920), .A2(new_n977), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(G197gat), .B1(new_n984), .B2(new_n604), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n982), .A2(new_n985), .ZN(G1352gat));
  OR2_X1    g785(.A1(new_n911), .A2(new_n885), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT57), .B1(new_n987), .B2(new_n719), .ZN(new_n988));
  INV_X1    g787(.A(new_n929), .ZN(new_n989));
  OAI21_X1  g788(.A(KEYINPUT124), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n990), .A2(new_n741), .A3(new_n977), .A4(new_n981), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n979), .A2(new_n993), .A3(new_n741), .A4(new_n981), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n992), .A2(G204gat), .A3(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(G204gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n984), .A2(new_n996), .A3(new_n741), .ZN(new_n997));
  NAND2_X1  g796(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n998));
  OR2_X1    g797(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n1000), .B1(new_n997), .B2(new_n998), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n995), .A2(new_n1001), .ZN(G1353gat));
  NAND3_X1  g801(.A1(new_n932), .A2(new_n736), .A3(new_n977), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G211gat), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1004), .A2(KEYINPUT63), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(KEYINPUT63), .ZN(new_n1006));
  NOR3_X1   g805(.A1(new_n983), .A2(G211gat), .A3(new_n679), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT127), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(G1354gat));
  AND4_X1   g808(.A1(G218gat), .A2(new_n979), .A3(new_n656), .A4(new_n981), .ZN(new_n1010));
  AOI21_X1  g809(.A(G218gat), .B1(new_n984), .B2(new_n656), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1355gat));
endmodule


