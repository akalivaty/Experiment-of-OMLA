//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G218gat), .ZN(new_n203));
  OR2_X1    g002(.A1(KEYINPUT78), .A2(G211gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT78), .A2(G211gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n206), .B2(KEYINPUT22), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n202), .B(new_n208), .C1(new_n206), .C2(KEYINPUT22), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G226gat), .ZN(new_n213));
  INV_X1    g012(.A(G233gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(KEYINPUT29), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n220), .B(KEYINPUT68), .C1(new_n222), .C2(KEYINPUT26), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n220), .A2(KEYINPUT26), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT27), .B(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(new_n231), .A3(new_n230), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n229), .A2(new_n234), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT25), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n221), .B1(new_n220), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n227), .B2(KEYINPUT23), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n220), .A2(KEYINPUT64), .A3(new_n246), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n238), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n256), .A3(new_n243), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n241), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT66), .A4(new_n243), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n251), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT25), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n263), .A3(KEYINPUT79), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n252), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n261), .B2(new_n251), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n217), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n249), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n222), .B1(KEYINPUT23), .B2(new_n227), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n260), .B2(new_n259), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n238), .B(new_n252), .C1(new_n274), .C2(new_n267), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n275), .A2(new_n213), .A3(new_n214), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n212), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G8gat), .B(G36gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n278), .B(new_n279), .Z(new_n280));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n269), .A3(new_n215), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n216), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n281), .A2(new_n211), .A3(new_n210), .A4(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n277), .A2(new_n283), .ZN(new_n287));
  INV_X1    g086(.A(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n277), .A2(new_n283), .A3(KEYINPUT30), .A4(new_n280), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G141gat), .B(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(G155gat), .B2(G162gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G155gat), .B(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT2), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G134gat), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n311), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(KEYINPUT69), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G120gat), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G113gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n316), .B2(new_n318), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n314), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n316), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT71), .B(G120gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(G113gat), .ZN(new_n327));
  INV_X1    g126(.A(G127gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G134gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n311), .A2(G127gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n321), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n327), .A2(KEYINPUT72), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G120gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n336), .A3(G113gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n316), .ZN(new_n338));
  INV_X1    g137(.A(new_n331), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n333), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n310), .B(new_n324), .C1(new_n332), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n299), .A2(new_n309), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n342), .B1(new_n299), .B2(new_n309), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT72), .B1(new_n327), .B2(new_n331), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n333), .A3(new_n339), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n316), .A2(new_n318), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(new_n321), .A3(new_n320), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n346), .A2(new_n347), .B1(new_n350), .B2(new_n314), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT4), .B(new_n341), .C1(new_n345), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n341), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  OAI21_X1  g163(.A(new_n324), .B1(new_n332), .B2(new_n340), .ZN(new_n365));
  INV_X1    g164(.A(new_n310), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT81), .A3(new_n341), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n368), .A2(new_n358), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n341), .A2(new_n354), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n343), .A2(new_n344), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n346), .A2(new_n347), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n310), .A4(new_n324), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n372), .A2(new_n374), .A3(new_n357), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n360), .B(new_n364), .C1(new_n371), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382));
  INV_X1    g181(.A(new_n364), .ZN(new_n383));
  INV_X1    g182(.A(new_n359), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n352), .B2(new_n355), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n358), .A3(new_n370), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT87), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n360), .B(new_n389), .C1(new_n371), .C2(new_n378), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n382), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n360), .B1(new_n371), .B2(new_n378), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n364), .B1(new_n394), .B2(KEYINPUT87), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT88), .A3(new_n391), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n381), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n383), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT82), .B1(new_n398), .B2(new_n380), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n394), .A2(new_n400), .A3(KEYINPUT6), .A4(new_n383), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n292), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT91), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT91), .B(new_n292), .C1(new_n397), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT73), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n351), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n275), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G227gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(new_n214), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n253), .A2(new_n263), .A3(KEYINPUT73), .A4(new_n365), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT32), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT74), .B(KEYINPUT33), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418));
  XNOR2_X1  g217(.A(G71gat), .B(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n414), .B(KEYINPUT32), .C1(new_n416), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n412), .B1(new_n410), .B2(new_n413), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT75), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT34), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT34), .B1(new_n425), .B2(KEYINPUT75), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n421), .A2(new_n429), .A3(new_n430), .A4(new_n423), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT92), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT31), .B(G50gat), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT29), .B1(new_n210), .B2(new_n211), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n366), .B1(new_n438), .B2(KEYINPUT3), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n343), .A2(KEYINPUT29), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n212), .ZN(new_n443));
  NAND2_X1  g242(.A1(G228gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n440), .A2(new_n441), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n212), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n310), .B1(new_n449), .B2(new_n342), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT84), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n443), .B1(new_n439), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n444), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n437), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n441), .A3(new_n446), .ZN(new_n456));
  INV_X1    g255(.A(new_n437), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n451), .A2(new_n453), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n444), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G22gat), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n455), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n455), .B2(new_n459), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT35), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n432), .A2(KEYINPUT92), .A3(new_n433), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n436), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n405), .A2(new_n406), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n434), .ZN(new_n468));
  INV_X1    g267(.A(new_n463), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n455), .A2(new_n459), .A3(new_n461), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n398), .A2(new_n380), .A3(new_n379), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n399), .A2(new_n474), .A3(new_n401), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n292), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT35), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT37), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n277), .B2(new_n283), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480));
  OR3_X1    g279(.A1(new_n479), .A2(new_n480), .A3(new_n280), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n479), .B2(new_n280), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n277), .A2(new_n478), .A3(new_n283), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT38), .ZN(new_n485));
  INV_X1    g284(.A(new_n381), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n394), .A2(KEYINPUT87), .ZN(new_n487));
  AND4_X1   g286(.A1(KEYINPUT88), .A2(new_n487), .A3(new_n383), .A4(new_n391), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT88), .B1(new_n395), .B2(new_n391), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n402), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n281), .A2(new_n212), .A3(new_n282), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n270), .A2(new_n276), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(KEYINPUT37), .C1(new_n493), .C2(new_n212), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n280), .A2(KEYINPUT38), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n483), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(new_n284), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n485), .A2(new_n490), .A3(new_n491), .A4(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n500), .A2(new_n374), .B1(new_n353), .B2(new_n354), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT85), .B1(new_n501), .B2(new_n358), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n352), .A2(new_n355), .A3(new_n358), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n499), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n368), .A2(new_n370), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT86), .B1(new_n507), .B2(new_n357), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  AOI211_X1 g308(.A(new_n509), .B(new_n358), .C1(new_n368), .C2(new_n370), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(KEYINPUT85), .A3(new_n358), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n503), .A2(new_n504), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT39), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n506), .B(new_n364), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT89), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n506), .A2(new_n364), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n511), .A2(new_n514), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(KEYINPUT40), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n393), .A2(new_n396), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n516), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n291), .A4(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n471), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n498), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n434), .A2(KEYINPUT36), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n529));
  NAND3_X1  g328(.A1(new_n432), .A2(new_n433), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(KEYINPUT77), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n476), .A2(new_n471), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n468), .A2(new_n533), .A3(new_n529), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n467), .A2(new_n477), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(G1gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(G1gat), .B2(new_n538), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n545));
  AOI21_X1  g344(.A(G36gat), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G29gat), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n547), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n548));
  OR3_X1    g347(.A1(new_n546), .A2(KEYINPUT15), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT15), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n543), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n541), .B(G8gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n553), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n537), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n552), .A3(new_n553), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n560), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n562), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n557), .A2(KEYINPUT18), .A3(new_n562), .A4(new_n560), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT11), .B(G169gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n564), .A2(new_n568), .A3(new_n575), .A4(new_n569), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G99gat), .B(G106gat), .ZN(new_n581));
  AND2_X1   g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(KEYINPUT96), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT96), .B1(new_n585), .B2(new_n583), .ZN(new_n586));
  MUX2_X1   g385(.A(new_n582), .B(new_n584), .S(new_n586), .Z(new_n587));
  INV_X1    g386(.A(KEYINPUT8), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(KEYINPUT97), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(KEYINPUT97), .B2(new_n589), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT98), .B(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n591), .B2(new_n594), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n581), .B(new_n587), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n591), .A2(new_n594), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT99), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n581), .B1(new_n603), .B2(new_n587), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n606));
  AOI211_X1 g405(.A(KEYINPUT100), .B(new_n581), .C1(new_n603), .C2(new_n587), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n599), .A2(new_n604), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n587), .B1(new_n596), .B2(new_n597), .ZN(new_n610));
  INV_X1    g409(.A(new_n581), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(KEYINPUT100), .A3(new_n598), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT101), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  OAI22_X1  g413(.A1(new_n608), .A2(new_n614), .B1(new_n556), .B2(new_n555), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n606), .B1(new_n605), .B2(new_n607), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n609), .A2(new_n613), .A3(KEYINPUT101), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n559), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n621), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n615), .A2(new_n618), .A3(new_n626), .A4(new_n619), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n622), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n622), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G183gat), .B(G211gat), .Z(new_n631));
  XNOR2_X1  g430(.A(G57gat), .B(G64gat), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G71gat), .B(G78gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n642), .B2(new_n645), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n631), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  INV_X1    g449(.A(new_n631), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n646), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n543), .B1(new_n637), .B2(new_n636), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n649), .A2(new_n652), .ZN(new_n657));
  INV_X1    g456(.A(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n630), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n636), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n598), .B1(new_n612), .B2(KEYINPUT102), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n604), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n661), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n636), .B1(new_n605), .B2(new_n607), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT104), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  INV_X1    g474(.A(new_n598), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n604), .B2(new_n663), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n612), .A2(KEYINPUT102), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n636), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n661), .B1(new_n609), .B2(new_n613), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n666), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(KEYINPUT103), .A3(new_n675), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n608), .A2(new_n614), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n636), .A2(new_n675), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n683), .A2(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n669), .B(new_n674), .C1(new_n688), .C2(new_n668), .ZN(new_n689));
  INV_X1    g488(.A(new_n669), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT103), .B1(new_n684), .B2(new_n675), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n682), .B(KEYINPUT10), .C1(new_n665), .C2(new_n666), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n667), .B(KEYINPUT105), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n690), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n689), .B1(new_n697), .B2(new_n674), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n660), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n536), .A2(new_n580), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n475), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n291), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT106), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT16), .B(G8gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(G8gat), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n706), .A2(new_n705), .A3(new_n708), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(G1325gat));
  INV_X1    g511(.A(new_n436), .ZN(new_n713));
  INV_X1    g512(.A(new_n465), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(G15gat), .B1(new_n701), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT107), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n531), .A2(new_n534), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n701), .A2(G15gat), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n717), .A2(new_n719), .ZN(G1326gat));
  NAND2_X1  g519(.A1(new_n701), .A2(new_n471), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT43), .B(G22gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1327gat));
  NAND2_X1  g522(.A1(new_n659), .A2(new_n656), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n579), .A3(new_n699), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT35), .ZN(new_n728));
  INV_X1    g527(.A(new_n476), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n472), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n436), .A2(new_n464), .A3(new_n465), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n403), .B2(new_n404), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n732), .B2(new_n406), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n524), .A2(new_n291), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n488), .A2(new_n489), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n471), .B1(new_n737), .B2(new_n522), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n734), .B1(new_n738), .B2(new_n498), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n630), .B(new_n727), .C1(new_n733), .C2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n740), .A2(G29gat), .A3(new_n475), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT45), .Z(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  INV_X1    g542(.A(new_n630), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n536), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(KEYINPUT44), .B(new_n630), .C1(new_n733), .C2(new_n739), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n727), .ZN(new_n748));
  OAI21_X1  g547(.A(G29gat), .B1(new_n748), .B2(new_n475), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n742), .A2(new_n749), .ZN(G1328gat));
  OAI21_X1  g549(.A(G36gat), .B1(new_n748), .B2(new_n292), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n740), .A2(G36gat), .A3(new_n292), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT46), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1329gat));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755));
  INV_X1    g554(.A(new_n715), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n740), .A2(G43gat), .A3(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT109), .Z(new_n758));
  INV_X1    g557(.A(new_n718), .ZN(new_n759));
  OAI21_X1  g558(.A(G43gat), .B1(new_n748), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n755), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT47), .Z(G1330gat));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n471), .A3(new_n746), .A4(new_n727), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G50gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n291), .B1(new_n490), .B2(new_n491), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n466), .B1(new_n765), .B2(KEYINPUT91), .ZN(new_n766));
  INV_X1    g565(.A(new_n406), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n477), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n527), .A2(new_n535), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n744), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT110), .B1(new_n770), .B2(new_n727), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n526), .A2(G50gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n740), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n764), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT48), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n774), .B2(new_n771), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n770), .A2(KEYINPUT110), .A3(new_n727), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n740), .A2(new_n773), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT111), .A4(new_n772), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n776), .B1(new_n763), .B2(G50gat), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT112), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND4_X1   g584(.A1(KEYINPUT112), .A2(new_n784), .A3(new_n782), .A4(new_n779), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT113), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n777), .C1(new_n785), .C2(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1331gat));
  INV_X1    g590(.A(new_n536), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n580), .A3(new_n660), .A4(new_n698), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n475), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g594(.A(new_n793), .B(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n291), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT49), .B(G64gat), .Z(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(G1333gat));
  NAND3_X1  g599(.A1(new_n796), .A2(G71gat), .A3(new_n718), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n793), .A2(new_n756), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(G71gat), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g603(.A1(new_n796), .A2(new_n471), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g605(.A1(new_n725), .A2(new_n580), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n536), .A2(new_n744), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n699), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n702), .A3(new_n592), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n807), .A2(new_n699), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n747), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n475), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n815), .B2(new_n592), .ZN(G1336gat));
  OAI21_X1  g615(.A(G92gat), .B1(new_n814), .B2(new_n292), .ZN(new_n817));
  INV_X1    g616(.A(new_n811), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n291), .A2(new_n593), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g620(.A(KEYINPUT115), .B1(new_n814), .B2(new_n759), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G99gat), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n814), .A2(KEYINPUT115), .A3(new_n759), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n756), .A2(G99gat), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n823), .A2(new_n824), .B1(new_n818), .B2(new_n825), .ZN(G1338gat));
  NAND3_X1  g625(.A1(new_n747), .A2(new_n471), .A3(new_n813), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G106gat), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT53), .B1(new_n828), .B2(KEYINPUT116), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n526), .A2(G106gat), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n811), .A2(new_n830), .B1(new_n827), .B2(G106gat), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n829), .B(new_n831), .ZN(G1339gat));
  NAND3_X1  g631(.A1(new_n660), .A2(new_n580), .A3(new_n699), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n695), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n837), .B(KEYINPUT54), .C1(new_n688), .C2(new_n668), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n694), .A2(new_n839), .A3(new_n696), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n673), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n841), .A2(KEYINPUT118), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT118), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n574), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n566), .A2(new_n567), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n561), .A2(new_n563), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n562), .B1(new_n557), .B2(new_n560), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n846), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n578), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT120), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n852), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n851), .A2(KEYINPUT119), .B1(new_n566), .B2(new_n567), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n574), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n578), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n628), .A3(new_n629), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n673), .A4(new_n840), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n689), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n836), .B1(new_n845), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n862), .A2(new_n863), .A3(new_n689), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n866), .B(KEYINPUT121), .C1(new_n844), .C2(new_n843), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n842), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n841), .A2(KEYINPUT118), .A3(new_n842), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n863), .A2(new_n579), .A3(new_n689), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n578), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n872), .A2(new_n874), .B1(new_n698), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n865), .B(new_n867), .C1(new_n877), .C2(new_n630), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n835), .B1(new_n878), .B2(new_n725), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n475), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n473), .A2(new_n291), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n579), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n867), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n872), .A2(new_n874), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n698), .A2(new_n876), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n630), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n725), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n835), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n756), .A2(new_n471), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n475), .A2(new_n291), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n580), .A2(new_n315), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n883), .B1(new_n895), .B2(new_n896), .ZN(G1340gat));
  NOR3_X1   g696(.A1(new_n879), .A2(new_n471), .A3(new_n756), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n893), .ZN(new_n899));
  OAI21_X1  g698(.A(G120gat), .B1(new_n899), .B2(new_n699), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n326), .A3(new_n698), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1341gat));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n328), .B1(new_n895), .B2(new_n724), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n725), .A2(G127gat), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n880), .A2(new_n881), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G127gat), .B1(new_n899), .B2(new_n725), .ZN(new_n908));
  INV_X1    g707(.A(new_n906), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(KEYINPUT122), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(G1342gat));
  NAND3_X1  g710(.A1(new_n882), .A2(new_n311), .A3(new_n630), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT56), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n882), .A2(new_n914), .A3(new_n311), .A4(new_n630), .ZN(new_n915));
  OAI21_X1  g714(.A(G134gat), .B1(new_n899), .B2(new_n744), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(G1343gat));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  INV_X1    g717(.A(new_n867), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT121), .B1(new_n872), .B2(new_n866), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n886), .B1(new_n845), .B2(new_n873), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n744), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n724), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n918), .B(new_n471), .C1(new_n924), .C2(new_n835), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n718), .A2(new_n894), .ZN(new_n926));
  INV_X1    g725(.A(new_n868), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n886), .B1(new_n927), .B2(new_n873), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n744), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n865), .A2(new_n867), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n835), .B1(new_n930), .B2(new_n725), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT57), .B1(new_n931), .B2(new_n526), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n925), .A2(new_n579), .A3(new_n926), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G141gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n718), .A2(new_n526), .A3(new_n291), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n880), .A2(new_n300), .A3(new_n579), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT58), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT58), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1344gat));
  NOR2_X1   g740(.A1(new_n699), .A2(G148gat), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n890), .A2(new_n702), .A3(new_n935), .A4(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT57), .B1(new_n879), .B2(new_n526), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n872), .A2(new_n866), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n724), .B1(new_n929), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n833), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n918), .B(new_n471), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n947), .A2(new_n698), .A3(new_n926), .A4(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(new_n302), .ZN(new_n954));
  AOI22_X1  g753(.A1(new_n945), .A2(new_n946), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n925), .A2(new_n926), .A3(new_n932), .ZN(new_n956));
  OAI21_X1  g755(.A(G148gat), .B1(new_n956), .B2(new_n699), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n953), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n958), .ZN(G1345gat));
  OAI21_X1  g758(.A(G155gat), .B1(new_n956), .B2(new_n725), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n880), .A2(new_n306), .A3(new_n724), .A4(new_n935), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1346gat));
  NAND4_X1  g761(.A1(new_n890), .A2(new_n702), .A3(new_n630), .A4(new_n935), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n307), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n630), .A2(G162gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT124), .ZN(G1347gat));
  NOR2_X1   g766(.A1(new_n473), .A2(new_n292), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n879), .A2(new_n702), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G169gat), .B1(new_n970), .B2(new_n579), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n702), .A2(new_n292), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n892), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n580), .A2(new_n218), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1348gat));
  NAND3_X1  g775(.A1(new_n970), .A2(new_n219), .A3(new_n698), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n892), .A2(new_n699), .A3(new_n973), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n219), .ZN(G1349gat));
  NAND4_X1  g778(.A1(new_n890), .A2(new_n724), .A3(new_n891), .A4(new_n972), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G183gat), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n724), .A2(new_n230), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n970), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n702), .B1(new_n888), .B2(new_n889), .ZN(new_n985));
  AND4_X1   g784(.A1(new_n982), .A2(new_n985), .A3(new_n968), .A4(new_n983), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT60), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT60), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n989), .B(new_n981), .C1(new_n984), .C2(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1350gat));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n231), .A3(new_n630), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n898), .A2(new_n630), .A3(new_n972), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n995));
  AND4_X1   g794(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(G190gat), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n231), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n997));
  AOI22_X1  g796(.A1(new_n994), .A2(new_n997), .B1(new_n993), .B2(new_n995), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n992), .B1(new_n996), .B2(new_n998), .ZN(G1351gat));
  NOR2_X1   g798(.A1(new_n718), .A2(new_n973), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n947), .A2(new_n951), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(G197gat), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n1001), .A2(new_n1002), .A3(new_n580), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n759), .A2(new_n471), .A3(new_n291), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT127), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n985), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g806(.A(G197gat), .B1(new_n1007), .B2(new_n579), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n1003), .A2(new_n1008), .ZN(G1352gat));
  NOR3_X1   g808(.A1(new_n1006), .A2(G204gat), .A3(new_n699), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT62), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g811(.A(G204gat), .B1(new_n1001), .B2(new_n699), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(G1353gat));
  NAND4_X1  g814(.A1(new_n1007), .A2(new_n204), .A3(new_n205), .A4(new_n724), .ZN(new_n1016));
  NAND4_X1  g815(.A1(new_n947), .A2(new_n724), .A3(new_n951), .A4(new_n1000), .ZN(new_n1017));
  AND3_X1   g816(.A1(new_n1017), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1018));
  AOI21_X1  g817(.A(KEYINPUT63), .B1(new_n1017), .B2(G211gat), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(G1354gat));
  OAI21_X1  g819(.A(G218gat), .B1(new_n1001), .B2(new_n744), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1007), .A2(new_n203), .A3(new_n630), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1021), .A2(new_n1022), .ZN(G1355gat));
endmodule


