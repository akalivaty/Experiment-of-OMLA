//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n203), .A2(new_n206), .A3(new_n207), .A4(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n204), .B(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(new_n208), .ZN(new_n213));
  OAI211_X1 g012(.A(KEYINPUT15), .B(new_n202), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT17), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G1gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  INV_X1    g023(.A(G15gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(G22gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G15gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n222), .A2(new_n223), .A3(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n230), .B(G8gat), .C1(new_n223), .C2(new_n222), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(KEYINPUT88), .ZN(new_n232));
  INV_X1    g031(.A(G8gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT88), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n220), .B(new_n234), .C1(new_n221), .C2(G1gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n229), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n215), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n241), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n240), .B(KEYINPUT13), .Z(new_n246));
  INV_X1    g045(.A(new_n241), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n237), .A2(new_n215), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G169gat), .B(G197gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT12), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n244), .A2(new_n245), .A3(new_n249), .A4(new_n256), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(G169gat), .B2(G176gat), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(G169gat), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT23), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT24), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n264), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT66), .B(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(new_n273), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n283), .A2(KEYINPUT25), .A3(new_n269), .A4(new_n264), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT26), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n287), .A2(new_n270), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G183gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n293), .A3(KEYINPUT27), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295));
  AOI21_X1  g094(.A(G190gat), .B1(new_n295), .B2(G183gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT28), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n280), .B1(new_n290), .B2(KEYINPUT27), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n295), .A2(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n289), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G226gat), .ZN(new_n303));
  INV_X1    g102(.A(G233gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT22), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n307), .A3(new_n311), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT73), .B1(new_n315), .B2(new_n316), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g122(.A(KEYINPUT67), .B(new_n289), .C1(new_n297), .C2(new_n301), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(new_n278), .B2(new_n284), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n305), .A2(KEYINPUT29), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n306), .B(new_n321), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n285), .A2(new_n302), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n325), .A2(new_n305), .B1(new_n329), .B2(new_n326), .ZN(new_n330));
  INV_X1    g129(.A(new_n317), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n328), .B(new_n335), .C1(new_n330), .C2(new_n331), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n338), .ZN(new_n339));
  OR3_X1    g138(.A1(new_n332), .A2(KEYINPUT30), .A3(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(G1gat), .B(G29gat), .Z(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT69), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G127gat), .B(G134gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT69), .ZN(new_n352));
  INV_X1    g151(.A(G120gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(G113gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(G127gat), .A2(G134gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT68), .B(G127gat), .ZN(new_n358));
  INV_X1    g157(.A(G134gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n347), .A2(KEYINPUT1), .ZN(new_n361));
  OAI22_X1  g160(.A1(new_n349), .A2(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(G155gat), .B2(G162gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G141gat), .B(G148gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(G155gat), .B2(G162gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G155gat), .B(G162gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n374));
  INV_X1    g173(.A(G141gat), .ZN(new_n375));
  INV_X1    g174(.A(G148gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n370), .A3(new_n365), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n379), .A2(new_n370), .A3(new_n365), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n370), .B1(new_n379), .B2(new_n365), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(KEYINPUT3), .A3(new_n380), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n362), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n384), .A2(new_n385), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n362), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n382), .A2(new_n388), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n355), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n348), .ZN(new_n399));
  INV_X1    g198(.A(new_n360), .ZN(new_n400));
  INV_X1    g199(.A(new_n361), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(new_n362), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n392), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n394), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n393), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n346), .B1(new_n397), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n382), .A2(new_n388), .A3(new_n391), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n406), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n411), .B(KEYINPUT39), .C1(new_n406), .C2(new_n405), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT39), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n413), .A3(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n414), .A2(new_n415), .A3(new_n346), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n414), .B2(new_n346), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT40), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n409), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT40), .B(new_n412), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n421), .A2(KEYINPUT82), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(KEYINPUT82), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n342), .B(new_n420), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(G50gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT77), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n427), .B(KEYINPUT31), .Z(new_n428));
  INV_X1    g227(.A(G228gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n304), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n315), .B2(new_n316), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n390), .B1(new_n432), .B2(KEYINPUT3), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n317), .B1(new_n386), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT78), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT3), .B1(new_n372), .B2(new_n380), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n331), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT78), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n431), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n316), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n313), .B1(new_n311), .B2(new_n307), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n434), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n381), .B1(new_n444), .B2(new_n383), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT79), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n433), .A2(new_n447), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n319), .A2(new_n320), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .A4(new_n430), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n227), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n428), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n445), .B1(new_n439), .B2(KEYINPUT78), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n436), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n430), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n450), .ZN(new_n457));
  OAI21_X1  g256(.A(G22gat), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n227), .A3(new_n450), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n458), .A2(new_n459), .A3(new_n452), .A4(new_n428), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n346), .ZN(new_n464));
  INV_X1    g263(.A(new_n408), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(new_n396), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n397), .A2(new_n408), .A3(new_n346), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n409), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n332), .A2(KEYINPUT37), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n336), .B1(new_n332), .B2(KEYINPUT37), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT38), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n466), .A2(new_n469), .A3(new_n467), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT83), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n306), .ZN(new_n481));
  INV_X1    g280(.A(new_n299), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT28), .A3(new_n296), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n298), .B1(new_n279), .B2(KEYINPUT27), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(KEYINPUT28), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT67), .B1(new_n485), .B2(new_n289), .ZN(new_n486));
  INV_X1    g285(.A(new_n324), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n285), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n488), .B2(new_n326), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n329), .A2(new_n326), .ZN(new_n490));
  INV_X1    g289(.A(new_n305), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n489), .A2(new_n321), .B1(new_n492), .B2(new_n317), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT38), .B1(new_n493), .B2(KEYINPUT37), .ZN(new_n494));
  INV_X1    g293(.A(new_n475), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n338), .C1(new_n476), .C2(KEYINPUT84), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n424), .B(new_n463), .C1(new_n480), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n488), .A2(new_n363), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n323), .A2(new_n324), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n362), .A3(new_n285), .ZN(new_n501));
  NAND2_X1  g300(.A1(G227gat), .A2(G233gat), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n502), .B(KEYINPUT64), .Z(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT32), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT33), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G71gat), .B(G99gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT70), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(new_n225), .ZN(new_n510));
  INV_X1    g309(.A(G43gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT32), .B(new_n504), .C1(new_n514), .C2(new_n506), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n503), .A2(KEYINPUT34), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n500), .A2(new_n362), .A3(new_n285), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n362), .B1(new_n500), .B2(new_n285), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n502), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n499), .B2(new_n501), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT34), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT71), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n520), .B(new_n526), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n515), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(new_n527), .A3(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT72), .B1(new_n516), .B2(new_n528), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n530), .A2(new_n536), .A3(new_n527), .A4(new_n525), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n535), .A2(KEYINPUT36), .A3(new_n529), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n463), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n478), .A2(new_n472), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n341), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n498), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n535), .A2(new_n529), .A3(new_n537), .A4(new_n463), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT35), .B1(new_n545), .B2(new_n542), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n531), .A2(new_n547), .A3(new_n341), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n473), .A2(new_n479), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n548), .A2(new_n529), .A3(new_n549), .A4(new_n463), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n261), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(G64gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G57gat), .ZN(new_n555));
  INV_X1    g354(.A(G57gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G64gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  OR2_X1    g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT89), .B1(new_n556), .B2(G64gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n554), .A3(G57gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n565), .A3(new_n557), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n563), .A2(new_n565), .A3(new_n568), .A4(new_n557), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n560), .B1(new_n561), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n562), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n575));
  NAND2_X1  g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(G99gat), .ZN(new_n578));
  INV_X1    g377(.A(G106gat), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT8), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(G85gat), .B(G92gat), .C1(KEYINPUT91), .C2(KEYINPUT7), .ZN(new_n582));
  AND2_X1   g381(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT96), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n573), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(new_n581), .B2(new_n584), .ZN(new_n589));
  INV_X1    g388(.A(new_n584), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n590), .A2(new_n587), .A3(new_n577), .A4(new_n580), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n589), .A2(new_n591), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n594), .A3(new_n585), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT10), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT92), .B1(new_n589), .B2(new_n591), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n589), .A2(new_n591), .A3(KEYINPUT92), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n570), .A2(new_n572), .ZN(new_n602));
  INV_X1    g401(.A(new_n562), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n553), .B1(new_n596), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n553), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n593), .A2(new_n607), .A3(new_n595), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n606), .A2(new_n608), .A3(new_n612), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n598), .A2(new_n215), .A3(new_n599), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n218), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n217), .B1(new_n211), .B2(new_n214), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n599), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n597), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT93), .B1(new_n219), .B2(new_n600), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n630), .B1(new_n627), .B2(new_n629), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n219), .A2(new_n600), .A3(KEYINPUT93), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n624), .A3(new_n636), .ZN(new_n642));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n638), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n636), .B1(new_n641), .B2(new_n624), .ZN(new_n648));
  AOI211_X1 g447(.A(new_n637), .B(new_n623), .C1(new_n639), .C2(new_n640), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(G231gat), .B(G233gat), .C1(new_n573), .C2(KEYINPUT21), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT21), .ZN(new_n652));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n604), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(G127gat), .ZN(new_n656));
  INV_X1    g455(.A(G127gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n651), .A2(new_n657), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n237), .B1(KEYINPUT21), .B2(new_n573), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n662), .A3(new_n658), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n664));
  INV_X1    g463(.A(G155gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(G183gat), .B(G211gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n661), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n661), .B2(new_n663), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n646), .B(new_n650), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n619), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n552), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n541), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n224), .ZN(G1324gat));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n341), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT99), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n681), .B(new_n683), .C1(new_n233), .C2(new_n676), .ZN(G1325gat));
  INV_X1    g483(.A(new_n673), .ZN(new_n685));
  INV_X1    g484(.A(new_n532), .ZN(new_n686));
  AOI21_X1  g485(.A(G15gat), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n539), .A2(new_n225), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT100), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n685), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n673), .A2(new_n463), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n498), .A2(new_n539), .A3(new_n543), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n551), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n546), .A2(KEYINPUT101), .A3(new_n550), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n648), .A2(new_n649), .A3(new_n647), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n645), .B1(new_n638), .B2(new_n642), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n694), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  AOI211_X1 g502(.A(new_n694), .B(new_n702), .C1(new_n544), .C2(new_n551), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n619), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n669), .A2(new_n670), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n260), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n711), .B2(new_n541), .ZN(new_n712));
  INV_X1    g511(.A(new_n702), .ZN(new_n713));
  AND4_X1   g512(.A1(new_n552), .A2(new_n708), .A3(new_n713), .A4(new_n707), .ZN(new_n714));
  INV_X1    g513(.A(G29gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n541), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n712), .A2(new_n718), .ZN(G1328gat));
  OAI21_X1  g518(.A(G36gat), .B1(new_n711), .B2(new_n341), .ZN(new_n720));
  INV_X1    g519(.A(G36gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n714), .A2(new_n721), .A3(new_n342), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT46), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(G1329gat));
  AOI21_X1  g523(.A(G43gat), .B1(new_n714), .B2(new_n686), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n539), .A2(new_n511), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n710), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g527(.A(G50gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n710), .B2(new_n540), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n729), .A3(new_n540), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT103), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT102), .B(KEYINPUT48), .Z(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(KEYINPUT48), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n733), .A2(new_n734), .B1(new_n730), .B2(new_n735), .ZN(G1331gat));
  AND3_X1   g535(.A1(new_n546), .A2(KEYINPUT101), .A3(new_n550), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT101), .B1(new_n546), .B2(new_n550), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n544), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n707), .A2(new_n260), .A3(new_n671), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n541), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(new_n556), .ZN(G1332gat));
  XNOR2_X1  g542(.A(new_n741), .B(KEYINPUT104), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n341), .B(KEYINPUT105), .Z(new_n745));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n554), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n554), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1333gat));
  NAND4_X1  g548(.A1(new_n744), .A2(G71gat), .A3(new_n534), .A4(new_n538), .ZN(new_n750));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n741), .B2(new_n532), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n540), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  INV_X1    g555(.A(new_n708), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n260), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n739), .A2(new_n713), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT106), .B(KEYINPUT51), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n739), .A2(new_n713), .A3(new_n758), .A4(new_n763), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n762), .A2(new_n619), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(G85gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(new_n716), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n739), .A2(new_n713), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n704), .B1(new_n768), .B2(new_n694), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n758), .A2(new_n619), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n541), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n767), .A2(new_n773), .ZN(G1336gat));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  INV_X1    g574(.A(new_n745), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n762), .A2(new_n619), .A3(new_n764), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n703), .A2(new_n705), .A3(new_n745), .A4(new_n771), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n775), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AND4_X1   g582(.A1(new_n775), .A2(new_n782), .A3(new_n779), .A4(new_n778), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n703), .A2(new_n342), .A3(new_n705), .A4(new_n771), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n778), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT107), .B1(new_n787), .B2(KEYINPUT52), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n789), .B(new_n779), .C1(new_n786), .C2(new_n778), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n783), .A2(new_n784), .B1(new_n788), .B2(new_n790), .ZN(G1337gat));
  NAND3_X1  g590(.A1(new_n765), .A2(new_n578), .A3(new_n686), .ZN(new_n792));
  OAI21_X1  g591(.A(G99gat), .B1(new_n772), .B2(new_n539), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n769), .A2(new_n540), .A3(new_n771), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT109), .B(G106gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(KEYINPUT53), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n765), .A2(new_n579), .A3(new_n540), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n798), .B2(new_n799), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n619), .A2(new_n671), .A3(new_n260), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n573), .A2(new_n594), .A3(new_n585), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n594), .B1(new_n573), .B2(new_n585), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n601), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n629), .A2(KEYINPUT10), .A3(new_n573), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n607), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n612), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n607), .A3(new_n809), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n606), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT55), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n247), .A2(new_n248), .A3(new_n246), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n255), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n259), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n700), .B2(new_n701), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n615), .B(new_n616), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n650), .A2(new_n646), .A3(new_n258), .A4(new_n259), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n819), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n619), .A2(new_n259), .A3(new_n702), .A4(new_n822), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n805), .B1(new_n829), .B2(new_n708), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n804), .B1(new_n830), .B2(new_n540), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n757), .B1(new_n827), .B2(new_n828), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT111), .B(new_n463), .C1(new_n832), .C2(new_n805), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n745), .A2(new_n541), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n834), .A2(new_n686), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(G113gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n261), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n830), .A2(new_n541), .ZN(new_n839));
  INV_X1    g638(.A(new_n545), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n776), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(new_n261), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n836), .A2(new_n838), .B1(new_n842), .B2(new_n837), .ZN(G1340gat));
  NOR2_X1   g642(.A1(new_n707), .A2(new_n353), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n841), .A2(new_n707), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n836), .A2(new_n844), .B1(new_n845), .B2(new_n353), .ZN(G1341gat));
  INV_X1    g645(.A(new_n358), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n841), .A2(new_n847), .A3(new_n708), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n836), .A2(new_n757), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n847), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT112), .Z(G1342gat));
  NAND2_X1  g650(.A1(new_n839), .A2(new_n840), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n713), .A2(new_n341), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n852), .A2(G134gat), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT56), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n836), .A2(new_n713), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n359), .B2(new_n856), .ZN(G1343gat));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n830), .B2(new_n463), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n540), .C1(new_n832), .C2(new_n805), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n835), .A2(new_n539), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G141gat), .B1(new_n864), .B2(new_n261), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n463), .B1(new_n534), .B2(new_n538), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n839), .A2(new_n776), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n375), .A3(new_n260), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n862), .B1(new_n859), .B2(new_n860), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(KEYINPUT113), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n874), .B(new_n862), .C1(new_n859), .C2(new_n860), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n873), .A2(new_n875), .A3(new_n261), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT114), .B1(new_n876), .B2(new_n375), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n864), .A2(new_n874), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n872), .A2(KEYINPUT113), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n878), .B(G141gat), .C1(new_n881), .C2(new_n261), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n877), .A2(new_n882), .A3(new_n870), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n871), .B1(new_n883), .B2(new_n866), .ZN(G1344gat));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n707), .B1(new_n862), .B2(KEYINPUT115), .ZN(new_n886));
  INV_X1    g685(.A(new_n860), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n859), .B1(new_n887), .B2(KEYINPUT116), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n860), .A2(new_n889), .ZN(new_n890));
  OAI221_X1 g689(.A(new_n886), .B1(KEYINPUT115), .B2(new_n862), .C1(new_n888), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G148gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n879), .A2(new_n619), .A3(new_n880), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n376), .A2(KEYINPUT59), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n892), .A2(KEYINPUT59), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n868), .A2(G148gat), .A3(new_n707), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n885), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n896), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n893), .A2(new_n894), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n891), .B2(G148gat), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT117), .B(new_n898), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(G155gat), .B1(new_n881), .B2(new_n708), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n869), .A2(new_n665), .A3(new_n757), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n881), .B2(new_n702), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n853), .A2(G162gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n839), .A2(new_n867), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1347gat));
  AND2_X1   g709(.A1(new_n831), .A2(new_n833), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n716), .A2(new_n341), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n686), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT119), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n831), .B2(new_n833), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(new_n265), .A3(new_n261), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n830), .A2(new_n716), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n840), .A3(new_n745), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n260), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n921), .A2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n920), .B2(new_n707), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n266), .A3(new_n619), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  NAND2_X1  g728(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n295), .A2(G183gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n757), .A2(new_n931), .A3(new_n482), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n757), .A3(new_n919), .ZN(new_n934));
  INV_X1    g733(.A(new_n279), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n924), .A2(new_n280), .A3(new_n713), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n917), .A2(new_n918), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT119), .B(new_n915), .C1(new_n831), .C2(new_n833), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n940), .A2(new_n941), .A3(new_n702), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT121), .B1(new_n942), .B2(new_n280), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n916), .A2(new_n713), .A3(new_n919), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n946), .A3(G190gat), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n943), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n939), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  OR2_X1    g749(.A1(new_n888), .A2(new_n890), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n539), .A2(new_n912), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(G197gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n953), .A2(new_n954), .A3(new_n261), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n867), .A2(new_n745), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n922), .B1(KEYINPUT122), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(KEYINPUT122), .B2(new_n956), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n260), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n955), .A2(new_n959), .ZN(G1352gat));
  XNOR2_X1  g759(.A(KEYINPUT123), .B(G204gat), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n707), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n953), .B2(new_n707), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT124), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(G1353gat));
  NAND3_X1  g768(.A1(new_n958), .A2(new_n309), .A3(new_n757), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n757), .A3(new_n952), .ZN(new_n972));
  AND4_X1   g771(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(G211gat), .B1(new_n971), .B2(KEYINPUT63), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI22_X1  g774(.A1(new_n972), .A2(new_n975), .B1(new_n971), .B2(KEYINPUT63), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n970), .B1(new_n973), .B2(new_n976), .ZN(G1354gat));
  AND2_X1   g776(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n713), .B1(new_n953), .B2(KEYINPUT127), .ZN(new_n979));
  OAI21_X1  g778(.A(G218gat), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n958), .A2(new_n310), .A3(new_n713), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1355gat));
endmodule


