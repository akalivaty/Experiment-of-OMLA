

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U555 ( .A(KEYINPUT94), .B(n755), .ZN(n711) );
  NOR2_X1 U556 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U557 ( .A1(n789), .A2(n775), .ZN(n776) );
  XOR2_X1 U558 ( .A(n744), .B(KEYINPUT29), .Z(n522) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(n715), .ZN(n719) );
  NOR2_X1 U560 ( .A1(n719), .A2(n718), .ZN(n722) );
  INV_X1 U561 ( .A(G2105), .ZN(n527) );
  NOR2_X1 U562 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U563 ( .A(KEYINPUT1), .B(n539), .Z(n652) );
  AND2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n855) );
  NAND2_X1 U565 ( .A1(n855), .A2(G113), .ZN(n525) );
  AND2_X4 U566 ( .A1(n527), .A2(G2104), .ZN(n858) );
  NAND2_X1 U567 ( .A1(G101), .A2(n858), .ZN(n523) );
  XOR2_X1 U568 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  NAND2_X1 U569 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U571 ( .A(KEYINPUT17), .B(n526), .Z(n859) );
  NAND2_X1 U572 ( .A1(G137), .A2(n859), .ZN(n529) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n527), .ZN(n854) );
  NAND2_X1 U574 ( .A1(G125), .A2(n854), .ZN(n528) );
  NAND2_X1 U575 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U576 ( .A1(n531), .A2(n530), .ZN(G160) );
  XNOR2_X1 U577 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U578 ( .A(G82), .ZN(G220) );
  INV_X1 U579 ( .A(G132), .ZN(G219) );
  XNOR2_X1 U580 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  NOR2_X1 U581 ( .A1(G220), .A2(G219), .ZN(n532) );
  XOR2_X1 U582 ( .A(KEYINPUT22), .B(n532), .Z(n533) );
  NOR2_X1 U583 ( .A1(G218), .A2(n533), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G96), .A2(n534), .ZN(n820) );
  NAND2_X1 U585 ( .A1(n820), .A2(G2106), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G108), .A2(G120), .ZN(n535) );
  NOR2_X1 U587 ( .A1(G237), .A2(n535), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G69), .A2(n536), .ZN(n821) );
  NAND2_X1 U589 ( .A1(n821), .A2(G567), .ZN(n537) );
  AND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(G319) );
  INV_X1 U591 ( .A(G651), .ZN(n543) );
  NOR2_X1 U592 ( .A1(G543), .A2(n543), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n652), .A2(G64), .ZN(n542) );
  XOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  NOR2_X1 U595 ( .A1(G651), .A2(n632), .ZN(n540) );
  XNOR2_X1 U596 ( .A(KEYINPUT64), .B(n540), .ZN(n645) );
  NAND2_X1 U597 ( .A1(G52), .A2(n645), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n548) );
  NOR2_X1 U599 ( .A1(n632), .A2(n543), .ZN(n648) );
  NAND2_X1 U600 ( .A1(G77), .A2(n648), .ZN(n545) );
  NOR2_X1 U601 ( .A1(G543), .A2(G651), .ZN(n644) );
  NAND2_X1 U602 ( .A1(G90), .A2(n644), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U605 ( .A1(n548), .A2(n547), .ZN(G171) );
  NAND2_X1 U606 ( .A1(G94), .A2(G452), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT66), .B(n549), .Z(G173) );
  NAND2_X1 U608 ( .A1(G7), .A2(G661), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U610 ( .A(G223), .B(KEYINPUT68), .Z(n813) );
  NAND2_X1 U611 ( .A1(n813), .A2(G567), .ZN(n551) );
  XOR2_X1 U612 ( .A(KEYINPUT11), .B(n551), .Z(G234) );
  NAND2_X1 U613 ( .A1(n644), .A2(G81), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n552), .B(KEYINPUT12), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G68), .A2(n648), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U617 ( .A(n555), .B(KEYINPUT13), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G43), .A2(n645), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n652), .A2(G56), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n558), .Z(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT69), .B(n561), .Z(n918) );
  NAND2_X1 U624 ( .A1(n918), .A2(G860), .ZN(G153) );
  INV_X1 U625 ( .A(G171), .ZN(G301) );
  NAND2_X1 U626 ( .A1(G868), .A2(G301), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n652), .A2(G66), .ZN(n563) );
  NAND2_X1 U628 ( .A1(G54), .A2(n645), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G79), .A2(n648), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G92), .A2(n644), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT15), .ZN(n917) );
  INV_X1 U635 ( .A(G868), .ZN(n594) );
  NAND2_X1 U636 ( .A1(n917), .A2(n594), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(G284) );
  NAND2_X1 U638 ( .A1(n652), .A2(G63), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G51), .A2(n645), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(KEYINPUT6), .B(n573), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n644), .A2(G89), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G76), .A2(n648), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U646 ( .A(KEYINPUT5), .B(n577), .Z(n578) );
  XNOR2_X1 U647 ( .A(KEYINPUT70), .B(n578), .ZN(n579) );
  NOR2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U649 ( .A(KEYINPUT7), .B(n581), .Z(G168) );
  XNOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .ZN(n582) );
  XNOR2_X1 U651 ( .A(n582), .B(KEYINPUT71), .ZN(G286) );
  NAND2_X1 U652 ( .A1(n652), .A2(G65), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G53), .A2(n645), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G78), .A2(n648), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G91), .A2(n644), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n902) );
  INV_X1 U659 ( .A(n902), .ZN(G299) );
  NOR2_X1 U660 ( .A1(G286), .A2(n594), .ZN(n590) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(G297) );
  INV_X1 U663 ( .A(G860), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n591), .A2(G559), .ZN(n592) );
  INV_X1 U665 ( .A(n917), .ZN(n880) );
  NAND2_X1 U666 ( .A1(n592), .A2(n880), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U668 ( .A1(n918), .A2(n594), .ZN(n595) );
  XOR2_X1 U669 ( .A(KEYINPUT72), .B(n595), .Z(n598) );
  NAND2_X1 U670 ( .A1(G868), .A2(n880), .ZN(n596) );
  NOR2_X1 U671 ( .A1(G559), .A2(n596), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G123), .A2(n854), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT18), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G135), .A2(n859), .ZN(n600) );
  XOR2_X1 U676 ( .A(KEYINPUT73), .B(n600), .Z(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G99), .A2(n858), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G111), .A2(n855), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n990) );
  XOR2_X1 U682 ( .A(G2096), .B(n990), .Z(n607) );
  NOR2_X1 U683 ( .A1(G2100), .A2(n607), .ZN(n608) );
  XOR2_X1 U684 ( .A(KEYINPUT74), .B(n608), .Z(G156) );
  NAND2_X1 U685 ( .A1(n652), .A2(G67), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G55), .A2(n645), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G80), .A2(n648), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G93), .A2(n644), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U691 ( .A(KEYINPUT77), .B(n613), .Z(n614) );
  NOR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n659) );
  NAND2_X1 U693 ( .A1(G559), .A2(n880), .ZN(n616) );
  XOR2_X1 U694 ( .A(n918), .B(n616), .Z(n662) );
  XOR2_X1 U695 ( .A(n662), .B(KEYINPUT75), .Z(n617) );
  NOR2_X1 U696 ( .A1(G860), .A2(n617), .ZN(n618) );
  XOR2_X1 U697 ( .A(KEYINPUT76), .B(n618), .Z(n619) );
  XOR2_X1 U698 ( .A(n659), .B(n619), .Z(G145) );
  NAND2_X1 U699 ( .A1(G61), .A2(n652), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G86), .A2(n644), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G48), .A2(n645), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n648), .A2(G73), .ZN(n622) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n627), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G49), .A2(n645), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n628), .B(KEYINPUT78), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U712 ( .A1(n652), .A2(n631), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G87), .A2(n632), .ZN(n633) );
  XOR2_X1 U714 ( .A(KEYINPUT79), .B(n633), .Z(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U716 ( .A1(n644), .A2(G88), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT81), .B(n636), .Z(n638) );
  NAND2_X1 U718 ( .A1(n648), .A2(G75), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U720 ( .A(KEYINPUT82), .B(n639), .Z(n643) );
  NAND2_X1 U721 ( .A1(n645), .A2(G50), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n652), .A2(G62), .ZN(n640) );
  AND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U725 ( .A(G303), .ZN(G166) );
  NAND2_X1 U726 ( .A1(G85), .A2(n644), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G47), .A2(n645), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G72), .A2(n648), .ZN(n649) );
  XNOR2_X1 U730 ( .A(KEYINPUT65), .B(n649), .ZN(n650) );
  NOR2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U732 ( .A1(n652), .A2(G60), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n654), .A2(n653), .ZN(G290) );
  NOR2_X1 U734 ( .A1(G868), .A2(n659), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(KEYINPUT83), .ZN(n665) );
  XNOR2_X1 U736 ( .A(G288), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n902), .B(G166), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n660), .B(G290), .ZN(n661) );
  XNOR2_X1 U741 ( .A(G305), .B(n661), .ZN(n879) );
  XNOR2_X1 U742 ( .A(n879), .B(n662), .ZN(n663) );
  NAND2_X1 U743 ( .A1(G868), .A2(n663), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n667), .ZN(n669) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G2072), .A2(n670), .ZN(G158) );
  NAND2_X1 U751 ( .A1(G661), .A2(G483), .ZN(n671) );
  XNOR2_X1 U752 ( .A(KEYINPUT85), .B(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n672), .A2(G319), .ZN(n673) );
  XOR2_X1 U754 ( .A(KEYINPUT86), .B(n673), .Z(n819) );
  NAND2_X1 U755 ( .A1(G36), .A2(n819), .ZN(G176) );
  NAND2_X1 U756 ( .A1(G102), .A2(n858), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G138), .A2(n859), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U759 ( .A1(G126), .A2(n854), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G114), .A2(n855), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U762 ( .A1(n679), .A2(n678), .ZN(G164) );
  XNOR2_X1 U763 ( .A(G1986), .B(G290), .ZN(n920) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n708) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n708), .A2(n707), .ZN(n808) );
  NAND2_X1 U767 ( .A1(n920), .A2(n808), .ZN(n795) );
  XNOR2_X1 U768 ( .A(KEYINPUT37), .B(G2067), .ZN(n806) );
  NAND2_X1 U769 ( .A1(G104), .A2(n858), .ZN(n681) );
  NAND2_X1 U770 ( .A1(G140), .A2(n859), .ZN(n680) );
  NAND2_X1 U771 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n682), .ZN(n689) );
  NAND2_X1 U773 ( .A1(n854), .A2(G128), .ZN(n683) );
  XNOR2_X1 U774 ( .A(KEYINPUT87), .B(n683), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n855), .A2(G116), .ZN(n684) );
  XOR2_X1 U776 ( .A(KEYINPUT88), .B(n684), .Z(n685) );
  NOR2_X1 U777 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U778 ( .A(n687), .B(KEYINPUT35), .ZN(n688) );
  NOR2_X1 U779 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U780 ( .A(KEYINPUT36), .B(n690), .ZN(n869) );
  NOR2_X1 U781 ( .A1(n806), .A2(n869), .ZN(n989) );
  NAND2_X1 U782 ( .A1(n808), .A2(n989), .ZN(n804) );
  NAND2_X1 U783 ( .A1(G105), .A2(n858), .ZN(n691) );
  XNOR2_X1 U784 ( .A(n691), .B(KEYINPUT38), .ZN(n698) );
  NAND2_X1 U785 ( .A1(G141), .A2(n859), .ZN(n693) );
  NAND2_X1 U786 ( .A1(G129), .A2(n854), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n855), .A2(G117), .ZN(n694) );
  XOR2_X1 U789 ( .A(KEYINPUT90), .B(n694), .Z(n695) );
  NOR2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U792 ( .A1(n872), .A2(G1996), .ZN(n991) );
  NAND2_X1 U793 ( .A1(G119), .A2(n854), .ZN(n700) );
  NAND2_X1 U794 ( .A1(G107), .A2(n855), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n705) );
  NAND2_X1 U796 ( .A1(G95), .A2(n858), .ZN(n702) );
  NAND2_X1 U797 ( .A1(G131), .A2(n859), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U799 ( .A(KEYINPUT89), .B(n703), .Z(n704) );
  NOR2_X1 U800 ( .A1(n705), .A2(n704), .ZN(n868) );
  INV_X1 U801 ( .A(G1991), .ZN(n797) );
  NOR2_X1 U802 ( .A1(n868), .A2(n797), .ZN(n998) );
  OR2_X1 U803 ( .A1(n991), .A2(n998), .ZN(n706) );
  NAND2_X1 U804 ( .A1(n808), .A2(n706), .ZN(n796) );
  NAND2_X1 U805 ( .A1(n804), .A2(n796), .ZN(n793) );
  XNOR2_X1 U806 ( .A(KEYINPUT91), .B(n707), .ZN(n709) );
  NAND2_X2 U807 ( .A1(n709), .A2(n708), .ZN(n755) );
  NAND2_X1 U808 ( .A1(G8), .A2(n755), .ZN(n789) );
  XOR2_X1 U809 ( .A(G1961), .B(KEYINPUT92), .Z(n932) );
  NAND2_X1 U810 ( .A1(n932), .A2(n755), .ZN(n710) );
  XNOR2_X1 U811 ( .A(n710), .B(KEYINPUT93), .ZN(n713) );
  XOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .Z(n972) );
  INV_X1 U813 ( .A(n711), .ZN(n723) );
  NOR2_X1 U814 ( .A1(n972), .A2(n711), .ZN(n712) );
  NOR2_X1 U815 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U816 ( .A(KEYINPUT95), .B(n714), .ZN(n749) );
  NAND2_X1 U817 ( .A1(n749), .A2(G171), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n711), .A2(G1956), .ZN(n715) );
  XOR2_X1 U819 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n717) );
  NAND2_X1 U820 ( .A1(n723), .A2(G2072), .ZN(n716) );
  XOR2_X1 U821 ( .A(n717), .B(n716), .Z(n718) );
  NOR2_X1 U822 ( .A1(n722), .A2(n902), .ZN(n721) );
  XOR2_X1 U823 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n720) );
  XNOR2_X1 U824 ( .A(n721), .B(n720), .ZN(n743) );
  NAND2_X1 U825 ( .A1(n722), .A2(n902), .ZN(n741) );
  NAND2_X1 U826 ( .A1(G2067), .A2(n723), .ZN(n724) );
  XNOR2_X1 U827 ( .A(KEYINPUT102), .B(n724), .ZN(n727) );
  NAND2_X1 U828 ( .A1(G1348), .A2(n755), .ZN(n725) );
  XOR2_X1 U829 ( .A(KEYINPUT101), .B(n725), .Z(n726) );
  NAND2_X1 U830 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U831 ( .A1(n917), .A2(n728), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n728), .A2(n917), .ZN(n733) );
  INV_X1 U833 ( .A(n755), .ZN(n729) );
  NAND2_X1 U834 ( .A1(n729), .A2(G1996), .ZN(n730) );
  XOR2_X1 U835 ( .A(KEYINPUT99), .B(n730), .Z(n731) );
  XNOR2_X1 U836 ( .A(n731), .B(KEYINPUT26), .ZN(n732) );
  NAND2_X1 U837 ( .A1(n733), .A2(n732), .ZN(n737) );
  NAND2_X1 U838 ( .A1(n755), .A2(G1341), .ZN(n734) );
  XNOR2_X1 U839 ( .A(n734), .B(KEYINPUT100), .ZN(n735) );
  NAND2_X1 U840 ( .A1(n735), .A2(n918), .ZN(n736) );
  NOR2_X1 U841 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U842 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U843 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U844 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U845 ( .A1(n745), .A2(n522), .ZN(n754) );
  NOR2_X1 U846 ( .A1(G1966), .A2(n789), .ZN(n765) );
  NOR2_X1 U847 ( .A1(G2084), .A2(n755), .ZN(n764) );
  NOR2_X1 U848 ( .A1(n765), .A2(n764), .ZN(n746) );
  NAND2_X1 U849 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U850 ( .A(KEYINPUT30), .B(n747), .ZN(n748) );
  NOR2_X1 U851 ( .A1(G168), .A2(n748), .ZN(n751) );
  NOR2_X1 U852 ( .A1(G171), .A2(n749), .ZN(n750) );
  NOR2_X1 U853 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U854 ( .A(KEYINPUT31), .B(n752), .Z(n753) );
  NAND2_X1 U855 ( .A1(n754), .A2(n753), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n768), .A2(G286), .ZN(n761) );
  NOR2_X1 U857 ( .A1(G2090), .A2(n755), .ZN(n757) );
  NOR2_X1 U858 ( .A1(G1971), .A2(n789), .ZN(n756) );
  NOR2_X1 U859 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U860 ( .A(n758), .B(KEYINPUT104), .ZN(n759) );
  NAND2_X1 U861 ( .A1(n759), .A2(G303), .ZN(n760) );
  NAND2_X1 U862 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U863 ( .A1(n762), .A2(G8), .ZN(n763) );
  XNOR2_X1 U864 ( .A(n763), .B(KEYINPUT32), .ZN(n771) );
  AND2_X1 U865 ( .A1(G8), .A2(n764), .ZN(n766) );
  NOR2_X1 U866 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U867 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U868 ( .A(KEYINPUT103), .B(n769), .ZN(n770) );
  NAND2_X1 U869 ( .A1(n771), .A2(n770), .ZN(n783) );
  NOR2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n906) );
  NOR2_X1 U871 ( .A1(G1971), .A2(G303), .ZN(n924) );
  NOR2_X1 U872 ( .A1(n906), .A2(n924), .ZN(n772) );
  XOR2_X1 U873 ( .A(KEYINPUT105), .B(n772), .Z(n773) );
  NAND2_X1 U874 ( .A1(n783), .A2(n773), .ZN(n774) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n907) );
  NAND2_X1 U876 ( .A1(n774), .A2(n907), .ZN(n775) );
  NOR2_X1 U877 ( .A1(KEYINPUT33), .A2(n776), .ZN(n779) );
  NAND2_X1 U878 ( .A1(n906), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U879 ( .A1(n777), .A2(n789), .ZN(n778) );
  XOR2_X1 U880 ( .A(G305), .B(G1981), .Z(n911) );
  NAND2_X1 U881 ( .A1(n780), .A2(n911), .ZN(n786) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U883 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U884 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U885 ( .A1(n784), .A2(n789), .ZN(n785) );
  NAND2_X1 U886 ( .A1(n786), .A2(n785), .ZN(n791) );
  NOR2_X1 U887 ( .A1(G305), .A2(G1981), .ZN(n787) );
  XOR2_X1 U888 ( .A(n787), .B(KEYINPUT24), .Z(n788) );
  NOR2_X1 U889 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U890 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n811) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n872), .ZN(n986) );
  INV_X1 U893 ( .A(n796), .ZN(n800) );
  AND2_X1 U894 ( .A1(n797), .A2(n868), .ZN(n994) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U896 ( .A1(n994), .A2(n798), .ZN(n799) );
  NOR2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U898 ( .A(n801), .B(KEYINPUT106), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n986), .A2(n802), .ZN(n803) );
  XNOR2_X1 U900 ( .A(n803), .B(KEYINPUT39), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n806), .A2(n869), .ZN(n1005) );
  NAND2_X1 U903 ( .A1(n807), .A2(n1005), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U906 ( .A(n812), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U907 ( .A1(n813), .A2(G2106), .ZN(n814) );
  XOR2_X1 U908 ( .A(KEYINPUT109), .B(n814), .Z(G217) );
  INV_X1 U909 ( .A(G661), .ZN(n816) );
  NAND2_X1 U910 ( .A1(G2), .A2(G15), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT110), .B(n817), .Z(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G108), .ZN(G238) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  XOR2_X1 U922 ( .A(G2100), .B(G2096), .Z(n823) );
  XNOR2_X1 U923 ( .A(KEYINPUT42), .B(G2678), .ZN(n822) );
  XNOR2_X1 U924 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U925 ( .A(KEYINPUT43), .B(G2090), .Z(n825) );
  XNOR2_X1 U926 ( .A(G2067), .B(G2072), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U928 ( .A(n827), .B(n826), .Z(n829) );
  XNOR2_X1 U929 ( .A(G2078), .B(G2084), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(G227) );
  XOR2_X1 U931 ( .A(G1981), .B(G1971), .Z(n831) );
  XNOR2_X1 U932 ( .A(G1986), .B(G1961), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U934 ( .A(n832), .B(G2474), .Z(n834) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U936 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U937 ( .A(KEYINPUT41), .B(G1976), .Z(n836) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1956), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(G229) );
  NAND2_X1 U941 ( .A1(n854), .A2(G124), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n839), .B(KEYINPUT44), .ZN(n841) );
  NAND2_X1 U943 ( .A1(G112), .A2(n855), .ZN(n840) );
  NAND2_X1 U944 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U945 ( .A1(G100), .A2(n858), .ZN(n843) );
  NAND2_X1 U946 ( .A1(G136), .A2(n859), .ZN(n842) );
  NAND2_X1 U947 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U948 ( .A1(n845), .A2(n844), .ZN(G162) );
  NAND2_X1 U949 ( .A1(G103), .A2(n858), .ZN(n847) );
  NAND2_X1 U950 ( .A1(G139), .A2(n859), .ZN(n846) );
  NAND2_X1 U951 ( .A1(n847), .A2(n846), .ZN(n848) );
  XOR2_X1 U952 ( .A(KEYINPUT111), .B(n848), .Z(n853) );
  NAND2_X1 U953 ( .A1(G127), .A2(n854), .ZN(n850) );
  NAND2_X1 U954 ( .A1(G115), .A2(n855), .ZN(n849) );
  NAND2_X1 U955 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U956 ( .A(KEYINPUT47), .B(n851), .Z(n852) );
  NOR2_X1 U957 ( .A1(n853), .A2(n852), .ZN(n1001) );
  XNOR2_X1 U958 ( .A(G162), .B(n990), .ZN(n866) );
  NAND2_X1 U959 ( .A1(G130), .A2(n854), .ZN(n857) );
  NAND2_X1 U960 ( .A1(G118), .A2(n855), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G106), .A2(n858), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G142), .A2(n859), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U965 ( .A(KEYINPUT45), .B(n862), .Z(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n1001), .B(n867), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n877) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n874) );
  XOR2_X1 U972 ( .A(G160), .B(n872), .Z(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(G164), .B(n875), .Z(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U976 ( .A1(G37), .A2(n878), .ZN(G395) );
  XOR2_X1 U977 ( .A(n879), .B(G286), .Z(n882) );
  XNOR2_X1 U978 ( .A(G171), .B(n880), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U980 ( .A(n918), .B(n883), .Z(n884) );
  NOR2_X1 U981 ( .A1(G37), .A2(n884), .ZN(G397) );
  XNOR2_X1 U982 ( .A(G2438), .B(G2443), .ZN(n894) );
  XOR2_X1 U983 ( .A(G2454), .B(G2430), .Z(n886) );
  XNOR2_X1 U984 ( .A(G2446), .B(KEYINPUT107), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U986 ( .A(G2451), .B(G2427), .Z(n888) );
  XNOR2_X1 U987 ( .A(G1341), .B(G1348), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n890), .B(n889), .Z(n892) );
  XNOR2_X1 U990 ( .A(G2435), .B(KEYINPUT108), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n895), .A2(G14), .ZN(n901) );
  NAND2_X1 U994 ( .A1(G319), .A2(n901), .ZN(n898) );
  NOR2_X1 U995 ( .A1(G227), .A2(G229), .ZN(n896) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(n901), .ZN(G401) );
  XNOR2_X1 U1002 ( .A(KEYINPUT56), .B(G16), .ZN(n931) );
  XNOR2_X1 U1003 ( .A(n902), .B(G1956), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(G171), .B(G1961), .ZN(n903) );
  NAND2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n905) );
  NOR2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n915) );
  XOR2_X1 U1008 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n913) );
  XNOR2_X1 U1009 ( .A(G1966), .B(G168), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(n909), .B(KEYINPUT118), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1012 ( .A(n913), .B(n912), .Z(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n929) );
  XOR2_X1 U1014 ( .A(G1348), .B(KEYINPUT120), .Z(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n922) );
  XOR2_X1 U1016 ( .A(n918), .B(G1341), .Z(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n927) );
  AND2_X1 U1019 ( .A1(G303), .A2(G1971), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(KEYINPUT121), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n1018) );
  XNOR2_X1 U1025 ( .A(G5), .B(n932), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(n933), .B(KEYINPUT122), .ZN(n956) );
  XNOR2_X1 U1027 ( .A(KEYINPUT59), .B(G1348), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(n934), .B(G4), .ZN(n942) );
  XOR2_X1 U1029 ( .A(G1341), .B(G19), .Z(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT123), .B(n935), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G6), .B(G1981), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT124), .B(n938), .Z(n940) );
  XNOR2_X1 U1034 ( .A(G1956), .B(G20), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(KEYINPUT60), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(KEYINPUT125), .ZN(n947) );
  XOR2_X1 U1039 ( .A(G1966), .B(KEYINPUT126), .Z(n945) );
  XNOR2_X1 U1040 ( .A(G21), .B(n945), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n954) );
  XNOR2_X1 U1042 ( .A(G1971), .B(G22), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G23), .B(G1976), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n951) );
  XOR2_X1 U1045 ( .A(G1986), .B(G24), .Z(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(KEYINPUT58), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n958), .B(n957), .ZN(n960) );
  INV_X1 U1052 ( .A(G16), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n961), .A2(G11), .ZN(n1016) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(KEYINPUT116), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n962), .B(G34), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G2084), .B(n963), .ZN(n981) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G35), .ZN(n978) );
  XNOR2_X1 U1059 ( .A(G1991), .B(G25), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n971) );
  XOR2_X1 U1062 ( .A(G2067), .B(G26), .Z(n966) );
  NAND2_X1 U1063 ( .A1(n966), .A2(G28), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(KEYINPUT114), .B(G1996), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(G32), .B(n967), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n975) );
  XOR2_X1 U1068 ( .A(G27), .B(n972), .Z(n973) );
  XNOR2_X1 U1069 ( .A(KEYINPUT113), .B(n973), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n976), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT115), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT55), .B(n982), .Z(n983) );
  NOR2_X1 U1076 ( .A1(G29), .A2(n983), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(n984), .B(KEYINPUT117), .ZN(n1014) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT51), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n1000) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n996) );
  XOR2_X1 U1083 ( .A(G160), .B(G2084), .Z(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT112), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1008) );
  XOR2_X1 U1089 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(n1004), .B(KEYINPUT50), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(n1009), .B(KEYINPUT52), .ZN(n1011) );
  INV_X1 U1096 ( .A(KEYINPUT55), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(G29), .A2(n1012), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

