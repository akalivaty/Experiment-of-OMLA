

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U549 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X2 U550 ( .A1(n1026), .A2(n629), .ZN(n644) );
  NOR2_X4 U551 ( .A1(n538), .A2(n537), .ZN(G160) );
  INV_X1 U552 ( .A(KEYINPUT17), .ZN(n532) );
  NOR2_X1 U553 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X2 U554 ( .A1(n520), .A2(n584), .ZN(n805) );
  NOR2_X2 U555 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XNOR2_X1 U556 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U557 ( .A(n600), .B(KEYINPUT95), .ZN(n601) );
  NOR2_X1 U558 ( .A1(n618), .A2(n617), .ZN(n619) );
  INV_X1 U559 ( .A(KEYINPUT23), .ZN(n527) );
  NOR2_X1 U560 ( .A1(n681), .A2(n680), .ZN(n516) );
  NOR2_X1 U561 ( .A1(n656), .A2(G299), .ZN(n653) );
  BUF_X2 U562 ( .A(n624), .Z(n664) );
  AND2_X1 U563 ( .A1(n677), .A2(n669), .ZN(n668) );
  INV_X1 U564 ( .A(KEYINPUT32), .ZN(n674) );
  AND2_X1 U565 ( .A1(n727), .A2(n516), .ZN(n728) );
  INV_X1 U566 ( .A(KEYINPUT70), .ZN(n614) );
  XNOR2_X1 U567 ( .A(n615), .B(n614), .ZN(n618) );
  XNOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n700), .A2(G138), .ZN(n543) );
  INV_X1 U570 ( .A(KEYINPUT82), .ZN(n544) );
  XNOR2_X1 U571 ( .A(n528), .B(n527), .ZN(n531) );
  INV_X1 U572 ( .A(KEYINPUT40), .ZN(n767) );
  NOR2_X1 U573 ( .A1(n766), .A2(n765), .ZN(n768) );
  XNOR2_X1 U574 ( .A(n545), .B(n544), .ZN(n546) );
  AND2_X1 U575 ( .A1(n547), .A2(n546), .ZN(G164) );
  INV_X1 U576 ( .A(G651), .ZN(n520) );
  NOR2_X1 U577 ( .A1(G543), .A2(n520), .ZN(n517) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n517), .Z(n810) );
  NAND2_X1 U579 ( .A1(G65), .A2(n810), .ZN(n522) );
  INV_X1 U580 ( .A(n518), .ZN(n519) );
  XNOR2_X1 U581 ( .A(KEYINPUT66), .B(n519), .ZN(n584) );
  NAND2_X1 U582 ( .A1(G78), .A2(n805), .ZN(n521) );
  NAND2_X1 U583 ( .A1(n522), .A2(n521), .ZN(n526) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n806) );
  NAND2_X1 U585 ( .A1(G91), .A2(n806), .ZN(n524) );
  NOR2_X1 U586 ( .A1(G651), .A2(n584), .ZN(n632) );
  BUF_X1 U587 ( .A(n632), .Z(n811) );
  NAND2_X1 U588 ( .A1(G53), .A2(n811), .ZN(n523) );
  NAND2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  OR2_X1 U590 ( .A1(n526), .A2(n525), .ZN(G299) );
  INV_X2 U591 ( .A(G2105), .ZN(n534) );
  AND2_X4 U592 ( .A1(n534), .A2(G2104), .ZN(n898) );
  NAND2_X1 U593 ( .A1(G101), .A2(n898), .ZN(n528) );
  NAND2_X1 U594 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(KEYINPUT65), .ZN(n696) );
  NAND2_X1 U596 ( .A1(n696), .A2(G113), .ZN(n530) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n538) );
  XNOR2_X2 U598 ( .A(n533), .B(n532), .ZN(n700) );
  NAND2_X1 U599 ( .A1(G137), .A2(n700), .ZN(n536) );
  NOR2_X2 U600 ( .A1(G2104), .A2(n534), .ZN(n902) );
  NAND2_X1 U601 ( .A1(G125), .A2(n902), .ZN(n535) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  AND2_X1 U603 ( .A1(n902), .A2(G126), .ZN(n541) );
  NAND2_X1 U604 ( .A1(G114), .A2(n696), .ZN(n539) );
  XNOR2_X1 U605 ( .A(KEYINPUT81), .B(n539), .ZN(n540) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n547) );
  NAND2_X1 U607 ( .A1(G102), .A2(n898), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n805), .A2(G72), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n810), .A2(G60), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G85), .A2(n806), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G47), .A2(n811), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U616 ( .A(KEYINPUT67), .B(n554), .ZN(G290) );
  NAND2_X1 U617 ( .A1(n806), .A2(G89), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G76), .A2(n805), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n558), .B(KEYINPUT5), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G63), .A2(n810), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G51), .A2(n811), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U628 ( .A1(G64), .A2(n810), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G52), .A2(n811), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n805), .A2(G77), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT68), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G90), .A2(n806), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(G171) );
  NAND2_X1 U637 ( .A1(G75), .A2(n805), .ZN(n574) );
  NAND2_X1 U638 ( .A1(G88), .A2(n806), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G62), .A2(n810), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G50), .A2(n811), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(G166) );
  INV_X1 U644 ( .A(G166), .ZN(G303) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(n811), .A2(G49), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT75), .B(n579), .Z(n581) );
  NAND2_X1 U648 ( .A1(G651), .A2(G74), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT76), .B(n582), .ZN(n583) );
  NOR2_X1 U651 ( .A1(n810), .A2(n583), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G87), .A2(n584), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U654 ( .A1(G73), .A2(n805), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT2), .ZN(n594) );
  NAND2_X1 U656 ( .A1(G61), .A2(n810), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G86), .A2(n806), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G48), .A2(n811), .ZN(n590) );
  XNOR2_X1 U660 ( .A(KEYINPUT77), .B(n590), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(G305) );
  XOR2_X1 U663 ( .A(G1986), .B(G290), .Z(n1006) );
  NOR2_X1 U664 ( .A1(G164), .A2(G1384), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G160), .A2(G40), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n598), .A2(n596), .ZN(n595) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT83), .ZN(n764) );
  NOR2_X1 U668 ( .A1(n1006), .A2(n764), .ZN(n749) );
  XOR2_X1 U669 ( .A(KEYINPUT86), .B(n596), .Z(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n624) );
  NAND2_X1 U671 ( .A1(G8), .A2(n624), .ZN(n738) );
  NOR2_X1 U672 ( .A1(G1966), .A2(n738), .ZN(n681) );
  NOR2_X1 U673 ( .A1(G2084), .A2(n664), .ZN(n679) );
  NOR2_X1 U674 ( .A1(n681), .A2(n679), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G8), .A2(n599), .ZN(n602) );
  INV_X1 U676 ( .A(KEYINPUT30), .ZN(n600) );
  NOR2_X1 U677 ( .A1(G168), .A2(n603), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n604), .B(KEYINPUT96), .ZN(n610) );
  INV_X1 U679 ( .A(n664), .ZN(n648) );
  NOR2_X1 U680 ( .A1(n648), .A2(G1961), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT88), .ZN(n607) );
  XOR2_X1 U682 ( .A(KEYINPUT25), .B(G2078), .Z(n930) );
  NOR2_X1 U683 ( .A1(n664), .A2(n930), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(KEYINPUT89), .ZN(n661) );
  NOR2_X1 U686 ( .A1(n661), .A2(G171), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT97), .B(n611), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT31), .ZN(n676) );
  NAND2_X1 U689 ( .A1(G56), .A2(n810), .ZN(n613) );
  XOR2_X1 U690 ( .A(KEYINPUT14), .B(n613), .Z(n621) );
  NAND2_X1 U691 ( .A1(n805), .A2(G68), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n806), .A2(G81), .ZN(n616) );
  XOR2_X1 U693 ( .A(KEYINPUT12), .B(n616), .Z(n617) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT13), .ZN(n620) );
  NOR2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n811), .A2(G43), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n1026) );
  INV_X1 U698 ( .A(G1996), .ZN(n927) );
  NOR2_X1 U699 ( .A1(n624), .A2(n927), .ZN(n626) );
  XOR2_X1 U700 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n625) );
  XNOR2_X1 U701 ( .A(n626), .B(n625), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n664), .A2(G1341), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G66), .A2(n810), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G79), .A2(n805), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n636) );
  NAND2_X1 U707 ( .A1(G92), .A2(n806), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G54), .A2(n632), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U711 ( .A(KEYINPUT15), .B(n637), .Z(n1005) );
  NAND2_X1 U712 ( .A1(n644), .A2(n1005), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n664), .A2(G1348), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n638), .B(KEYINPUT92), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n648), .A2(G2067), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(KEYINPUT93), .ZN(n646) );
  NOR2_X1 U719 ( .A1(n1005), .A2(n644), .ZN(n645) );
  NOR2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n655) );
  NAND2_X1 U721 ( .A1(G1956), .A2(n664), .ZN(n647) );
  XOR2_X1 U722 ( .A(KEYINPUT91), .B(n647), .Z(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT90), .B(KEYINPUT27), .Z(n650) );
  NAND2_X1 U724 ( .A1(G2072), .A2(n648), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n653), .B(KEYINPUT94), .ZN(n654) );
  NOR2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n656), .A2(G299), .ZN(n657) );
  XOR2_X1 U730 ( .A(KEYINPUT28), .B(n657), .Z(n658) );
  NOR2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(KEYINPUT29), .ZN(n663) );
  NAND2_X1 U733 ( .A1(G171), .A2(n661), .ZN(n662) );
  NAND2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n677) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n738), .ZN(n666) );
  NOR2_X1 U736 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n667), .A2(G303), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n676), .A2(n668), .ZN(n673) );
  INV_X1 U740 ( .A(n669), .ZN(n670) );
  OR2_X1 U741 ( .A1(n670), .A2(G286), .ZN(n671) );
  AND2_X1 U742 ( .A1(G8), .A2(n671), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(n729) );
  NAND2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n1018) );
  AND2_X1 U746 ( .A1(n677), .A2(n1018), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n676), .A2(n678), .ZN(n683) );
  INV_X1 U748 ( .A(n1018), .ZN(n687) );
  AND2_X1 U749 ( .A1(G8), .A2(n679), .ZN(n680) );
  OR2_X1 U750 ( .A1(n687), .A2(n516), .ZN(n682) );
  AND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n729), .A2(n684), .ZN(n689) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  NOR2_X1 U755 ( .A1(n685), .A2(n1013), .ZN(n686) );
  NOR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n690), .B(KEYINPUT98), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n691), .A2(n738), .ZN(n692) );
  NOR2_X1 U760 ( .A1(KEYINPUT33), .A2(n692), .ZN(n695) );
  NAND2_X1 U761 ( .A1(n1013), .A2(KEYINPUT33), .ZN(n693) );
  NOR2_X1 U762 ( .A1(n693), .A2(n738), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n726) );
  XOR2_X1 U764 ( .A(G1981), .B(G305), .Z(n1021) );
  BUF_X1 U765 ( .A(n696), .Z(n901) );
  NAND2_X1 U766 ( .A1(G116), .A2(n901), .ZN(n698) );
  NAND2_X1 U767 ( .A1(G128), .A2(n902), .ZN(n697) );
  NAND2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U769 ( .A(n699), .B(KEYINPUT35), .ZN(n705) );
  NAND2_X1 U770 ( .A1(G104), .A2(n898), .ZN(n702) );
  NAND2_X1 U771 ( .A1(G140), .A2(n700), .ZN(n701) );
  NAND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U773 ( .A(KEYINPUT34), .B(n703), .Z(n704) );
  NAND2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n706), .B(KEYINPUT36), .ZN(n894) );
  XOR2_X1 U776 ( .A(G2067), .B(KEYINPUT37), .Z(n751) );
  NAND2_X1 U777 ( .A1(n894), .A2(n751), .ZN(n990) );
  NOR2_X1 U778 ( .A1(n764), .A2(n990), .ZN(n761) );
  INV_X1 U779 ( .A(n761), .ZN(n742) );
  AND2_X1 U780 ( .A1(n1021), .A2(n742), .ZN(n724) );
  NAND2_X1 U781 ( .A1(G95), .A2(n898), .ZN(n708) );
  NAND2_X1 U782 ( .A1(G119), .A2(n902), .ZN(n707) );
  NAND2_X1 U783 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U784 ( .A1(n901), .A2(G107), .ZN(n709) );
  XOR2_X1 U785 ( .A(KEYINPUT84), .B(n709), .Z(n710) );
  NOR2_X1 U786 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U787 ( .A1(n700), .A2(G131), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n893) );
  AND2_X1 U789 ( .A1(n893), .A2(G1991), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G105), .A2(n898), .ZN(n714) );
  XOR2_X1 U791 ( .A(KEYINPUT38), .B(n714), .Z(n719) );
  NAND2_X1 U792 ( .A1(G117), .A2(n901), .ZN(n716) );
  NAND2_X1 U793 ( .A1(G129), .A2(n902), .ZN(n715) );
  NAND2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U795 ( .A(KEYINPUT85), .B(n717), .Z(n718) );
  NOR2_X1 U796 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U797 ( .A1(n700), .A2(G141), .ZN(n720) );
  NAND2_X1 U798 ( .A1(n721), .A2(n720), .ZN(n908) );
  AND2_X1 U799 ( .A1(n908), .A2(G1996), .ZN(n722) );
  NOR2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n987) );
  NOR2_X1 U801 ( .A1(n987), .A2(n764), .ZN(n756) );
  INV_X1 U802 ( .A(n756), .ZN(n744) );
  AND2_X1 U803 ( .A1(n724), .A2(n744), .ZN(n725) );
  AND2_X1 U804 ( .A1(n726), .A2(n725), .ZN(n747) );
  NAND2_X1 U805 ( .A1(n676), .A2(n677), .ZN(n727) );
  NOR2_X1 U806 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U807 ( .A1(G166), .A2(G8), .ZN(n730) );
  NOR2_X1 U808 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U809 ( .A1(n732), .A2(n731), .ZN(n734) );
  INV_X1 U810 ( .A(n738), .ZN(n733) );
  NOR2_X2 U811 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U812 ( .A(n735), .B(KEYINPUT99), .ZN(n741) );
  NOR2_X1 U813 ( .A1(G1981), .A2(G305), .ZN(n736) );
  XOR2_X1 U814 ( .A(n736), .B(KEYINPUT24), .Z(n737) );
  NOR2_X1 U815 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U816 ( .A(KEYINPUT87), .B(n739), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n741), .A2(n740), .ZN(n743) );
  AND2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n745) );
  AND2_X2 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U821 ( .A(n750), .B(KEYINPUT100), .ZN(n766) );
  NOR2_X1 U822 ( .A1(n894), .A2(n751), .ZN(n752) );
  XOR2_X1 U823 ( .A(KEYINPUT103), .B(n752), .Z(n992) );
  NOR2_X1 U824 ( .A1(G1996), .A2(n908), .ZN(n753) );
  XOR2_X1 U825 ( .A(KEYINPUT101), .B(n753), .Z(n980) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n754) );
  NOR2_X1 U827 ( .A1(G1991), .A2(n893), .ZN(n985) );
  NOR2_X1 U828 ( .A1(n754), .A2(n985), .ZN(n755) );
  NOR2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U830 ( .A1(n980), .A2(n757), .ZN(n758) );
  XOR2_X1 U831 ( .A(n758), .B(KEYINPUT102), .Z(n759) );
  XNOR2_X1 U832 ( .A(KEYINPUT39), .B(n759), .ZN(n760) );
  NOR2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U834 ( .A1(n992), .A2(n762), .ZN(n763) );
  NOR2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n768), .B(n767), .ZN(G329) );
  XOR2_X1 U837 ( .A(G2438), .B(G2454), .Z(n770) );
  XNOR2_X1 U838 ( .A(G2435), .B(G2430), .ZN(n769) );
  XNOR2_X1 U839 ( .A(n770), .B(n769), .ZN(n771) );
  XOR2_X1 U840 ( .A(n771), .B(KEYINPUT104), .Z(n773) );
  XNOR2_X1 U841 ( .A(G1341), .B(G1348), .ZN(n772) );
  XNOR2_X1 U842 ( .A(n773), .B(n772), .ZN(n777) );
  XOR2_X1 U843 ( .A(G2427), .B(G2443), .Z(n775) );
  XNOR2_X1 U844 ( .A(G2451), .B(G2446), .ZN(n774) );
  XNOR2_X1 U845 ( .A(n775), .B(n774), .ZN(n776) );
  XOR2_X1 U846 ( .A(n777), .B(n776), .Z(n778) );
  AND2_X1 U847 ( .A1(G14), .A2(n778), .ZN(G401) );
  AND2_X1 U848 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U849 ( .A(G57), .ZN(G237) );
  INV_X1 U850 ( .A(G132), .ZN(G219) );
  INV_X1 U851 ( .A(G82), .ZN(G220) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n779) );
  XNOR2_X1 U853 ( .A(n779), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U854 ( .A(G223), .ZN(n843) );
  NAND2_X1 U855 ( .A1(n843), .A2(G567), .ZN(n780) );
  XNOR2_X1 U856 ( .A(n780), .B(KEYINPUT11), .ZN(n781) );
  XNOR2_X1 U857 ( .A(KEYINPUT69), .B(n781), .ZN(G234) );
  INV_X1 U858 ( .A(G860), .ZN(n786) );
  OR2_X1 U859 ( .A1(n1026), .A2(n786), .ZN(G153) );
  INV_X1 U860 ( .A(G171), .ZN(G301) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n783) );
  OR2_X1 U862 ( .A1(n1005), .A2(G868), .ZN(n782) );
  NAND2_X1 U863 ( .A1(n783), .A2(n782), .ZN(G284) );
  INV_X1 U864 ( .A(G868), .ZN(n826) );
  NOR2_X1 U865 ( .A1(G286), .A2(n826), .ZN(n785) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n784) );
  NOR2_X1 U867 ( .A1(n785), .A2(n784), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n786), .A2(G559), .ZN(n787) );
  NAND2_X1 U869 ( .A1(n787), .A2(n1005), .ZN(n788) );
  XNOR2_X1 U870 ( .A(n788), .B(KEYINPUT71), .ZN(n789) );
  XOR2_X1 U871 ( .A(KEYINPUT16), .B(n789), .Z(G148) );
  NAND2_X1 U872 ( .A1(n1005), .A2(G868), .ZN(n790) );
  XNOR2_X1 U873 ( .A(KEYINPUT72), .B(n790), .ZN(n791) );
  NOR2_X1 U874 ( .A1(G559), .A2(n791), .ZN(n793) );
  NOR2_X1 U875 ( .A1(G868), .A2(n1026), .ZN(n792) );
  NOR2_X1 U876 ( .A1(n793), .A2(n792), .ZN(G282) );
  NAND2_X1 U877 ( .A1(G99), .A2(n898), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G111), .A2(n901), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n796), .B(KEYINPUT73), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G135), .A2(n700), .ZN(n797) );
  NAND2_X1 U882 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U883 ( .A1(n902), .A2(G123), .ZN(n799) );
  XOR2_X1 U884 ( .A(KEYINPUT18), .B(n799), .Z(n800) );
  NOR2_X1 U885 ( .A1(n801), .A2(n800), .ZN(n989) );
  XNOR2_X1 U886 ( .A(n989), .B(G2096), .ZN(n803) );
  INV_X1 U887 ( .A(G2100), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n803), .A2(n802), .ZN(G156) );
  NAND2_X1 U889 ( .A1(G559), .A2(n1005), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n1026), .B(n804), .ZN(n823) );
  NOR2_X1 U891 ( .A1(n823), .A2(G860), .ZN(n816) );
  NAND2_X1 U892 ( .A1(G80), .A2(n805), .ZN(n808) );
  NAND2_X1 U893 ( .A1(G93), .A2(n806), .ZN(n807) );
  NAND2_X1 U894 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U895 ( .A(KEYINPUT74), .B(n809), .ZN(n815) );
  NAND2_X1 U896 ( .A1(G67), .A2(n810), .ZN(n813) );
  NAND2_X1 U897 ( .A1(G55), .A2(n811), .ZN(n812) );
  NAND2_X1 U898 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U899 ( .A1(n815), .A2(n814), .ZN(n825) );
  XNOR2_X1 U900 ( .A(n816), .B(n825), .ZN(G145) );
  XNOR2_X1 U901 ( .A(n825), .B(G288), .ZN(n822) );
  XNOR2_X1 U902 ( .A(KEYINPUT19), .B(KEYINPUT78), .ZN(n818) );
  XNOR2_X1 U903 ( .A(G305), .B(G166), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U905 ( .A(n819), .B(G290), .Z(n820) );
  XNOR2_X1 U906 ( .A(G299), .B(n820), .ZN(n821) );
  XNOR2_X1 U907 ( .A(n822), .B(n821), .ZN(n849) );
  XOR2_X1 U908 ( .A(n823), .B(n849), .Z(n824) );
  NAND2_X1 U909 ( .A1(n824), .A2(G868), .ZN(n828) );
  NAND2_X1 U910 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U911 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U912 ( .A(KEYINPUT79), .B(n829), .ZN(G295) );
  NAND2_X1 U913 ( .A1(G2078), .A2(G2084), .ZN(n830) );
  XOR2_X1 U914 ( .A(KEYINPUT20), .B(n830), .Z(n831) );
  NAND2_X1 U915 ( .A1(G2090), .A2(n831), .ZN(n833) );
  XNOR2_X1 U916 ( .A(KEYINPUT21), .B(KEYINPUT80), .ZN(n832) );
  XNOR2_X1 U917 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U918 ( .A1(G2072), .A2(n834), .ZN(G158) );
  XNOR2_X1 U919 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U920 ( .A1(G220), .A2(G219), .ZN(n835) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U922 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U923 ( .A1(G96), .A2(n837), .ZN(n847) );
  NAND2_X1 U924 ( .A1(n847), .A2(G2106), .ZN(n841) );
  NAND2_X1 U925 ( .A1(G69), .A2(G120), .ZN(n838) );
  NOR2_X1 U926 ( .A1(G237), .A2(n838), .ZN(n839) );
  NAND2_X1 U927 ( .A1(G108), .A2(n839), .ZN(n848) );
  NAND2_X1 U928 ( .A1(n848), .A2(G567), .ZN(n840) );
  NAND2_X1 U929 ( .A1(n841), .A2(n840), .ZN(n923) );
  NAND2_X1 U930 ( .A1(G661), .A2(G483), .ZN(n842) );
  NOR2_X1 U931 ( .A1(n923), .A2(n842), .ZN(n846) );
  NAND2_X1 U932 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U935 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U937 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n848), .A2(n847), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  XOR2_X1 U944 ( .A(n849), .B(G286), .Z(n851) );
  XNOR2_X1 U945 ( .A(G171), .B(n1005), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n852), .B(n1026), .ZN(n853) );
  NOR2_X1 U948 ( .A1(G37), .A2(n853), .ZN(G397) );
  XOR2_X1 U949 ( .A(G1961), .B(G1971), .Z(n855) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1976), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n865) );
  XOR2_X1 U952 ( .A(G2474), .B(KEYINPUT108), .Z(n857) );
  XNOR2_X1 U953 ( .A(G1991), .B(KEYINPUT41), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U955 ( .A(G1956), .B(G1966), .Z(n859) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1981), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U958 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U959 ( .A(KEYINPUT109), .B(KEYINPUT107), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U961 ( .A(n865), .B(n864), .Z(G229) );
  XOR2_X1 U962 ( .A(G2100), .B(KEYINPUT106), .Z(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U965 ( .A(KEYINPUT42), .B(G2090), .Z(n869) );
  XNOR2_X1 U966 ( .A(G2067), .B(G2072), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U968 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U969 ( .A(G2678), .B(G2096), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U971 ( .A(G2078), .B(G2084), .Z(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(G227) );
  NAND2_X1 U973 ( .A1(G100), .A2(n898), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G136), .A2(n700), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U976 ( .A1(G124), .A2(n902), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n878), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G112), .A2(n901), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n879), .B(KEYINPUT110), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U982 ( .A1(G118), .A2(n901), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G130), .A2(n902), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U985 ( .A1(n898), .A2(G106), .ZN(n886) );
  XOR2_X1 U986 ( .A(KEYINPUT111), .B(n886), .Z(n888) );
  NAND2_X1 U987 ( .A1(n700), .A2(G142), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(KEYINPUT45), .B(n889), .Z(n890) );
  NOR2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U991 ( .A(G164), .B(n892), .ZN(n897) );
  XOR2_X1 U992 ( .A(n894), .B(n893), .Z(n895) );
  XNOR2_X1 U993 ( .A(n895), .B(G162), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n915) );
  NAND2_X1 U995 ( .A1(G103), .A2(n898), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G139), .A2(n700), .ZN(n899) );
  NAND2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n907) );
  NAND2_X1 U998 ( .A1(G115), .A2(n901), .ZN(n904) );
  NAND2_X1 U999 ( .A1(G127), .A2(n902), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1001 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n975) );
  XOR2_X1 U1003 ( .A(n908), .B(n975), .Z(n913) );
  XOR2_X1 U1004 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n910) );
  XNOR2_X1 U1005 ( .A(n989), .B(KEYINPUT112), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(G160), .B(n911), .Z(n912) );
  XOR2_X1 U1008 ( .A(n913), .B(n912), .Z(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G397), .A2(n918), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n923), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT113), .B(n919), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G395), .A2(n920), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n923), .ZN(G319) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(G29), .B(KEYINPUT117), .ZN(n945) );
  XNOR2_X1 U1022 ( .A(G2084), .B(G34), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(KEYINPUT54), .ZN(n942) );
  XNOR2_X1 U1024 ( .A(G2090), .B(G35), .ZN(n939) );
  XOR2_X1 U1025 ( .A(G2072), .B(G33), .Z(n925) );
  NAND2_X1 U1026 ( .A1(n925), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1027 ( .A(KEYINPUT115), .B(G2067), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(n926), .B(G26), .ZN(n934) );
  XOR2_X1 U1029 ( .A(G1991), .B(G25), .Z(n929) );
  XNOR2_X1 U1030 ( .A(n927), .B(G32), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G27), .B(n930), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(KEYINPUT53), .B(n937), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1038 ( .A(KEYINPUT116), .B(n940), .Z(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(KEYINPUT55), .B(n943), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT118), .B(n946), .ZN(n1004) );
  XOR2_X1 U1043 ( .A(G1961), .B(G5), .Z(n959) );
  XOR2_X1 U1044 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n947) );
  XNOR2_X1 U1045 ( .A(KEYINPUT60), .B(n947), .ZN(n957) );
  XOR2_X1 U1046 ( .A(G1348), .B(KEYINPUT59), .Z(n948) );
  XNOR2_X1 U1047 ( .A(G4), .B(n948), .ZN(n955) );
  XOR2_X1 U1048 ( .A(G1956), .B(G20), .Z(n952) );
  XNOR2_X1 U1049 ( .A(G1981), .B(G6), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(G19), .B(G1341), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1053 ( .A(KEYINPUT123), .B(n953), .Z(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(n957), .B(n956), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G21), .B(G1966), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(KEYINPUT126), .B(n962), .ZN(n969) );
  XOR2_X1 U1060 ( .A(G1976), .B(G23), .Z(n966) );
  XNOR2_X1 U1061 ( .A(G1986), .B(G24), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G22), .ZN(n963) );
  NOR2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1065 ( .A(KEYINPUT58), .B(n967), .Z(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(n970), .B(KEYINPUT127), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT61), .B(n971), .ZN(n973) );
  INV_X1 U1069 ( .A(G16), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n974), .A2(G11), .ZN(n1002) );
  XOR2_X1 U1072 ( .A(G2072), .B(n975), .Z(n977) );
  XOR2_X1 U1073 ( .A(G164), .B(G2078), .Z(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1075 ( .A(KEYINPUT50), .B(n978), .Z(n983) );
  XOR2_X1 U1076 ( .A(G2090), .B(G162), .Z(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1078 ( .A(KEYINPUT51), .B(n981), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n995) );
  XOR2_X1 U1080 ( .A(G160), .B(G2084), .Z(n984) );
  NOR2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT114), .B(n996), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(KEYINPUT52), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(KEYINPUT55), .A2(n998), .ZN(n1000) );
  INV_X1 U1090 ( .A(G29), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1033) );
  XOR2_X1 U1094 ( .A(G16), .B(KEYINPUT56), .Z(n1031) );
  XNOR2_X1 U1095 ( .A(n1005), .B(G1348), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G166), .B(G1971), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(G1956), .B(G299), .Z(n1008) );
  XNOR2_X1 U1099 ( .A(KEYINPUT119), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(n1013), .B(KEYINPUT120), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(G1961), .B(G171), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT121), .B(n1020), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(G1966), .B(G168), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(n1023), .B(KEYINPUT57), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(G1341), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(KEYINPUT122), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1117 ( .A(n1034), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

