//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n451, new_n453,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n450));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  INV_X1    g027(.A(new_n451), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n453), .A2(G567), .ZN(G234));
  NAND2_X1  g029(.A1(new_n453), .A2(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  AOI22_X1  g037(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n465), .A3(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(new_n468), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G137), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND3_X1  g057(.A1(new_n476), .A2(G2105), .A3(new_n478), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n479), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n478), .A2(new_n475), .A3(new_n468), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(new_n477), .A3(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n469), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT3), .B(G2104), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT68), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n493), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n477), .A2(G114), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n483), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n502), .A2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  AND2_X1   g084(.A1(G75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT69), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n512), .A2(new_n515), .A3(G50), .A4(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n508), .A2(new_n512), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G88), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n517), .A2(KEYINPUT70), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT70), .B1(new_n517), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(G76), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n508), .B(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n527), .B1(new_n530), .B2(G63), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n526), .B1(new_n525), .B2(new_n532), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT72), .B(G89), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n534), .B1(new_n535), .B2(new_n536), .C1(new_n518), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n533), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n532), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT73), .B(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n518), .A2(new_n542), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n541), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n532), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT74), .B(G81), .Z(new_n549));
  INV_X1    g124(.A(new_n535), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n519), .A2(new_n549), .B1(new_n550), .B2(G43), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n550), .A2(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n519), .A2(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n560), .C1(new_n532), .C2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G168), .ZN(G286));
  OAI21_X1  g138(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  INV_X1    g141(.A(G49), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n518), .A2(new_n566), .B1(new_n535), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G288));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  INV_X1    g146(.A(G48), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n518), .A2(new_n571), .B1(new_n535), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n532), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(G85), .A2(new_n519), .B1(new_n550), .B2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n532), .ZN(G290));
  NAND2_X1  g155(.A1(new_n519), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT10), .Z(new_n582));
  NAND2_X1  g157(.A1(new_n508), .A2(G66), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n532), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(G54), .B2(new_n550), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(G171), .B2(new_n588), .ZN(G284));
  OAI21_X1  g165(.A(new_n589), .B1(G171), .B2(new_n588), .ZN(G321));
  NAND2_X1  g166(.A1(G299), .A2(new_n588), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(G168), .B2(new_n588), .ZN(G297));
  XOR2_X1   g168(.A(G297), .B(KEYINPUT75), .Z(G280));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n582), .B(new_n586), .C1(new_n595), .C2(G860), .ZN(G148));
  INV_X1    g171(.A(new_n552), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(G868), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n587), .A2(G559), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT76), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n598), .B1(new_n600), .B2(G868), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n498), .A2(new_n472), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT12), .Z(new_n604));
  INV_X1    g179(.A(G2100), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n604), .A2(KEYINPUT13), .B1(KEYINPUT77), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(KEYINPUT13), .B2(new_n604), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(KEYINPUT77), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G123), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n477), .A2(G111), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n483), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G135), .B2(new_n488), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT78), .B(G2096), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n616), .ZN(G156));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n620), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n623), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n630), .A2(G14), .A3(new_n631), .ZN(G401));
  XOR2_X1   g207(.A(G2084), .B(G2090), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g212(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT18), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n635), .A2(KEYINPUT79), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(KEYINPUT79), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(new_n637), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n635), .B(KEYINPUT17), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n642), .B(new_n634), .C1(new_n643), .C2(new_n637), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n637), .A3(new_n633), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n639), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(KEYINPUT80), .B(KEYINPUT19), .Z(new_n649));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1956), .B(G2474), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1961), .B(G1966), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT20), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n654), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n656), .B(new_n659), .C1(new_n651), .C2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT81), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G5), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(G171), .B2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT96), .Z(new_n674));
  INV_X1    g249(.A(G1961), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT97), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NAND3_X1  g253(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT26), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n681), .A2(new_n682), .B1(G105), .B2(new_n472), .ZN(new_n683));
  INV_X1    g258(.A(G141), .ZN(new_n684));
  INV_X1    g259(.A(G129), .ZN(new_n685));
  OAI221_X1 g260(.A(new_n683), .B1(new_n479), .B2(new_n684), .C1(new_n685), .C2(new_n483), .ZN(new_n686));
  MUX2_X1   g261(.A(G32), .B(new_n686), .S(G29), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT27), .B(G1996), .Z(new_n688));
  INV_X1    g263(.A(G2084), .ZN(new_n689));
  INV_X1    g264(.A(G34), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(KEYINPUT24), .ZN(new_n691));
  AOI21_X1  g266(.A(G29), .B1(new_n690), .B2(KEYINPUT24), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(KEYINPUT91), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(KEYINPUT91), .B2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n481), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n687), .A2(new_n688), .B1(new_n689), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n678), .A2(KEYINPUT98), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n677), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT89), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(G26), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  INV_X1    g278(.A(G140), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT86), .Z(new_n706));
  INV_X1    g281(.A(G128), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n477), .A2(G116), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n483), .A2(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(new_n695), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(KEYINPUT87), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(KEYINPUT87), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n703), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2067), .ZN(new_n717));
  AOI21_X1  g292(.A(KEYINPUT98), .B1(new_n678), .B2(new_n697), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n699), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G6), .A2(G16), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n576), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT32), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1981), .Z(new_n723));
  NAND2_X1  g298(.A1(G166), .A2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G16), .B2(G22), .ZN(new_n725));
  INV_X1    g300(.A(G1971), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n671), .A2(G23), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n569), .B2(new_n671), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT33), .B(G1976), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n723), .A2(new_n727), .A3(new_n728), .A4(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n695), .A2(G25), .ZN(new_n736));
  INV_X1    g311(.A(G119), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n477), .A2(G107), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n483), .A2(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G131), .B2(new_n488), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n736), .B1(new_n741), .B2(new_n695), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  MUX2_X1   g319(.A(G24), .B(G290), .S(G16), .Z(new_n745));
  INV_X1    g320(.A(G1986), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n734), .A2(new_n735), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT36), .Z(new_n749));
  NAND3_X1  g324(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT25), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n488), .B2(G139), .ZN(new_n752));
  NAND2_X1  g327(.A1(G115), .A2(G2104), .ZN(new_n753));
  INV_X1    g328(.A(G127), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n469), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n477), .B1(new_n755), .B2(KEYINPUT90), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT90), .B2(new_n755), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n695), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n695), .B2(G33), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n442), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT92), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n442), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n695), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n695), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n764), .B1(G2078), .B2(new_n766), .C1(new_n687), .C2(new_n688), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n695), .A2(G35), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n695), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2090), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n763), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n671), .A2(G19), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT83), .Z(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n552), .B2(new_n671), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT85), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT84), .B(G1341), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G4), .A2(G16), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT82), .Z(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n587), .B2(new_n671), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1348), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n783), .A2(KEYINPUT95), .A3(G28), .ZN(new_n784));
  AOI21_X1  g359(.A(KEYINPUT95), .B1(new_n783), .B2(G28), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n695), .B1(new_n783), .B2(G28), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT31), .B(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n614), .B2(G29), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n782), .B(new_n789), .C1(new_n696), .C2(new_n689), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n766), .A2(G2078), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n671), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT23), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n790), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(G168), .A2(G16), .ZN(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G21), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(KEYINPUT93), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(KEYINPUT93), .B2(new_n798), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT94), .B(G1966), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n801), .B(new_n802), .Z(new_n803));
  NAND4_X1  g378(.A1(new_n772), .A2(new_n778), .A3(new_n797), .A4(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n719), .A2(new_n749), .A3(new_n804), .ZN(G311));
  INV_X1    g380(.A(G311), .ZN(G150));
  NAND2_X1  g381(.A1(G80), .A2(G543), .ZN(new_n807));
  INV_X1    g382(.A(G67), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n529), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n532), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n810), .B2(new_n809), .ZN(new_n812));
  AOI22_X1  g387(.A1(G93), .A2(new_n519), .B1(new_n550), .B2(G55), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT101), .B(G860), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n812), .A2(new_n813), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(KEYINPUT100), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n552), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n822), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n595), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n818), .B1(new_n829), .B2(new_n815), .ZN(G145));
  INV_X1    g405(.A(G37), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n488), .A2(G142), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n476), .A2(G2105), .A3(new_n478), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G130), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n477), .A2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n832), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT105), .ZN(new_n838));
  INV_X1    g413(.A(new_n604), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n741), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT106), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n501), .A2(KEYINPUT103), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n494), .B1(new_n469), .B2(new_n496), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n498), .A2(KEYINPUT68), .A3(new_n499), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n493), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n506), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n711), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n686), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n851), .B1(new_n854), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n842), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n614), .B(new_n481), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n831), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n841), .B1(new_n856), .B2(KEYINPUT107), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(KEYINPUT107), .B2(new_n856), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n853), .A2(new_n855), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n859), .B1(new_n865), .B2(new_n842), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n862), .A2(KEYINPUT40), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT40), .B1(new_n862), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(G395));
  INV_X1    g445(.A(KEYINPUT110), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n825), .B(new_n600), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n587), .B(G299), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(KEYINPUT41), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n569), .B(G290), .ZN(new_n880));
  NAND2_X1  g455(.A1(G166), .A2(new_n576), .ZN(new_n881));
  NAND2_X1  g456(.A1(G303), .A2(G305), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT108), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n882), .A3(new_n881), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT109), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n887), .A2(KEYINPUT42), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(KEYINPUT42), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n879), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n875), .A3(new_n878), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G868), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n819), .A2(G868), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n871), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI211_X1 g472(.A(KEYINPUT110), .B(new_n895), .C1(new_n893), .C2(G868), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(G295));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n896), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT112), .ZN(new_n902));
  OAI21_X1  g477(.A(G168), .B1(G301), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G301), .A2(new_n902), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n825), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n874), .ZN(new_n907));
  INV_X1    g482(.A(new_n905), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n825), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n823), .B2(new_n824), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n876), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n884), .A2(new_n886), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(KEYINPUT113), .A3(new_n831), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n907), .A2(new_n887), .A3(new_n911), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT113), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n887), .B1(new_n907), .B2(new_n911), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(G37), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n914), .A2(new_n831), .A3(new_n916), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n901), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n915), .A2(new_n916), .A3(new_n921), .ZN(new_n926));
  INV_X1    g501(.A(new_n917), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n920), .A2(G37), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n926), .A2(new_n927), .B1(new_n928), .B2(new_n918), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n925), .B1(new_n929), .B2(new_n901), .ZN(G397));
  NOR2_X1   g505(.A1(new_n504), .A2(new_n505), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n833), .B2(G126), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n846), .A2(new_n847), .A3(new_n493), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n847), .B1(new_n846), .B2(new_n493), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(G160), .A2(G40), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n941), .A2(KEYINPUT114), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(KEYINPUT114), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT46), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n711), .B(G2067), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n944), .B1(new_n686), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  INV_X1    g527(.A(new_n944), .ZN(new_n953));
  OR3_X1    g528(.A1(new_n953), .A2(G1986), .A3(G290), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n686), .B(new_n945), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n741), .A2(new_n743), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n741), .A2(new_n743), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n948), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n954), .A2(new_n955), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n954), .A2(new_n955), .ZN(new_n962));
  AND4_X1   g537(.A1(new_n743), .A2(new_n948), .A3(new_n741), .A4(new_n956), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n711), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n961), .A2(new_n962), .B1(new_n953), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n952), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n849), .B2(G1384), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n935), .A2(KEYINPUT115), .A3(new_n936), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n932), .B2(new_n501), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT116), .B1(new_n973), .B2(new_n970), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n936), .B1(new_n502), .B2(new_n506), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT50), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n938), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n675), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n935), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(new_n938), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G2078), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n937), .B2(new_n939), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n975), .A2(new_n939), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n981), .A2(new_n938), .A3(new_n443), .A4(new_n987), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n982), .A2(new_n986), .B1(new_n988), .B2(new_n983), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n980), .A2(new_n989), .A3(G301), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n979), .A2(new_n675), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n849), .A2(new_n968), .A3(G1384), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n935), .B2(new_n936), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n939), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G160), .A2(G40), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(KEYINPUT45), .B2(new_n973), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n997), .A3(new_n984), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n988), .A2(new_n983), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(G171), .B1(new_n992), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT124), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n980), .A2(new_n989), .A3(new_n1002), .A4(G301), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n991), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT125), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(KEYINPUT125), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n969), .B2(new_n971), .ZN(new_n1011));
  INV_X1    g586(.A(new_n997), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n802), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT118), .B(G2084), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n996), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n972), .A2(new_n1014), .A3(new_n978), .A4(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n972), .A2(new_n978), .A3(new_n1016), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT119), .ZN(new_n1020));
  AOI21_X1  g595(.A(G168), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(G168), .A3(new_n1013), .A4(new_n1017), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT51), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1025), .A3(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT122), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n980), .A2(G301), .A3(new_n999), .A4(new_n998), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n980), .A2(new_n989), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT54), .B(new_n1029), .C1(new_n1030), .C2(G301), .ZN(new_n1031));
  AND3_X1   g606(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n973), .A2(new_n1035), .A3(new_n970), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n970), .B(new_n936), .C1(new_n502), .C2(new_n506), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT117), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n938), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n970), .B1(new_n969), .B2(new_n971), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G2090), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n981), .A2(new_n938), .A3(new_n987), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1042), .A2(new_n1043), .B1(new_n726), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n972), .A2(new_n1043), .A3(new_n938), .A4(new_n978), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(new_n726), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1046), .B(new_n1034), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n969), .A2(new_n938), .A3(new_n971), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n569), .A2(G1976), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(G8), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n576), .B(G1981), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1055), .A2(KEYINPUT49), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(KEYINPUT49), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1051), .A2(new_n1056), .A3(G8), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n569), .B2(G1976), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1054), .B(new_n1058), .C1(new_n1053), .C2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1050), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1031), .A2(new_n1047), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1348), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n979), .A2(new_n1064), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n964), .A2(new_n969), .A3(new_n938), .A4(new_n971), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(KEYINPUT60), .A3(new_n587), .A4(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(G1341), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1051), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(G1996), .B2(new_n1044), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(KEYINPUT59), .A3(new_n552), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n981), .A2(new_n938), .A3(new_n987), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1075), .A2(new_n945), .B1(new_n1051), .B2(new_n1070), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1076), .B2(new_n597), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1068), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1066), .B1(new_n979), .B2(new_n1064), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n587), .B1(new_n1082), .B2(KEYINPUT60), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT61), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n795), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1086));
  XOR2_X1   g661(.A(G299), .B(KEYINPUT57), .Z(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1075), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1087), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1078), .A2(new_n1084), .A3(new_n1092), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1082), .A2(new_n587), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1099), .B2(new_n1091), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1063), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1024), .A2(new_n1026), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1010), .A2(new_n1028), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1050), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1051), .A2(G8), .ZN(new_n1106));
  NOR2_X1   g681(.A1(G305), .A2(G1981), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G288), .A2(G1976), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1058), .B2(new_n1108), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1105), .A2(new_n1061), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1046), .B(G286), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1062), .A2(new_n1047), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1034), .B1(new_n1116), .B2(new_n1046), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1112), .A2(KEYINPUT63), .A3(new_n1062), .A4(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1110), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1104), .A2(KEYINPUT126), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT126), .B1(new_n1104), .B2(new_n1119), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1024), .A2(new_n1026), .A3(new_n1102), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1102), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1028), .A2(KEYINPUT62), .A3(new_n1103), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1114), .A2(new_n1001), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1120), .A2(new_n1121), .A3(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(G290), .B(new_n746), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n953), .B1(new_n960), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n967), .B1(new_n1129), .B2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g707(.A(G319), .ZN(new_n1134));
  NOR3_X1   g708(.A1(G401), .A2(new_n1134), .A3(G227), .ZN(new_n1135));
  NAND3_X1  g709(.A1(new_n668), .A2(new_n669), .A3(new_n1135), .ZN(new_n1136));
  XOR2_X1   g710(.A(new_n1136), .B(KEYINPUT127), .Z(new_n1137));
  INV_X1    g711(.A(new_n867), .ZN(new_n1138));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1138), .B2(new_n861), .ZN(new_n1139));
  NOR2_X1   g713(.A1(new_n929), .A2(new_n1139), .ZN(G308));
  OR2_X1    g714(.A1(new_n929), .A2(new_n1139), .ZN(G225));
endmodule


