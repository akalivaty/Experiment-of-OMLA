

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810;

  AND2_X1 U378 ( .A1(n437), .A2(n436), .ZN(n435) );
  BUF_X1 U379 ( .A(n639), .Z(n358) );
  XNOR2_X1 U380 ( .A(n580), .B(n579), .ZN(n615) );
  NAND2_X1 U381 ( .A1(n659), .A2(n709), .ZN(n660) );
  XNOR2_X1 U382 ( .A(n661), .B(n498), .ZN(n727) );
  NOR2_X1 U383 ( .A1(n381), .A2(n639), .ZN(n657) );
  XNOR2_X1 U384 ( .A(G472), .B(KEYINPUT6), .ZN(n360) );
  NOR2_X1 U385 ( .A1(n773), .A2(G902), .ZN(n558) );
  XNOR2_X1 U386 ( .A(n566), .B(n428), .ZN(n597) );
  INV_X1 U387 ( .A(KEYINPUT75), .ZN(n459) );
  INV_X1 U388 ( .A(G113), .ZN(n460) );
  NAND2_X1 U389 ( .A1(n359), .A2(n393), .ZN(n690) );
  NAND2_X1 U390 ( .A1(n391), .A2(n392), .ZN(n359) );
  AND2_X2 U391 ( .A1(n448), .A2(n462), .ZN(n461) );
  XNOR2_X1 U392 ( .A(n540), .B(n360), .ZN(n656) );
  INV_X2 U393 ( .A(G125), .ZN(n430) );
  XNOR2_X2 U394 ( .A(n495), .B(KEYINPUT40), .ZN(n808) );
  XNOR2_X1 U395 ( .A(n597), .B(n551), .ZN(n791) );
  XNOR2_X2 U396 ( .A(G110), .B(KEYINPUT94), .ZN(n423) );
  NOR2_X1 U397 ( .A1(n358), .A2(n452), .ZN(n618) );
  NAND2_X1 U398 ( .A1(n368), .A2(n369), .ZN(n567) );
  INV_X1 U399 ( .A(G953), .ZN(n798) );
  NOR2_X1 U400 ( .A1(n507), .A2(n506), .ZN(n508) );
  NOR2_X1 U401 ( .A1(n509), .A2(n522), .ZN(n507) );
  XNOR2_X1 U402 ( .A(n501), .B(n382), .ZN(n625) );
  XNOR2_X2 U403 ( .A(n543), .B(n780), .ZN(n562) );
  INV_X1 U404 ( .A(G128), .ZN(n367) );
  INV_X1 U405 ( .A(KEYINPUT68), .ZN(n472) );
  INV_X1 U406 ( .A(G143), .ZN(n366) );
  NOR2_X1 U407 ( .A1(n625), .A2(n482), .ZN(n481) );
  NOR2_X1 U408 ( .A1(n625), .A2(n622), .ZN(n623) );
  XNOR2_X1 U409 ( .A(KEYINPUT96), .B(n583), .ZN(n700) );
  NOR2_X1 U410 ( .A1(n615), .A2(n735), .ZN(n516) );
  INV_X1 U411 ( .A(n473), .ZN(n708) );
  NAND2_X1 U412 ( .A1(n727), .A2(n726), .ZN(n730) );
  XNOR2_X1 U413 ( .A(n612), .B(n611), .ZN(n735) );
  XNOR2_X1 U414 ( .A(n658), .B(KEYINPUT104), .ZN(n711) );
  NOR2_X1 U415 ( .A1(n617), .A2(n616), .ZN(n645) );
  NOR2_X1 U416 ( .A1(n737), .A2(n738), .ZN(n582) );
  AND2_X1 U417 ( .A1(n397), .A2(n398), .ZN(n391) );
  NAND2_X1 U418 ( .A1(n530), .A2(n529), .ZN(n793) );
  XNOR2_X1 U419 ( .A(n488), .B(n590), .ZN(n771) );
  XNOR2_X1 U420 ( .A(G134), .B(n567), .ZN(n528) );
  XNOR2_X1 U421 ( .A(n555), .B(KEYINPUT88), .ZN(n675) );
  XNOR2_X1 U422 ( .A(n429), .B(KEYINPUT70), .ZN(n428) );
  XNOR2_X1 U423 ( .A(n459), .B(KEYINPUT16), .ZN(n458) );
  XNOR2_X1 U424 ( .A(G110), .B(G104), .ZN(n541) );
  INV_X1 U425 ( .A(KEYINPUT47), .ZN(n470) );
  XOR2_X1 U426 ( .A(G116), .B(G107), .Z(n589) );
  XNOR2_X1 U427 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n552) );
  NAND2_X1 U428 ( .A1(n435), .A2(n433), .ZN(n361) );
  NAND2_X1 U429 ( .A1(n435), .A2(n433), .ZN(n717) );
  BUF_X1 U430 ( .A(n690), .Z(n362) );
  AND2_X1 U431 ( .A1(n363), .A2(n364), .ZN(n490) );
  XNOR2_X1 U432 ( .A(n403), .B(n670), .ZN(n363) );
  XOR2_X1 U433 ( .A(KEYINPUT80), .B(n677), .Z(n364) );
  INV_X1 U434 ( .A(n720), .ZN(n365) );
  NAND2_X1 U435 ( .A1(G143), .A2(n367), .ZN(n368) );
  NAND2_X1 U436 ( .A1(n366), .A2(G128), .ZN(n369) );
  BUF_X1 U437 ( .A(n773), .Z(n370) );
  XNOR2_X1 U438 ( .A(n660), .B(KEYINPUT107), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n660), .B(KEYINPUT107), .ZN(n664) );
  BUF_X1 U440 ( .A(n672), .Z(n372) );
  BUF_X1 U441 ( .A(n661), .Z(n373) );
  BUF_X1 U442 ( .A(n809), .Z(n374) );
  XNOR2_X1 U443 ( .A(n654), .B(KEYINPUT108), .ZN(n809) );
  XNOR2_X1 U444 ( .A(n540), .B(G472), .ZN(n609) );
  INV_X1 U445 ( .A(n624), .ZN(n521) );
  INV_X1 U446 ( .A(KEYINPUT10), .ZN(n429) );
  INV_X1 U447 ( .A(KEYINPUT84), .ZN(n496) );
  AND2_X1 U448 ( .A1(n662), .A2(n439), .ZN(n438) );
  XNOR2_X1 U449 ( .A(n460), .B(G122), .ZN(n602) );
  XNOR2_X1 U450 ( .A(n600), .B(n599), .ZN(n601) );
  INV_X1 U451 ( .A(G140), .ZN(n599) );
  XNOR2_X1 U452 ( .A(G104), .B(KEYINPUT11), .ZN(n594) );
  XOR2_X1 U453 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n595) );
  XNOR2_X1 U454 ( .A(n597), .B(n603), .ZN(n494) );
  INV_X1 U455 ( .A(G113), .ZN(n390) );
  XNOR2_X1 U456 ( .A(KEYINPUT71), .B(G131), .ZN(n604) );
  XNOR2_X1 U457 ( .A(n569), .B(n568), .ZN(n570) );
  INV_X1 U458 ( .A(n730), .ZN(n464) );
  INV_X1 U459 ( .A(KEYINPUT30), .ZN(n487) );
  XNOR2_X1 U460 ( .A(KEYINPUT21), .B(n560), .ZN(n738) );
  XNOR2_X1 U461 ( .A(G137), .B(G113), .ZN(n535) );
  INV_X1 U462 ( .A(G953), .ZN(n478) );
  XNOR2_X1 U463 ( .A(G122), .B(KEYINPUT99), .ZN(n585) );
  XOR2_X1 U464 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n586) );
  INV_X1 U465 ( .A(KEYINPUT39), .ZN(n636) );
  NOR2_X1 U466 ( .A1(n741), .A2(n379), .ZN(n436) );
  INV_X1 U467 ( .A(KEYINPUT106), .ZN(n512) );
  INV_X1 U468 ( .A(KEYINPUT1), .ZN(n517) );
  XNOR2_X1 U469 ( .A(G478), .B(n593), .ZN(n613) );
  OR2_X1 U470 ( .A1(n685), .A2(G902), .ZN(n492) );
  INV_X1 U471 ( .A(KEYINPUT25), .ZN(n484) );
  XNOR2_X1 U472 ( .A(G902), .B(KEYINPUT15), .ZN(n555) );
  AND2_X1 U473 ( .A1(G953), .A2(G902), .ZN(n575) );
  INV_X1 U474 ( .A(n589), .ZN(n400) );
  XNOR2_X1 U475 ( .A(n476), .B(n574), .ZN(n576) );
  NAND2_X1 U476 ( .A1(G234), .A2(G237), .ZN(n574) );
  XNOR2_X1 U477 ( .A(KEYINPUT14), .B(KEYINPUT90), .ZN(n476) );
  OR2_X1 U478 ( .A1(G237), .A2(G902), .ZN(n571) );
  INV_X1 U479 ( .A(KEYINPUT41), .ZN(n467) );
  NOR2_X1 U480 ( .A1(n729), .A2(n467), .ZN(n463) );
  INV_X1 U481 ( .A(KEYINPUT38), .ZN(n498) );
  INV_X1 U482 ( .A(n738), .ZN(n503) );
  XNOR2_X1 U483 ( .A(n494), .B(n493), .ZN(n606) );
  XNOR2_X1 U484 ( .A(n596), .B(n601), .ZN(n493) );
  XOR2_X1 U485 ( .A(G137), .B(G140), .Z(n551) );
  XNOR2_X1 U486 ( .A(n547), .B(n546), .ZN(n549) );
  XNOR2_X1 U487 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U488 ( .A(KEYINPUT92), .ZN(n544) );
  XNOR2_X1 U489 ( .A(n475), .B(n474), .ZN(n759) );
  INV_X1 U490 ( .A(KEYINPUT91), .ZN(n474) );
  NAND2_X1 U491 ( .A1(n576), .A2(G952), .ZN(n475) );
  NOR2_X1 U492 ( .A1(n753), .A2(n432), .ZN(n754) );
  XNOR2_X1 U493 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n611) );
  NOR2_X1 U494 ( .A1(n720), .A2(n479), .ZN(n721) );
  INV_X1 U495 ( .A(n510), .ZN(n723) );
  XNOR2_X1 U496 ( .A(n644), .B(KEYINPUT110), .ZN(n647) );
  AND2_X1 U497 ( .A1(n466), .A2(n465), .ZN(n448) );
  NAND2_X1 U498 ( .A1(n464), .A2(n463), .ZN(n462) );
  NAND2_X1 U499 ( .A1(n729), .A2(n467), .ZN(n465) );
  NOR2_X1 U500 ( .A1(n427), .A2(n640), .ZN(n634) );
  OR2_X2 U501 ( .A1(n647), .A2(n477), .ZN(n473) );
  NAND2_X1 U502 ( .A1(n617), .A2(n613), .ZN(n658) );
  XOR2_X1 U503 ( .A(n539), .B(KEYINPUT62), .Z(n681) );
  XNOR2_X1 U504 ( .A(n591), .B(n592), .ZN(n488) );
  XNOR2_X1 U505 ( .A(n685), .B(KEYINPUT59), .ZN(n687) );
  NAND2_X1 U506 ( .A1(n434), .A2(KEYINPUT36), .ZN(n433) );
  XNOR2_X1 U507 ( .A(n514), .B(n485), .ZN(n803) );
  XNOR2_X1 U508 ( .A(n614), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U509 ( .A(n623), .B(KEYINPUT32), .ZN(n806) );
  INV_X1 U510 ( .A(KEYINPUT102), .ZN(n480) );
  NAND2_X1 U511 ( .A1(n741), .A2(n618), .ZN(n482) );
  NAND2_X1 U512 ( .A1(n389), .A2(n451), .ZN(n450) );
  AND2_X1 U513 ( .A1(n510), .A2(n679), .ZN(n376) );
  XOR2_X1 U514 ( .A(KEYINPUT73), .B(G469), .Z(n377) );
  NOR2_X2 U515 ( .A1(n741), .A2(n742), .ZN(n610) );
  AND2_X1 U516 ( .A1(n388), .A2(n376), .ZN(n378) );
  NOR2_X1 U517 ( .A1(n662), .A2(n439), .ZN(n379) );
  XOR2_X1 U518 ( .A(KEYINPUT13), .B(G475), .Z(n380) );
  OR2_X1 U519 ( .A1(n640), .A2(n738), .ZN(n381) );
  XOR2_X1 U520 ( .A(KEYINPUT74), .B(KEYINPUT22), .Z(n382) );
  XNOR2_X1 U521 ( .A(n768), .B(n767), .ZN(n383) );
  XNOR2_X1 U522 ( .A(n771), .B(KEYINPUT121), .ZN(n384) );
  XOR2_X1 U523 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n385) );
  XOR2_X1 U524 ( .A(KEYINPUT72), .B(KEYINPUT48), .Z(n386) );
  INV_X1 U525 ( .A(KEYINPUT44), .ZN(n522) );
  XOR2_X1 U526 ( .A(KEYINPUT87), .B(n682), .Z(n778) );
  AND2_X1 U527 ( .A1(KEYINPUT65), .A2(n674), .ZN(n387) );
  NAND2_X1 U528 ( .A1(n420), .A2(n675), .ZN(n388) );
  OR2_X1 U529 ( .A1(n615), .A2(n450), .ZN(n583) );
  INV_X1 U530 ( .A(n582), .ZN(n742) );
  XNOR2_X1 U531 ( .A(n619), .B(KEYINPUT25), .ZN(n737) );
  AND2_X1 U532 ( .A1(n806), .A2(KEYINPUT44), .ZN(n506) );
  NAND2_X1 U533 ( .A1(n582), .A2(n643), .ZN(n427) );
  XNOR2_X1 U534 ( .A(n602), .B(n458), .ZN(n457) );
  NAND2_X1 U535 ( .A1(n416), .A2(n440), .ZN(n769) );
  AND2_X1 U536 ( .A1(n650), .A2(n649), .ZN(n418) );
  INV_X1 U537 ( .A(n647), .ZN(n469) );
  AND2_X1 U538 ( .A1(n582), .A2(n643), .ZN(n389) );
  NAND2_X1 U539 ( .A1(n419), .A2(n570), .ZN(n393) );
  INV_X1 U540 ( .A(n570), .ZN(n392) );
  NAND2_X1 U541 ( .A1(n411), .A2(n410), .ZN(n397) );
  NAND2_X1 U542 ( .A1(n395), .A2(n396), .ZN(n398) );
  NAND2_X1 U543 ( .A1(n397), .A2(n398), .ZN(n419) );
  INV_X1 U544 ( .A(n411), .ZN(n395) );
  INV_X1 U545 ( .A(n410), .ZN(n396) );
  NAND2_X1 U546 ( .A1(n457), .A2(n589), .ZN(n401) );
  NAND2_X1 U547 ( .A1(n399), .A2(n400), .ZN(n402) );
  NAND2_X1 U548 ( .A1(n401), .A2(n402), .ZN(n500) );
  INV_X1 U549 ( .A(n457), .ZN(n399) );
  INV_X1 U550 ( .A(n562), .ZN(n410) );
  BUF_X1 U551 ( .A(n748), .Z(n452) );
  INV_X1 U552 ( .A(n452), .ZN(n451) );
  BUF_X1 U553 ( .A(n671), .Z(n403) );
  BUF_X1 U554 ( .A(n411), .Z(n404) );
  XNOR2_X1 U555 ( .A(n390), .B(G122), .ZN(n405) );
  NAND2_X1 U556 ( .A1(n453), .A2(n719), .ZN(n671) );
  XNOR2_X2 U557 ( .A(n619), .B(n484), .ZN(n639) );
  BUF_X1 U558 ( .A(n808), .Z(n406) );
  XNOR2_X1 U559 ( .A(n671), .B(n670), .ZN(n676) );
  NAND2_X1 U560 ( .A1(n416), .A2(n440), .ZN(n407) );
  BUF_X1 U561 ( .A(n805), .Z(n408) );
  INV_X1 U562 ( .A(n479), .ZN(n409) );
  XNOR2_X1 U563 ( .A(n481), .B(n480), .ZN(n805) );
  XNOR2_X1 U564 ( .A(n404), .B(G101), .ZN(n779) );
  XNOR2_X2 U565 ( .A(n500), .B(n412), .ZN(n411) );
  INV_X1 U566 ( .A(n561), .ZN(n412) );
  AND2_X1 U567 ( .A1(n413), .A2(n694), .ZN(G54) );
  XNOR2_X1 U568 ( .A(n770), .B(n383), .ZN(n413) );
  AND2_X1 U569 ( .A1(n414), .A2(n694), .ZN(G63) );
  XNOR2_X1 U570 ( .A(n772), .B(n384), .ZN(n414) );
  NAND2_X1 U571 ( .A1(n461), .A2(n469), .ZN(n468) );
  NAND2_X1 U572 ( .A1(n730), .A2(n467), .ZN(n466) );
  NAND2_X1 U573 ( .A1(n415), .A2(n694), .ZN(n684) );
  XNOR2_X1 U574 ( .A(n680), .B(n681), .ZN(n415) );
  XNOR2_X1 U575 ( .A(n454), .B(n386), .ZN(n453) );
  AND2_X2 U576 ( .A1(n442), .A2(n443), .ZN(n416) );
  XNOR2_X1 U577 ( .A(n511), .B(n417), .ZN(n554) );
  NAND2_X1 U578 ( .A1(n584), .A2(G221), .ZN(n417) );
  NOR2_X1 U579 ( .A1(n418), .A2(n446), .ZN(n456) );
  NAND2_X1 U580 ( .A1(n490), .A2(n678), .ZN(n510) );
  NAND2_X1 U581 ( .A1(n794), .A2(KEYINPUT83), .ZN(n420) );
  NAND2_X1 U582 ( .A1(n421), .A2(n694), .ZN(n689) );
  XNOR2_X1 U583 ( .A(n686), .B(n687), .ZN(n421) );
  INV_X1 U584 ( .A(n609), .ZN(n748) );
  NAND2_X1 U585 ( .A1(n445), .A2(KEYINPUT65), .ZN(n443) );
  XNOR2_X1 U586 ( .A(n646), .B(n385), .ZN(n455) );
  XNOR2_X1 U587 ( .A(n423), .B(n422), .ZN(n426) );
  XNOR2_X2 U588 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n422) );
  XNOR2_X1 U589 ( .A(n424), .B(G128), .ZN(n425) );
  XNOR2_X2 U590 ( .A(G119), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U591 ( .A(n426), .B(n425), .ZN(n511) );
  XNOR2_X2 U592 ( .A(n430), .B(G146), .ZN(n566) );
  AND2_X1 U593 ( .A1(n461), .A2(n431), .ZN(n724) );
  INV_X1 U594 ( .A(n735), .ZN(n431) );
  INV_X1 U595 ( .A(n461), .ZN(n432) );
  INV_X1 U596 ( .A(n371), .ZN(n434) );
  NAND2_X1 U597 ( .A1(n664), .A2(n438), .ZN(n437) );
  INV_X1 U598 ( .A(KEYINPUT36), .ZN(n439) );
  NAND2_X1 U599 ( .A1(n388), .A2(n510), .ZN(n445) );
  NAND2_X1 U600 ( .A1(n441), .A2(n378), .ZN(n440) );
  NAND2_X1 U601 ( .A1(n444), .A2(n674), .ZN(n441) );
  NAND2_X1 U602 ( .A1(n444), .A2(n387), .ZN(n442) );
  NAND2_X1 U603 ( .A1(n673), .A2(n794), .ZN(n444) );
  NAND2_X1 U604 ( .A1(n717), .A2(n663), .ZN(n446) );
  AND2_X2 U605 ( .A1(n509), .A2(n505), .ZN(n504) );
  XNOR2_X2 U606 ( .A(n558), .B(n557), .ZN(n619) );
  BUF_X1 U607 ( .A(n806), .Z(n447) );
  NOR2_X2 U608 ( .A1(n473), .A2(n472), .ZN(n471) );
  NOR2_X1 U609 ( .A1(n504), .A2(n520), .ZN(n483) );
  NOR2_X1 U610 ( .A1(n626), .A2(n656), .ZN(n627) );
  NAND2_X1 U611 ( .A1(n521), .A2(n698), .ZN(n520) );
  NOR2_X2 U612 ( .A1(n539), .A2(G902), .ZN(n540) );
  XNOR2_X1 U613 ( .A(n471), .B(n470), .ZN(n650) );
  NAND2_X1 U614 ( .A1(n449), .A2(n643), .ZN(n644) );
  XNOR2_X1 U615 ( .A(n641), .B(n642), .ZN(n449) );
  NAND2_X1 U616 ( .A1(n809), .A2(n655), .ZN(n489) );
  XNOR2_X1 U617 ( .A(n629), .B(n487), .ZN(n486) );
  NAND2_X1 U618 ( .A1(n456), .A2(n455), .ZN(n454) );
  NAND2_X1 U619 ( .A1(n672), .A2(n638), .ZN(n495) );
  XNOR2_X1 U620 ( .A(n637), .B(n636), .ZN(n672) );
  XNOR2_X2 U621 ( .A(n468), .B(KEYINPUT42), .ZN(n810) );
  NOR2_X2 U622 ( .A1(n477), .A2(n578), .ZN(n580) );
  XNOR2_X2 U623 ( .A(n572), .B(n573), .ZN(n477) );
  AND2_X1 U624 ( .A1(n409), .A2(n798), .ZN(n783) );
  INV_X1 U625 ( .A(n678), .ZN(n479) );
  XNOR2_X1 U626 ( .A(n678), .B(KEYINPUT83), .ZN(n491) );
  XNOR2_X2 U627 ( .A(n519), .B(KEYINPUT45), .ZN(n678) );
  NOR2_X1 U628 ( .A1(n652), .A2(n668), .ZN(n653) );
  NAND2_X1 U629 ( .A1(n634), .A2(n486), .ZN(n652) );
  NAND2_X1 U630 ( .A1(n483), .A2(n508), .ZN(n519) );
  NOR2_X1 U631 ( .A1(n806), .A2(KEYINPUT44), .ZN(n505) );
  NAND2_X1 U632 ( .A1(n407), .A2(G475), .ZN(n686) );
  NAND2_X1 U633 ( .A1(n657), .A2(n656), .ZN(n513) );
  XNOR2_X1 U634 ( .A(n489), .B(KEYINPUT81), .ZN(n663) );
  XNOR2_X2 U635 ( .A(n643), .B(n517), .ZN(n741) );
  XNOR2_X1 U636 ( .A(n513), .B(n512), .ZN(n659) );
  NAND2_X1 U637 ( .A1(n491), .A2(n628), .ZN(n673) );
  XNOR2_X2 U638 ( .A(n492), .B(n380), .ZN(n617) );
  NAND2_X1 U639 ( .A1(n810), .A2(n808), .ZN(n646) );
  XNOR2_X2 U640 ( .A(n497), .B(n496), .ZN(n794) );
  NAND2_X1 U641 ( .A1(n676), .A2(n718), .ZN(n497) );
  XNOR2_X2 U642 ( .A(n499), .B(n523), .ZN(n661) );
  NAND2_X1 U643 ( .A1(n690), .A2(n675), .ZN(n499) );
  NOR2_X1 U644 ( .A1(n615), .A2(n502), .ZN(n501) );
  NAND2_X1 U645 ( .A1(n645), .A2(n503), .ZN(n502) );
  AND2_X2 U646 ( .A1(n805), .A2(n803), .ZN(n509) );
  NAND2_X1 U647 ( .A1(n515), .A2(n524), .ZN(n514) );
  XNOR2_X1 U648 ( .A(n516), .B(KEYINPUT34), .ZN(n515) );
  XNOR2_X2 U649 ( .A(n518), .B(n377), .ZN(n643) );
  OR2_X2 U650 ( .A1(n768), .A2(G902), .ZN(n518) );
  NAND2_X1 U651 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U652 ( .A(n693), .B(n692), .ZN(n695) );
  XNOR2_X1 U653 ( .A(n561), .B(G146), .ZN(n542) );
  AND2_X1 U654 ( .A1(G210), .A2(n571), .ZN(n523) );
  AND2_X1 U655 ( .A1(n617), .A2(n616), .ZN(n524) );
  XOR2_X1 U656 ( .A(n793), .B(n542), .Z(n525) );
  INV_X1 U657 ( .A(KEYINPUT86), .ZN(n670) );
  XNOR2_X1 U658 ( .A(n604), .B(KEYINPUT98), .ZN(n605) );
  INV_X1 U659 ( .A(KEYINPUT65), .ZN(n679) );
  XNOR2_X1 U660 ( .A(n606), .B(n605), .ZN(n685) );
  INV_X1 U661 ( .A(KEYINPUT60), .ZN(n688) );
  XNOR2_X2 U662 ( .A(G101), .B(KEYINPUT67), .ZN(n526) );
  XNOR2_X2 U663 ( .A(n526), .B(KEYINPUT4), .ZN(n543) );
  XNOR2_X1 U664 ( .A(KEYINPUT3), .B(G119), .ZN(n780) );
  XNOR2_X1 U665 ( .A(n562), .B(G146), .ZN(n531) );
  INV_X1 U666 ( .A(n528), .ZN(n588) );
  INV_X1 U667 ( .A(n604), .ZN(n527) );
  NAND2_X1 U668 ( .A1(n588), .A2(n527), .ZN(n530) );
  NAND2_X1 U669 ( .A1(n604), .A2(n528), .ZN(n529) );
  XNOR2_X1 U670 ( .A(n531), .B(n793), .ZN(n538) );
  XOR2_X1 U671 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n533) );
  NOR2_X1 U672 ( .A1(G953), .A2(G237), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n598), .A2(G210), .ZN(n532) );
  XNOR2_X1 U674 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U675 ( .A(n534), .B(G116), .Z(n536) );
  XNOR2_X1 U676 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U677 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U678 ( .A(n541), .B(KEYINPUT76), .Z(n561) );
  XNOR2_X1 U679 ( .A(n543), .B(KEYINPUT77), .ZN(n547) );
  AND2_X1 U680 ( .A1(G227), .A2(n798), .ZN(n545) );
  XNOR2_X1 U681 ( .A(G107), .B(n551), .ZN(n548) );
  XNOR2_X1 U682 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U683 ( .A(n525), .B(n550), .ZN(n768) );
  NAND2_X1 U684 ( .A1(n478), .A2(G234), .ZN(n553) );
  XNOR2_X1 U685 ( .A(n553), .B(n552), .ZN(n584) );
  XNOR2_X1 U686 ( .A(n554), .B(n791), .ZN(n773) );
  NAND2_X1 U687 ( .A1(G234), .A2(n675), .ZN(n556) );
  XNOR2_X1 U688 ( .A(n556), .B(KEYINPUT20), .ZN(n559) );
  AND2_X1 U689 ( .A1(G217), .A2(n559), .ZN(n557) );
  NAND2_X1 U690 ( .A1(n559), .A2(G221), .ZN(n560) );
  NAND2_X1 U691 ( .A1(n452), .A2(n610), .ZN(n750) );
  XOR2_X1 U692 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n573) );
  XOR2_X1 U693 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n564) );
  NAND2_X1 U694 ( .A1(G224), .A2(n798), .ZN(n563) );
  XNOR2_X1 U695 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U696 ( .A(n565), .B(KEYINPUT89), .Z(n569) );
  XNOR2_X1 U697 ( .A(n566), .B(n567), .ZN(n568) );
  NAND2_X1 U698 ( .A1(G214), .A2(n571), .ZN(n726) );
  NAND2_X1 U699 ( .A1(n661), .A2(n726), .ZN(n572) );
  NOR2_X1 U700 ( .A1(G953), .A2(n759), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n576), .A2(n575), .ZN(n630) );
  NOR2_X1 U702 ( .A1(G898), .A2(n630), .ZN(n577) );
  NOR2_X1 U703 ( .A1(n632), .A2(n577), .ZN(n578) );
  INV_X1 U704 ( .A(KEYINPUT0), .ZN(n579) );
  NOR2_X1 U705 ( .A1(n750), .A2(n615), .ZN(n581) );
  XNOR2_X1 U706 ( .A(n581), .B(KEYINPUT31), .ZN(n713) );
  NAND2_X1 U707 ( .A1(n713), .A2(n700), .ZN(n607) );
  NAND2_X1 U708 ( .A1(n584), .A2(G217), .ZN(n592) );
  XNOR2_X1 U709 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U710 ( .A(n587), .B(KEYINPUT7), .Z(n591) );
  XNOR2_X1 U711 ( .A(n588), .B(n589), .ZN(n590) );
  NOR2_X1 U712 ( .A1(G902), .A2(n771), .ZN(n593) );
  XNOR2_X1 U713 ( .A(n595), .B(n594), .ZN(n596) );
  NAND2_X1 U714 ( .A1(G214), .A2(n598), .ZN(n600) );
  XNOR2_X1 U715 ( .A(n405), .B(G143), .ZN(n603) );
  NOR2_X1 U716 ( .A1(n617), .A2(n613), .ZN(n704) );
  INV_X1 U717 ( .A(n704), .ZN(n714) );
  NAND2_X1 U718 ( .A1(n658), .A2(n714), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n607), .A2(n648), .ZN(n608) );
  XNOR2_X1 U720 ( .A(n608), .B(KEYINPUT101), .ZN(n624) );
  NAND2_X1 U721 ( .A1(n610), .A2(n656), .ZN(n612) );
  INV_X1 U722 ( .A(n613), .ZN(n616) );
  XNOR2_X1 U723 ( .A(KEYINPUT78), .B(KEYINPUT85), .ZN(n614) );
  INV_X1 U724 ( .A(n741), .ZN(n666) );
  OR2_X1 U725 ( .A1(n358), .A2(n656), .ZN(n620) );
  NOR2_X1 U726 ( .A1(n741), .A2(n620), .ZN(n621) );
  XNOR2_X1 U727 ( .A(n621), .B(KEYINPUT79), .ZN(n622) );
  OR2_X1 U728 ( .A1(n666), .A2(n625), .ZN(n626) );
  NAND2_X1 U729 ( .A1(n627), .A2(n358), .ZN(n698) );
  INV_X1 U730 ( .A(n675), .ZN(n628) );
  NAND2_X1 U731 ( .A1(n748), .A2(n726), .ZN(n629) );
  XOR2_X1 U732 ( .A(n630), .B(KEYINPUT105), .Z(n631) );
  NOR2_X1 U733 ( .A1(G900), .A2(n631), .ZN(n633) );
  NOR2_X1 U734 ( .A1(n633), .A2(n632), .ZN(n640) );
  INV_X1 U735 ( .A(n727), .ZN(n635) );
  NOR2_X2 U736 ( .A1(n652), .A2(n635), .ZN(n637) );
  INV_X1 U737 ( .A(n658), .ZN(n638) );
  XNOR2_X1 U738 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n642) );
  NAND2_X1 U739 ( .A1(n657), .A2(n748), .ZN(n641) );
  INV_X1 U740 ( .A(n645), .ZN(n729) );
  INV_X1 U741 ( .A(n648), .ZN(n731) );
  NAND2_X1 U742 ( .A1(n731), .A2(n708), .ZN(n649) );
  NAND2_X1 U743 ( .A1(KEYINPUT47), .A2(n731), .ZN(n651) );
  XNOR2_X1 U744 ( .A(KEYINPUT82), .B(n651), .ZN(n655) );
  INV_X1 U745 ( .A(n373), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n653), .A2(n524), .ZN(n654) );
  INV_X1 U747 ( .A(n711), .ZN(n709) );
  AND2_X1 U748 ( .A1(n726), .A2(n373), .ZN(n662) );
  NAND2_X1 U749 ( .A1(n371), .A2(n726), .ZN(n665) );
  NOR2_X1 U750 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U751 ( .A(KEYINPUT43), .B(n667), .Z(n669) );
  NAND2_X1 U752 ( .A1(n669), .A2(n668), .ZN(n719) );
  NAND2_X1 U753 ( .A1(n372), .A2(n704), .ZN(n718) );
  INV_X1 U754 ( .A(KEYINPUT2), .ZN(n674) );
  NAND2_X1 U755 ( .A1(KEYINPUT2), .A2(n718), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n407), .A2(G472), .ZN(n680) );
  NOR2_X1 U757 ( .A1(G952), .A2(n798), .ZN(n682) );
  INV_X1 U758 ( .A(n778), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT63), .B(KEYINPUT111), .Z(n683) );
  XNOR2_X1 U760 ( .A(n684), .B(n683), .ZN(G57) );
  XNOR2_X1 U761 ( .A(n689), .B(n688), .ZN(G60) );
  NAND2_X1 U762 ( .A1(n769), .A2(G210), .ZN(n693) );
  XOR2_X1 U763 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n691) );
  XNOR2_X1 U764 ( .A(n362), .B(n691), .ZN(n692) );
  INV_X1 U765 ( .A(KEYINPUT56), .ZN(n696) );
  XNOR2_X1 U766 ( .A(n697), .B(n696), .ZN(G51) );
  XNOR2_X1 U767 ( .A(G101), .B(n698), .ZN(G3) );
  NOR2_X1 U768 ( .A1(n711), .A2(n700), .ZN(n699) );
  XOR2_X1 U769 ( .A(G104), .B(n699), .Z(G6) );
  NOR2_X1 U770 ( .A1(n700), .A2(n714), .ZN(n702) );
  XNOR2_X1 U771 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n701) );
  XNOR2_X1 U772 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U773 ( .A(G107), .B(n703), .ZN(G9) );
  XOR2_X1 U774 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U775 ( .A1(n708), .A2(n704), .ZN(n705) );
  XNOR2_X1 U776 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U777 ( .A(G128), .B(n707), .ZN(G30) );
  NAND2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U779 ( .A(n710), .B(G146), .ZN(G48) );
  NOR2_X1 U780 ( .A1(n711), .A2(n713), .ZN(n712) );
  XOR2_X1 U781 ( .A(G113), .B(n712), .Z(G15) );
  NOR2_X1 U782 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U783 ( .A(G116), .B(n715), .Z(G18) );
  XOR2_X1 U784 ( .A(G125), .B(KEYINPUT37), .Z(n716) );
  XNOR2_X1 U785 ( .A(n361), .B(n716), .ZN(G27) );
  XNOR2_X1 U786 ( .A(G134), .B(n718), .ZN(G36) );
  XNOR2_X1 U787 ( .A(G140), .B(n719), .ZN(G42) );
  INV_X1 U788 ( .A(n794), .ZN(n720) );
  NOR2_X1 U789 ( .A1(KEYINPUT2), .A2(n721), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n725) );
  NOR2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n762) );
  NOR2_X1 U792 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n734) );
  NOR2_X1 U794 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U795 ( .A(n732), .B(KEYINPUT116), .ZN(n733) );
  NOR2_X1 U796 ( .A1(n734), .A2(n733), .ZN(n736) );
  NOR2_X1 U797 ( .A1(n736), .A2(n735), .ZN(n755) );
  NAND2_X1 U798 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U799 ( .A(n739), .B(KEYINPUT49), .ZN(n740) );
  XNOR2_X1 U800 ( .A(KEYINPUT113), .B(n740), .ZN(n746) );
  NAND2_X1 U801 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U802 ( .A(n743), .B(KEYINPUT114), .ZN(n744) );
  XNOR2_X1 U803 ( .A(KEYINPUT50), .B(n744), .ZN(n745) );
  NAND2_X1 U804 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U805 ( .A1(n452), .A2(n747), .ZN(n749) );
  XNOR2_X1 U806 ( .A(n749), .B(KEYINPUT115), .ZN(n751) );
  NAND2_X1 U807 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U808 ( .A(KEYINPUT51), .B(n752), .ZN(n753) );
  NOR2_X1 U809 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U810 ( .A(n756), .B(KEYINPUT117), .Z(n757) );
  XNOR2_X1 U811 ( .A(KEYINPUT52), .B(n757), .ZN(n758) );
  NOR2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U813 ( .A1(G953), .A2(n760), .ZN(n761) );
  NAND2_X1 U814 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U815 ( .A(KEYINPUT118), .B(n763), .ZN(n764) );
  XOR2_X1 U816 ( .A(KEYINPUT53), .B(n764), .Z(G75) );
  XOR2_X1 U817 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n766) );
  XNOR2_X1 U818 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n765) );
  XNOR2_X1 U819 ( .A(n766), .B(n765), .ZN(n767) );
  BUF_X2 U820 ( .A(n769), .Z(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(G469), .ZN(n770) );
  NAND2_X1 U822 ( .A1(n774), .A2(G478), .ZN(n772) );
  XNOR2_X1 U823 ( .A(n370), .B(KEYINPUT122), .ZN(n776) );
  NAND2_X1 U824 ( .A1(G217), .A2(n774), .ZN(n775) );
  XNOR2_X1 U825 ( .A(n775), .B(n776), .ZN(n777) );
  NOR2_X1 U826 ( .A1(n778), .A2(n777), .ZN(G66) );
  XNOR2_X1 U827 ( .A(n780), .B(n779), .ZN(n782) );
  NOR2_X1 U828 ( .A1(G898), .A2(n798), .ZN(n781) );
  NOR2_X1 U829 ( .A1(n782), .A2(n781), .ZN(n790) );
  XNOR2_X1 U830 ( .A(KEYINPUT123), .B(n783), .ZN(n787) );
  NAND2_X1 U831 ( .A1(G953), .A2(G224), .ZN(n784) );
  XNOR2_X1 U832 ( .A(KEYINPUT61), .B(n784), .ZN(n785) );
  NAND2_X1 U833 ( .A1(n785), .A2(G898), .ZN(n786) );
  NAND2_X1 U834 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U835 ( .A(n788), .B(KEYINPUT124), .ZN(n789) );
  XNOR2_X1 U836 ( .A(n790), .B(n789), .ZN(G69) );
  XNOR2_X1 U837 ( .A(n791), .B(KEYINPUT4), .ZN(n792) );
  XOR2_X1 U838 ( .A(n793), .B(n792), .Z(n796) );
  XOR2_X1 U839 ( .A(n796), .B(n365), .Z(n795) );
  NAND2_X1 U840 ( .A1(n795), .A2(n798), .ZN(n801) );
  XNOR2_X1 U841 ( .A(n796), .B(G227), .ZN(n797) );
  NOR2_X1 U842 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U843 ( .A1(G900), .A2(n799), .ZN(n800) );
  NAND2_X1 U844 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U845 ( .A(KEYINPUT125), .B(n802), .ZN(G72) );
  XNOR2_X1 U846 ( .A(n803), .B(G122), .ZN(n804) );
  XNOR2_X1 U847 ( .A(n804), .B(KEYINPUT126), .ZN(G24) );
  XNOR2_X1 U848 ( .A(n408), .B(G110), .ZN(G12) );
  XNOR2_X1 U849 ( .A(G119), .B(KEYINPUT127), .ZN(n807) );
  XNOR2_X1 U850 ( .A(n807), .B(n447), .ZN(G21) );
  XNOR2_X1 U851 ( .A(n406), .B(G131), .ZN(G33) );
  XNOR2_X1 U852 ( .A(n374), .B(G143), .ZN(G45) );
  XNOR2_X1 U853 ( .A(n810), .B(G137), .ZN(G39) );
endmodule

