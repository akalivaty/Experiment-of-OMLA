//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n193), .A3(new_n197), .A4(new_n191), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(KEYINPUT65), .A3(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT80), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G104), .ZN(new_n206));
  AOI21_X1  g020(.A(G107), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT3), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n205), .A2(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(KEYINPUT80), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT3), .A2(G107), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(G104), .B2(new_n212), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n208), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n216), .A2(KEYINPUT81), .A3(new_n218), .A4(new_n208), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n211), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n226), .A3(G143), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n228), .B(G146), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n223), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n233), .ZN(new_n235));
  AOI211_X1 g049(.A(new_n235), .B(new_n211), .C1(new_n221), .C2(new_n222), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n202), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(KEYINPUT12), .B(new_n202), .C1(new_n234), .C2(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n211), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n212), .B1(new_n204), .B2(new_n206), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n209), .A3(G104), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT3), .A2(G107), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT81), .B1(new_n248), .B2(new_n208), .ZN(new_n249));
  NOR4_X1   g063(.A1(new_n243), .A2(new_n247), .A3(new_n220), .A4(G101), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n233), .B(new_n242), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT10), .B1(new_n223), .B2(new_n233), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n216), .A2(new_n218), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G101), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n221), .A2(new_n222), .ZN(new_n261));
  OAI21_X1  g075(.A(G101), .B1(new_n243), .B2(new_n247), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n260), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n227), .A2(new_n229), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT0), .B(G128), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n256), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n263), .B1(new_n221), .B2(new_n222), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n269), .A2(new_n272), .ZN(new_n276));
  NOR4_X1   g090(.A1(new_n275), .A2(KEYINPUT82), .A3(new_n260), .A4(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n255), .B(new_n201), .C1(new_n274), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n241), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT78), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G227), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G953), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT77), .B(G110), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n285), .A2(KEYINPUT79), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(KEYINPUT79), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n251), .A2(new_n252), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n233), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n261), .A2(new_n264), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n273), .A3(new_n259), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT82), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n265), .A2(new_n256), .A3(new_n273), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n289), .B1(new_n297), .B2(new_n201), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n274), .A2(new_n277), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n202), .B1(new_n299), .B2(new_n292), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n288), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G469), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n187), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n278), .A2(KEYINPUT84), .A3(new_n285), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT84), .B1(new_n278), .B2(new_n285), .ZN(new_n307));
  INV_X1    g121(.A(new_n241), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n285), .B1(new_n300), .B2(new_n278), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n303), .B(new_n305), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n241), .A2(new_n278), .B1(KEYINPUT79), .B2(new_n285), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n312), .A2(new_n286), .B1(new_n300), .B2(new_n298), .ZN(new_n313));
  OAI211_X1 g127(.A(KEYINPUT83), .B(G469), .C1(new_n313), .C2(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n304), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n316));
  XNOR2_X1  g130(.A(G113), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n203), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT90), .A3(G146), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT90), .B1(new_n323), .B2(new_n226), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n226), .B2(new_n323), .ZN(new_n327));
  NOR2_X1   g141(.A1(G237), .A2(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G214), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n228), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n328), .B(G214), .C1(KEYINPUT89), .C2(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT18), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n333), .A2(new_n334), .A3(new_n197), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n331), .A2(new_n332), .B1(KEYINPUT18), .B2(G131), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n325), .B(new_n327), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(G131), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT17), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n331), .A2(new_n197), .A3(new_n332), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT92), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(KEYINPUT17), .A3(G131), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n338), .A2(new_n344), .A3(new_n339), .A4(new_n340), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT16), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n350), .A2(new_n319), .A3(KEYINPUT72), .A4(G125), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n226), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n349), .A3(G146), .A4(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT91), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(KEYINPUT91), .A3(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n318), .B(new_n337), .C1(new_n346), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n338), .A2(new_n340), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n323), .B(KEYINPUT19), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(G146), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n354), .B(KEYINPUT73), .Z(new_n365));
  OAI21_X1  g179(.A(new_n337), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n318), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G475), .A2(G902), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT93), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n316), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI211_X1 g188(.A(KEYINPUT20), .B(new_n371), .C1(new_n360), .C2(new_n368), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n337), .B1(new_n346), .B2(new_n359), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n367), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n379), .B2(new_n360), .ZN(new_n380));
  INV_X1    g194(.A(G475), .ZN(new_n381));
  OR2_X1    g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT94), .ZN(new_n383));
  OAI22_X1  g197(.A1(new_n373), .A2(new_n375), .B1(new_n380), .B2(new_n381), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT9), .B(G234), .Z(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n389), .A2(new_n390), .A3(G953), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G116), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n228), .A2(G128), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT95), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n224), .A2(G143), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n228), .A2(KEYINPUT13), .A3(G128), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT95), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n395), .A2(new_n401), .A3(new_n396), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n394), .B1(G134), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n399), .A2(new_n395), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n189), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n405), .B(new_n189), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n393), .A2(new_n209), .ZN(new_n410));
  INV_X1    g224(.A(G116), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT14), .A3(G122), .ZN(new_n412));
  INV_X1    g226(.A(new_n393), .ZN(new_n413));
  OAI211_X1 g227(.A(G107), .B(new_n412), .C1(new_n413), .C2(KEYINPUT14), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n392), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n415), .A3(new_n391), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(KEYINPUT96), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT96), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n392), .C1(new_n408), .C2(new_n416), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n305), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n422), .B(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n387), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G214), .B1(G237), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(G953), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G952), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(G234), .B2(G237), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT21), .B(G898), .Z(new_n432));
  NAND2_X1  g246(.A1(G234), .A2(G237), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(G902), .A3(G953), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G119), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT67), .B1(new_n436), .B2(G116), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT67), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n411), .A3(G119), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n437), .A2(new_n439), .B1(G116), .B2(new_n436), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT66), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT2), .B(G113), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n440), .B2(new_n441), .ZN(new_n446));
  INV_X1    g260(.A(new_n262), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n444), .A2(new_n446), .B1(new_n447), .B2(new_n258), .ZN(new_n448));
  INV_X1    g262(.A(G113), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n440), .B2(KEYINPUT5), .ZN(new_n450));
  OR3_X1    g264(.A1(new_n411), .A2(KEYINPUT5), .A3(G119), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n450), .A2(new_n451), .B1(new_n440), .B2(new_n445), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n293), .A2(new_n448), .B1(new_n223), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G122), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT85), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n456), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(KEYINPUT6), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n233), .A2(new_n321), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n276), .B2(new_n321), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT88), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n428), .A2(G224), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n463), .B(KEYINPUT87), .Z(new_n464));
  XNOR2_X1  g278(.A(new_n462), .B(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n453), .A2(new_n456), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR4_X1   g283(.A1(new_n453), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n456), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n459), .B(new_n465), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G210), .B1(G237), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n464), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n461), .B(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n223), .B(new_n452), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n455), .B(KEYINPUT8), .Z(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n478), .B2(new_n458), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n471), .A2(new_n472), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n472), .B1(new_n471), .B2(new_n479), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n427), .B(new_n435), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n315), .A2(new_n426), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n436), .B2(G128), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n488), .B(new_n489), .C1(G119), .C2(new_n224), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G110), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  XOR2_X1   g306(.A(G119), .B(G128), .Z(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n355), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n354), .B(KEYINPUT73), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n490), .A2(G110), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n494), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n497), .A2(new_n498), .B1(new_n226), .B2(new_n323), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(G137), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n428), .A2(G221), .A3(G234), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n495), .A2(new_n500), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n504), .B(KEYINPUT75), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n305), .B(new_n505), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n510), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(KEYINPUT76), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT76), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n514), .A3(new_n510), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n390), .B1(G234), .B2(new_n305), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n507), .A2(new_n508), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n507), .B2(new_n504), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n516), .A2(G902), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n513), .A2(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT32), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n444), .A2(new_n446), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n199), .A2(new_n200), .A3(new_n273), .ZN(new_n526));
  INV_X1    g340(.A(new_n191), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n189), .A2(G137), .ZN(new_n528));
  OAI21_X1  g342(.A(G131), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n233), .A2(new_n198), .A3(new_n529), .ZN(new_n530));
  AOI211_X1 g344(.A(KEYINPUT68), .B(new_n525), .C1(new_n526), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(KEYINPUT68), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT30), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n526), .A2(new_n532), .A3(new_n530), .A4(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n524), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n526), .A2(new_n446), .A3(new_n444), .A4(new_n530), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(G101), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n328), .A2(G210), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n537), .A2(new_n538), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n537), .A2(new_n546), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT31), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT28), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n526), .A2(new_n530), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n524), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n554), .B2(new_n539), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n539), .A2(new_n552), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n545), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n537), .A2(KEYINPUT69), .A3(new_n538), .A4(new_n546), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n549), .A2(new_n551), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n560), .A2(KEYINPUT70), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT70), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n523), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n555), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n565), .A2(KEYINPUT29), .A3(new_n544), .A4(new_n556), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n544), .A3(new_n556), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT29), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n553), .A2(new_n533), .A3(KEYINPUT30), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n535), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n540), .B1(new_n571), .B2(new_n524), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n544), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n305), .B(new_n566), .C1(new_n569), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n522), .B1(new_n564), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n486), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G101), .ZN(G3));
  NAND2_X1  g394(.A1(new_n315), .A2(new_n484), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n560), .A2(new_n305), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G472), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n521), .B(new_n583), .C1(new_n563), .C2(new_n562), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n422), .A2(new_n423), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n419), .A2(new_n587), .A3(new_n421), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n417), .A2(KEYINPUT33), .A3(new_n418), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n588), .A2(G478), .A3(new_n305), .A4(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n383), .A2(new_n386), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n483), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT34), .B(G104), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  OR3_X1    g409(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT97), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT97), .B1(new_n373), .B2(new_n375), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n596), .A2(new_n597), .A3(new_n382), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n425), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n482), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n585), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  OAI21_X1  g417(.A(new_n583), .B1(new_n562), .B2(new_n563), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n508), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n508), .A2(new_n605), .A3(new_n606), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n507), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n609), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n611), .A2(new_n506), .A3(new_n607), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n517), .A2(new_n513), .B1(new_n613), .B2(new_n520), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n604), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n485), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT37), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G110), .ZN(G12));
  AOI21_X1  g432(.A(new_n614), .B1(new_n564), .B2(new_n577), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n427), .B1(new_n480), .B2(new_n481), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n619), .A2(new_n621), .A3(new_n484), .A4(new_n315), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n434), .A2(G900), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n431), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n599), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n224), .ZN(G30));
  INV_X1    g443(.A(new_n427), .ZN(new_n630));
  INV_X1    g444(.A(new_n581), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n624), .B(KEYINPUT39), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n630), .B1(new_n633), .B2(KEYINPUT40), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n572), .A2(new_n545), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n554), .A2(new_n539), .A3(new_n545), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n305), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n564), .A2(new_n576), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n634), .A2(new_n614), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n480), .A2(new_n481), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT38), .Z(new_n642));
  AOI21_X1  g456(.A(KEYINPUT94), .B1(new_n377), .B2(new_n382), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n384), .A2(new_n385), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n425), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n642), .B(new_n646), .C1(new_n633), .C2(KEYINPUT40), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n228), .ZN(G45));
  NAND2_X1  g463(.A1(new_n591), .A2(new_n624), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n622), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n226), .ZN(G48));
  OAI21_X1  g466(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G469), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n484), .A3(new_n311), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n654), .A2(KEYINPUT99), .A3(new_n484), .A4(new_n311), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n592), .A3(new_n578), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT41), .B(G113), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G15));
  NAND4_X1  g475(.A1(new_n657), .A2(new_n578), .A3(new_n600), .A4(new_n658), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G116), .ZN(G18));
  NAND4_X1  g477(.A1(new_n657), .A2(new_n621), .A3(new_n435), .A4(new_n658), .ZN(new_n664));
  INV_X1    g478(.A(new_n426), .ZN(new_n665));
  INV_X1    g479(.A(new_n619), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n436), .ZN(G21));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n645), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n387), .A2(KEYINPUT102), .A3(new_n425), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n560), .A2(new_n561), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT100), .B1(new_n582), .B2(G472), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  INV_X1    g489(.A(G472), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n675), .B(new_n676), .C1(new_n560), .C2(new_n305), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n521), .B(new_n673), .C1(new_n674), .C2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n672), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(new_n664), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  AND2_X1   g498(.A1(new_n591), .A2(new_n624), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n657), .A2(new_n621), .A3(new_n685), .A4(new_n658), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n674), .A2(new_n677), .ZN(new_n687));
  INV_X1    g501(.A(new_n673), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n614), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n321), .ZN(G27));
  INV_X1    g507(.A(new_n484), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n313), .B2(G902), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n694), .B1(new_n311), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n480), .A2(new_n481), .A3(new_n630), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n673), .A2(new_n523), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n522), .B1(new_n577), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n699), .A2(new_n701), .A3(KEYINPUT42), .A4(new_n685), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n564), .A2(new_n577), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n521), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n704), .A2(new_n698), .A3(new_n650), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n702), .B1(new_n705), .B2(KEYINPUT42), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G131), .ZN(G33));
  NAND3_X1  g521(.A1(new_n699), .A2(new_n578), .A3(new_n626), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  AOI21_X1  g523(.A(new_n387), .B1(new_n586), .B2(new_n590), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT43), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n590), .A2(new_n586), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n590), .A2(KEYINPUT104), .A3(new_n586), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n383), .A2(new_n714), .A3(new_n386), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n717), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n711), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n604), .B(new_n690), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n726));
  OR3_X1    g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n288), .A2(new_n301), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT103), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n303), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n313), .A2(new_n732), .A3(KEYINPUT45), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(G469), .A2(G902), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n735), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n311), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n484), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n632), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n726), .B1(new_n724), .B2(new_n725), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n727), .A2(new_n697), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  NAND2_X1  g560(.A1(new_n742), .A2(KEYINPUT47), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n703), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n522), .A3(new_n685), .A4(new_n697), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G140), .ZN(G42));
  AND2_X1   g566(.A1(new_n657), .A2(new_n658), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n430), .A2(new_n753), .A3(new_n697), .A4(new_n722), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n701), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n639), .A2(new_n431), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n521), .A2(new_n753), .A3(new_n697), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n429), .B1(new_n760), .B2(new_n591), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n678), .B(new_n679), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n762), .A2(new_n430), .A3(new_n722), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n621), .A3(new_n753), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n758), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n763), .A2(new_n697), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n747), .A2(new_n749), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n654), .A2(new_n311), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n484), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT115), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n766), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n722), .A2(new_n430), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n642), .A2(new_n427), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n753), .A3(new_n762), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n763), .A2(KEYINPUT50), .A3(new_n753), .A4(new_n773), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n387), .A2(new_n712), .ZN(new_n779));
  INV_X1    g593(.A(new_n691), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n760), .A2(new_n779), .B1(new_n754), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n771), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n757), .B(new_n765), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n778), .A2(new_n786), .A3(new_n781), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n786), .B1(new_n778), .B2(new_n781), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT51), .B(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n784), .A2(KEYINPUT117), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT117), .B1(new_n784), .B2(new_n789), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n584), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n383), .A2(new_n425), .A3(new_n386), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(new_n591), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n631), .A2(new_n483), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n579), .A2(new_n616), .A3(new_n796), .A4(KEYINPUT107), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT107), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n485), .B1(new_n704), .B2(new_n615), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n483), .B1(new_n794), .B2(new_n591), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n581), .A3(new_n584), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n798), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n657), .A2(new_n621), .A3(new_n658), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n435), .A3(new_n426), .A4(new_n619), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n659), .A2(new_n662), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n683), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n315), .A2(new_n621), .A3(new_n484), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n809), .B(new_n619), .C1(new_n626), .C2(new_n685), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n620), .B1(new_n670), .B2(new_n671), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n694), .B(new_n625), .C1(new_n311), .C2(new_n695), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n614), .A3(new_n639), .A4(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n810), .B(new_n813), .C1(new_n691), .C2(new_n686), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n689), .A2(new_n685), .A3(new_n697), .A4(new_n696), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT108), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n697), .A2(new_n598), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n425), .A2(new_n625), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n697), .A2(new_n598), .A3(new_n818), .A4(new_n820), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n703), .A3(new_n484), .A4(new_n315), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n817), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n690), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n825), .A2(new_n706), .A3(new_n708), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n808), .A2(new_n816), .A3(KEYINPUT53), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT111), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT109), .B1(new_n814), .B2(new_n815), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n815), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n622), .B1(new_n627), .B2(new_n650), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n692), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT109), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT52), .A4(new_n813), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n814), .A2(KEYINPUT110), .A3(new_n815), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n830), .A2(new_n833), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n659), .B(new_n662), .C1(new_n682), .C2(new_n664), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n667), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n797), .A2(new_n802), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n826), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n829), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n827), .A2(KEYINPUT111), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n828), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n814), .B(KEYINPUT52), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n829), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n825), .A2(new_n706), .A3(KEYINPUT53), .A4(new_n708), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n803), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n840), .B2(new_n667), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n683), .A2(new_n805), .A3(KEYINPUT112), .A4(new_n806), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n848), .B1(new_n839), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n846), .A2(KEYINPUT54), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(G952), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n792), .A2(new_n860), .B1(new_n861), .B2(new_n428), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n710), .A2(new_n427), .A3(new_n484), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n642), .A2(new_n863), .A3(new_n639), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n768), .B(KEYINPUT49), .Z(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n521), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT118), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n784), .A2(new_n789), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n784), .A2(KEYINPUT117), .A3(new_n789), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n860), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n861), .A2(new_n428), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n866), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n868), .A2(new_n877), .ZN(G75));
  NOR2_X1   g692(.A1(new_n428), .A2(G952), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(new_n465), .Z(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n856), .A2(G210), .A3(G902), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n884), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n882), .B1(new_n884), .B2(KEYINPUT119), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT120), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n879), .B(new_n886), .C1(new_n892), .C2(new_n894), .ZN(G51));
  NAND2_X1  g709(.A1(new_n856), .A2(new_n858), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n833), .A2(new_n837), .A3(new_n830), .A4(new_n838), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n854), .A3(new_n850), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n848), .A3(new_n859), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n857), .A2(KEYINPUT121), .A3(new_n859), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n735), .B(KEYINPUT57), .Z(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n309), .A2(new_n310), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT122), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n857), .A2(new_n305), .A3(new_n734), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n879), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n856), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  INV_X1    g725(.A(new_n369), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n879), .ZN(G60));
  NAND2_X1  g729(.A1(new_n901), .A2(new_n902), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n588), .A2(new_n589), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT59), .Z(new_n919));
  NOR3_X1   g733(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n860), .A2(new_n919), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n879), .B(new_n920), .C1(new_n921), .C2(new_n917), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n857), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n613), .ZN(new_n926));
  INV_X1    g740(.A(new_n879), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n519), .B(KEYINPUT123), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n857), .B2(new_n924), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g745(.A1(new_n432), .A2(G224), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G953), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT124), .B(new_n933), .C1(new_n808), .C2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(KEYINPUT124), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n880), .B1(G898), .B2(new_n428), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT125), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  XNOR2_X1  g752(.A(new_n571), .B(new_n363), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n751), .A2(new_n745), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n835), .B1(new_n640), .B2(new_n647), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT62), .Z(new_n943));
  INV_X1    g757(.A(new_n633), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n578), .A3(new_n697), .A4(new_n795), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n940), .B1(new_n946), .B2(new_n428), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n706), .A2(new_n708), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n743), .A2(new_n701), .A3(new_n811), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n941), .A2(new_n948), .A3(new_n835), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n428), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(G900), .B2(new_n428), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n952), .B2(new_n940), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n428), .B1(G227), .B2(G900), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT126), .Z(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G72));
  INV_X1    g770(.A(new_n808), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n572), .A2(new_n545), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n941), .A2(new_n943), .A3(new_n808), .A4(new_n945), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n960), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n965), .A2(KEYINPUT127), .A3(new_n635), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT127), .B1(new_n965), .B2(new_n635), .ZN(new_n967));
  OAI221_X1 g781(.A(new_n927), .B1(new_n962), .B2(new_n963), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n846), .B(new_n960), .C1(new_n545), .C2(new_n572), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n968), .B1(new_n963), .B2(new_n970), .ZN(G57));
endmodule


