

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(KEYINPUT66), .B(n541), .ZN(n794) );
  XOR2_X1 U553 ( .A(n644), .B(KEYINPUT29), .Z(n517) );
  NAND2_X1 U554 ( .A1(n679), .A2(n678), .ZN(n723) );
  AND2_X2 U555 ( .A1(n533), .A2(n532), .ZN(G160) );
  BUF_X1 U556 ( .A(n612), .Z(n540) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n660) );
  XNOR2_X1 U558 ( .A(n659), .B(KEYINPUT102), .ZN(n673) );
  AND2_X1 U559 ( .A1(n648), .A2(G1996), .ZN(n594) );
  INV_X1 U560 ( .A(KEYINPUT99), .ZN(n622) );
  XNOR2_X1 U561 ( .A(n661), .B(n660), .ZN(n669) );
  OR2_X1 U562 ( .A1(n649), .A2(n648), .ZN(n732) );
  AND2_X1 U563 ( .A1(n530), .A2(n518), .ZN(n533) );
  AND2_X2 U564 ( .A1(n592), .A2(n714), .ZN(n648) );
  AND2_X1 U565 ( .A1(n529), .A2(n528), .ZN(n518) );
  XNOR2_X1 U566 ( .A(KEYINPUT31), .B(n657), .ZN(n519) );
  XOR2_X1 U567 ( .A(n680), .B(n723), .Z(n520) );
  XNOR2_X1 U568 ( .A(n591), .B(KEYINPUT64), .ZN(n714) );
  AND2_X2 U569 ( .A1(n526), .A2(G2105), .ZN(n885) );
  NOR2_X1 U570 ( .A1(G2105), .A2(n526), .ZN(n694) );
  OR2_X1 U571 ( .A1(G301), .A2(n654), .ZN(n521) );
  XOR2_X1 U572 ( .A(KEYINPUT79), .B(n600), .Z(n522) );
  INV_X1 U573 ( .A(KEYINPUT100), .ZN(n625) );
  NOR2_X1 U574 ( .A1(n652), .A2(G168), .ZN(n653) );
  NAND2_X1 U575 ( .A1(n517), .A2(n521), .ZN(n658) );
  NAND2_X1 U576 ( .A1(n658), .A2(n519), .ZN(n659) );
  XNOR2_X1 U577 ( .A(n671), .B(KEYINPUT32), .ZN(n679) );
  INV_X1 U578 ( .A(n975), .ZN(n684) );
  AND2_X1 U579 ( .A1(n685), .A2(n684), .ZN(n686) );
  BUF_X1 U580 ( .A(n694), .Z(n890) );
  XNOR2_X1 U581 ( .A(n523), .B(KEYINPUT69), .ZN(n524) );
  XNOR2_X1 U582 ( .A(G2104), .B(KEYINPUT67), .ZN(n526) );
  NAND2_X1 U583 ( .A1(G101), .A2(n694), .ZN(n523) );
  XNOR2_X1 U584 ( .A(n524), .B(KEYINPUT23), .ZN(n530) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U586 ( .A1(G113), .A2(n886), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(KEYINPUT70), .ZN(n529) );
  NAND2_X1 U588 ( .A1(G125), .A2(n885), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT68), .ZN(n528) );
  NOR2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  XOR2_X1 U591 ( .A(KEYINPUT17), .B(n531), .Z(n549) );
  BUF_X1 U592 ( .A(n549), .Z(n889) );
  NAND2_X1 U593 ( .A1(G137), .A2(n889), .ZN(n532) );
  NOR2_X2 U594 ( .A1(G543), .A2(G651), .ZN(n798) );
  NAND2_X1 U595 ( .A1(n798), .A2(G89), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT4), .ZN(n536) );
  XOR2_X2 U597 ( .A(G543), .B(KEYINPUT0), .Z(n570) );
  XNOR2_X1 U598 ( .A(KEYINPUT71), .B(G651), .ZN(n538) );
  NOR2_X4 U599 ( .A1(n570), .A2(n538), .ZN(n797) );
  NAND2_X1 U600 ( .A1(G76), .A2(n797), .ZN(n535) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT5), .ZN(n546) );
  NOR2_X1 U603 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT1), .B(n539), .Z(n612) );
  NAND2_X1 U605 ( .A1(n540), .A2(G63), .ZN(n543) );
  NOR2_X1 U606 ( .A1(G651), .A2(n570), .ZN(n541) );
  NAND2_X1 U607 ( .A1(G51), .A2(n794), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n544), .Z(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U612 ( .A1(n885), .A2(G126), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(KEYINPUT90), .ZN(n551) );
  NAND2_X1 U614 ( .A1(G138), .A2(n549), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G114), .A2(n886), .ZN(n553) );
  NAND2_X1 U617 ( .A1(G102), .A2(n694), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X2 U619 ( .A1(n555), .A2(n554), .ZN(G164) );
  NAND2_X1 U620 ( .A1(n540), .A2(G64), .ZN(n557) );
  NAND2_X1 U621 ( .A1(G52), .A2(n794), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G77), .A2(n797), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G90), .A2(n798), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(G171) );
  INV_X1 U628 ( .A(G171), .ZN(G301) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G75), .A2(n797), .ZN(n564) );
  NAND2_X1 U631 ( .A1(G88), .A2(n798), .ZN(n563) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n540), .A2(G62), .ZN(n566) );
  NAND2_X1 U634 ( .A1(G50), .A2(n794), .ZN(n565) );
  NAND2_X1 U635 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(G166) );
  INV_X1 U637 ( .A(G166), .ZN(G303) );
  NAND2_X1 U638 ( .A1(n794), .A2(G49), .ZN(n569) );
  XNOR2_X1 U639 ( .A(n569), .B(KEYINPUT86), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G87), .A2(n570), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U643 ( .A1(n540), .A2(n573), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(G288) );
  NAND2_X1 U645 ( .A1(G86), .A2(n798), .ZN(n577) );
  NAND2_X1 U646 ( .A1(G48), .A2(n794), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G73), .A2(n797), .ZN(n578) );
  XOR2_X1 U649 ( .A(KEYINPUT2), .B(n578), .Z(n579) );
  NOR2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n540), .A2(G61), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(G305) );
  NAND2_X1 U653 ( .A1(G47), .A2(n794), .ZN(n583) );
  XNOR2_X1 U654 ( .A(n583), .B(KEYINPUT72), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G60), .A2(n540), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U657 ( .A(KEYINPUT73), .B(n586), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n797), .A2(G72), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G85), .A2(n798), .ZN(n587) );
  AND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(G290) );
  INV_X1 U662 ( .A(KEYINPUT106), .ZN(n680) );
  NAND2_X1 U663 ( .A1(G160), .A2(G40), .ZN(n713) );
  INV_X1 U664 ( .A(n713), .ZN(n592) );
  NOR2_X1 U665 ( .A1(G1384), .A2(G164), .ZN(n591) );
  XNOR2_X1 U666 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n594), .B(n593), .ZN(n596) );
  INV_X1 U668 ( .A(n648), .ZN(n662) );
  NAND2_X1 U669 ( .A1(n662), .A2(G1341), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n609) );
  XOR2_X1 U671 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n598) );
  NAND2_X1 U672 ( .A1(G81), .A2(n798), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U674 ( .A(KEYINPUT77), .B(n599), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n797), .A2(G68), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n522), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT13), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G43), .A2(n794), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n612), .A2(G56), .ZN(n605) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n605), .Z(n606) );
  NOR2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X2 U683 ( .A(KEYINPUT80), .B(n608), .Z(n978) );
  NOR2_X2 U684 ( .A1(n609), .A2(n978), .ZN(n624) );
  NAND2_X1 U685 ( .A1(G79), .A2(n797), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G92), .A2(n798), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n612), .A2(G66), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G54), .A2(n794), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U692 ( .A(KEYINPUT15), .B(n617), .Z(n990) );
  NAND2_X1 U693 ( .A1(n624), .A2(n990), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n648), .A2(G1348), .ZN(n619) );
  NOR2_X1 U695 ( .A1(G2067), .A2(n662), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(n628) );
  NOR2_X1 U699 ( .A1(n990), .A2(n624), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n639) );
  NAND2_X1 U702 ( .A1(n540), .A2(G65), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G53), .A2(n794), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U705 ( .A1(G78), .A2(n797), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G91), .A2(n798), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n809) );
  NAND2_X1 U709 ( .A1(n648), .A2(G2072), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n635), .B(KEYINPUT27), .ZN(n637) );
  AND2_X1 U711 ( .A1(G1956), .A2(n662), .ZN(n636) );
  NOR2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n809), .A2(n640), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n809), .A2(n640), .ZN(n641) );
  XOR2_X1 U716 ( .A(n641), .B(KEYINPUT28), .Z(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U718 ( .A1(n648), .A2(G1961), .ZN(n647) );
  XOR2_X1 U719 ( .A(G2078), .B(KEYINPUT25), .Z(n645) );
  XNOR2_X1 U720 ( .A(KEYINPUT98), .B(n645), .ZN(n955) );
  NOR2_X1 U721 ( .A1(n662), .A2(n955), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n654) );
  INV_X1 U723 ( .A(G8), .ZN(n649) );
  NOR2_X1 U724 ( .A1(G1966), .A2(n732), .ZN(n675) );
  NOR2_X1 U725 ( .A1(G2084), .A2(n662), .ZN(n672) );
  NOR2_X1 U726 ( .A1(n675), .A2(n672), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n653), .B(KEYINPUT101), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n654), .A2(G301), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n673), .A2(G286), .ZN(n661) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XOR2_X1 U734 ( .A(KEYINPUT104), .B(n663), .Z(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(G303), .ZN(n666) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n732), .ZN(n665) );
  NOR2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U738 ( .A(KEYINPUT105), .B(n667), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n670), .A2(G8), .ZN(n671) );
  NAND2_X1 U741 ( .A1(G8), .A2(n672), .ZN(n677) );
  INV_X1 U742 ( .A(n673), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U745 ( .A1(G1971), .A2(G303), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n681), .B(KEYINPUT107), .ZN(n683) );
  INV_X1 U747 ( .A(KEYINPUT33), .ZN(n682) );
  AND2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NAND2_X1 U750 ( .A1(n520), .A2(n686), .ZN(n722) );
  INV_X1 U751 ( .A(n732), .ZN(n687) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n981) );
  AND2_X1 U753 ( .A1(n687), .A2(n981), .ZN(n688) );
  OR2_X1 U754 ( .A1(KEYINPUT33), .A2(n688), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n975), .A2(KEYINPUT33), .ZN(n689) );
  OR2_X1 U756 ( .A1(n732), .A2(n689), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n720) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n985) );
  XOR2_X1 U759 ( .A(KEYINPUT95), .B(G1991), .Z(n956) );
  INV_X1 U760 ( .A(n956), .ZN(n702) );
  NAND2_X1 U761 ( .A1(G119), .A2(n885), .ZN(n693) );
  NAND2_X1 U762 ( .A1(G107), .A2(n886), .ZN(n692) );
  NAND2_X1 U763 ( .A1(n693), .A2(n692), .ZN(n699) );
  NAND2_X1 U764 ( .A1(G131), .A2(n889), .ZN(n696) );
  NAND2_X1 U765 ( .A1(G95), .A2(n890), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U767 ( .A(KEYINPUT93), .B(n697), .Z(n698) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U769 ( .A(KEYINPUT94), .B(n700), .Z(n875) );
  INV_X1 U770 ( .A(n875), .ZN(n701) );
  NOR2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n712) );
  XOR2_X1 U772 ( .A(KEYINPUT38), .B(KEYINPUT96), .Z(n704) );
  NAND2_X1 U773 ( .A1(G105), .A2(n890), .ZN(n703) );
  XNOR2_X1 U774 ( .A(n704), .B(n703), .ZN(n708) );
  NAND2_X1 U775 ( .A1(G141), .A2(n889), .ZN(n706) );
  NAND2_X1 U776 ( .A1(G117), .A2(n886), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n885), .A2(G129), .ZN(n709) );
  NAND2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n882) );
  AND2_X1 U781 ( .A1(n882), .A2(G1996), .ZN(n711) );
  NOR2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n938) );
  NOR2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n761) );
  INV_X1 U784 ( .A(n761), .ZN(n715) );
  NOR2_X1 U785 ( .A1(n938), .A2(n715), .ZN(n753) );
  INV_X1 U786 ( .A(n753), .ZN(n718) );
  XNOR2_X1 U787 ( .A(G1986), .B(G290), .ZN(n995) );
  NAND2_X1 U788 ( .A1(n761), .A2(n995), .ZN(n716) );
  XOR2_X1 U789 ( .A(KEYINPUT91), .B(n716), .Z(n717) );
  AND2_X1 U790 ( .A1(n718), .A2(n717), .ZN(n736) );
  NAND2_X1 U791 ( .A1(n985), .A2(n736), .ZN(n719) );
  NOR2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n739) );
  XNOR2_X1 U794 ( .A(KEYINPUT106), .B(n723), .ZN(n731) );
  NOR2_X1 U795 ( .A1(G2090), .A2(G303), .ZN(n724) );
  NAND2_X1 U796 ( .A1(G8), .A2(n724), .ZN(n729) );
  NOR2_X1 U797 ( .A1(G1981), .A2(G305), .ZN(n725) );
  XOR2_X1 U798 ( .A(n725), .B(KEYINPUT24), .Z(n726) );
  NOR2_X1 U799 ( .A1(n732), .A2(n726), .ZN(n727) );
  XOR2_X1 U800 ( .A(KEYINPUT97), .B(n727), .Z(n733) );
  INV_X1 U801 ( .A(n733), .ZN(n728) );
  AND2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n735) );
  OR2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n750) );
  NAND2_X1 U808 ( .A1(n889), .A2(G140), .ZN(n740) );
  XNOR2_X1 U809 ( .A(n740), .B(KEYINPUT92), .ZN(n742) );
  NAND2_X1 U810 ( .A1(G104), .A2(n890), .ZN(n741) );
  NAND2_X1 U811 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U812 ( .A(KEYINPUT34), .B(n743), .ZN(n748) );
  NAND2_X1 U813 ( .A1(G128), .A2(n885), .ZN(n745) );
  NAND2_X1 U814 ( .A1(G116), .A2(n886), .ZN(n744) );
  NAND2_X1 U815 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U816 ( .A(KEYINPUT35), .B(n746), .Z(n747) );
  NOR2_X1 U817 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U818 ( .A(KEYINPUT36), .B(n749), .ZN(n874) );
  XNOR2_X1 U819 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NOR2_X1 U820 ( .A1(n874), .A2(n758), .ZN(n940) );
  NAND2_X1 U821 ( .A1(n761), .A2(n940), .ZN(n756) );
  NAND2_X1 U822 ( .A1(n750), .A2(n756), .ZN(n763) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n882), .ZN(n931) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U825 ( .A1(n956), .A2(n875), .ZN(n926) );
  NOR2_X1 U826 ( .A1(n751), .A2(n926), .ZN(n752) );
  NOR2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U828 ( .A1(n931), .A2(n754), .ZN(n755) );
  XNOR2_X1 U829 ( .A(KEYINPUT39), .B(n755), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n874), .A2(n758), .ZN(n941) );
  NAND2_X1 U832 ( .A1(n759), .A2(n941), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U835 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U836 ( .A(G860), .ZN(n776) );
  OR2_X1 U837 ( .A1(n776), .A2(n978), .ZN(G153) );
  INV_X1 U838 ( .A(G57), .ZN(G237) );
  INV_X1 U839 ( .A(G132), .ZN(G219) );
  INV_X1 U840 ( .A(G82), .ZN(G220) );
  INV_X1 U841 ( .A(n809), .ZN(G299) );
  NAND2_X1 U842 ( .A1(G94), .A2(G452), .ZN(n765) );
  XOR2_X1 U843 ( .A(KEYINPUT74), .B(n765), .Z(G173) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U845 ( .A(n766), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U846 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n768) );
  INV_X1 U847 ( .A(G223), .ZN(n832) );
  NAND2_X1 U848 ( .A1(G567), .A2(n832), .ZN(n767) );
  XNOR2_X1 U849 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U850 ( .A(KEYINPUT75), .B(n769), .Z(G234) );
  INV_X1 U851 ( .A(G868), .ZN(n814) );
  NOR2_X1 U852 ( .A1(n814), .A2(G171), .ZN(n770) );
  XNOR2_X1 U853 ( .A(n770), .B(KEYINPUT81), .ZN(n772) );
  OR2_X1 U854 ( .A1(G868), .A2(n990), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U856 ( .A(KEYINPUT82), .B(n773), .ZN(G284) );
  NOR2_X1 U857 ( .A1(G286), .A2(n814), .ZN(n775) );
  NOR2_X1 U858 ( .A1(G868), .A2(G299), .ZN(n774) );
  NOR2_X1 U859 ( .A1(n775), .A2(n774), .ZN(G297) );
  NAND2_X1 U860 ( .A1(n776), .A2(G559), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n777), .A2(n990), .ZN(n778) );
  XNOR2_X1 U862 ( .A(n778), .B(KEYINPUT83), .ZN(n779) );
  XOR2_X1 U863 ( .A(KEYINPUT16), .B(n779), .Z(G148) );
  NOR2_X1 U864 ( .A1(n978), .A2(G868), .ZN(n782) );
  NAND2_X1 U865 ( .A1(G868), .A2(n990), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(G282) );
  XNOR2_X1 U868 ( .A(G2100), .B(KEYINPUT85), .ZN(n792) );
  NAND2_X1 U869 ( .A1(G123), .A2(n885), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT18), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(KEYINPUT84), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G111), .A2(n886), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G135), .A2(n889), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G99), .A2(n890), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n925) );
  XNOR2_X1 U878 ( .A(n925), .B(G2096), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(G156) );
  NAND2_X1 U880 ( .A1(G559), .A2(n990), .ZN(n793) );
  XNOR2_X1 U881 ( .A(n793), .B(n978), .ZN(n811) );
  NOR2_X1 U882 ( .A1(G860), .A2(n811), .ZN(n803) );
  NAND2_X1 U883 ( .A1(n540), .A2(G67), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G55), .A2(n794), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G80), .A2(n797), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G93), .A2(n798), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n813) );
  XOR2_X1 U890 ( .A(n803), .B(n813), .Z(G145) );
  XOR2_X1 U891 ( .A(n813), .B(G288), .Z(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(G290), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT19), .B(n805), .ZN(n807) );
  XNOR2_X1 U894 ( .A(G305), .B(KEYINPUT87), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U896 ( .A(n809), .B(n808), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n810), .B(G303), .ZN(n902) );
  XNOR2_X1 U898 ( .A(n902), .B(n811), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n812), .A2(G868), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n816), .A2(n815), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n817) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n817), .Z(n818) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n818), .ZN(n819) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n819), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n821) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U910 ( .A1(G218), .A2(n822), .ZN(n823) );
  NAND2_X1 U911 ( .A1(G96), .A2(n823), .ZN(n836) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n836), .ZN(n827) );
  NAND2_X1 U913 ( .A1(G120), .A2(G108), .ZN(n824) );
  NOR2_X1 U914 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G69), .A2(n825), .ZN(n837) );
  NAND2_X1 U916 ( .A1(G567), .A2(n837), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U918 ( .A(KEYINPUT88), .B(n828), .Z(G319) );
  INV_X1 U919 ( .A(G319), .ZN(n830) );
  NAND2_X1 U920 ( .A1(G661), .A2(G483), .ZN(n829) );
  NOR2_X1 U921 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U922 ( .A(KEYINPUT89), .B(n831), .Z(n835) );
  NAND2_X1 U923 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U926 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U929 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XOR2_X1 U935 ( .A(G2096), .B(G2100), .Z(n839) );
  XNOR2_X1 U936 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U938 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U941 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2084), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U944 ( .A(KEYINPUT41), .B(G1956), .Z(n847) );
  XNOR2_X1 U945 ( .A(G1976), .B(G1961), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U947 ( .A(n848), .B(KEYINPUT112), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U950 ( .A(G1986), .B(G1971), .Z(n852) );
  XNOR2_X1 U951 ( .A(G1981), .B(G1966), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U954 ( .A(KEYINPUT111), .B(G2474), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n885), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G112), .A2(n886), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G100), .A2(n890), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(KEYINPUT114), .B(n860), .Z(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G136), .A2(n889), .ZN(n863) );
  XNOR2_X1 U964 ( .A(KEYINPUT113), .B(n863), .ZN(n864) );
  NOR2_X1 U965 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G127), .A2(n885), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G115), .A2(n886), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n868), .B(KEYINPUT47), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G103), .A2(n890), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G139), .A2(n889), .ZN(n871) );
  XNOR2_X1 U973 ( .A(KEYINPUT115), .B(n871), .ZN(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n933) );
  XNOR2_X1 U975 ( .A(n874), .B(n933), .ZN(n877) );
  XNOR2_X1 U976 ( .A(G160), .B(n875), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n881) );
  XOR2_X1 U978 ( .A(KEYINPUT116), .B(KEYINPUT48), .Z(n879) );
  XNOR2_X1 U979 ( .A(n925), .B(KEYINPUT46), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(n881), .B(n880), .Z(n884) );
  XOR2_X1 U982 ( .A(G164), .B(n882), .Z(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n898) );
  NAND2_X1 U984 ( .A1(G130), .A2(n885), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G118), .A2(n886), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U987 ( .A1(G142), .A2(n889), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G106), .A2(n890), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(KEYINPUT45), .B(n893), .Z(n894) );
  NOR2_X1 U991 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U992 ( .A(G162), .B(n896), .Z(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U994 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U995 ( .A(G286), .B(n978), .Z(n901) );
  XNOR2_X1 U996 ( .A(G171), .B(n990), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U999 ( .A1(G37), .A2(n904), .ZN(G397) );
  XOR2_X1 U1000 ( .A(G2443), .B(G2451), .Z(n906) );
  XNOR2_X1 U1001 ( .A(KEYINPUT109), .B(G2427), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1003 ( .A(KEYINPUT110), .B(G2438), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G2435), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1006 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1007 ( .A(G2446), .B(KEYINPUT108), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n915) );
  XOR2_X1 U1009 ( .A(G1348), .B(G1341), .Z(n913) );
  XNOR2_X1 U1010 ( .A(G2430), .B(n913), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1012 ( .A1(G14), .A2(n916), .ZN(n923) );
  NAND2_X1 U1013 ( .A1(n923), .A2(G319), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n917) );
  XOR2_X1 U1015 ( .A(KEYINPUT49), .B(n917), .Z(n918) );
  XNOR2_X1 U1016 ( .A(n918), .B(KEYINPUT117), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  INV_X1 U1022 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT119), .B(n924), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT120), .B(n929), .ZN(n948) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n932), .Z(n946) );
  XNOR2_X1 U1031 ( .A(G2072), .B(n933), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(G164), .B(G2078), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(n936), .B(KEYINPUT50), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n937), .B(KEYINPUT121), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n944) );
  INV_X1 U1037 ( .A(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(n949), .ZN(n950) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n970), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n951), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1046 ( .A(G2090), .B(G35), .ZN(n965) );
  XOR2_X1 U1047 ( .A(G2067), .B(G26), .Z(n952) );
  NAND2_X1 U1048 ( .A1(n952), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1049 ( .A(G1996), .B(G32), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n955), .B(G27), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G25), .B(n956), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n966), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n970), .B(n969), .ZN(n972) );
  INV_X1 U1063 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n973), .ZN(n1028) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XNOR2_X1 U1067 ( .A(G166), .B(G1971), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G1956), .B(G299), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(KEYINPUT57), .B(KEYINPUT123), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G168), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT122), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n987), .B(n986), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n997) );
  XOR2_X1 U1080 ( .A(G1348), .B(n990), .Z(n992) );
  XOR2_X1 U1081 ( .A(G171), .B(G1961), .Z(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT124), .B(n993), .Z(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1026) );
  INV_X1 U1087 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(n1000), .B(G4), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G1956), .B(G20), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT125), .B(G1981), .Z(n1005) );
  XNOR2_X1 U1095 ( .A(G6), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(KEYINPUT126), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G21), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  XNOR2_X1 U1103 ( .A(G1976), .B(G23), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G1986), .B(KEYINPUT127), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(n1016), .B(G24), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

