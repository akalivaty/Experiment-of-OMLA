//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n212), .B1(new_n213), .B2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n215), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT0), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(new_n219), .B2(new_n218), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n213), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n222), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n224), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n248), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G274), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n260), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(G226), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n255), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G222), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n269), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n267), .B2(new_n268), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT69), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n276), .B2(G223), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n265), .B(G190), .C1(new_n277), .C2(new_n257), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n278), .B(KEYINPUT72), .Z(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n280), .A2(new_n208), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n255), .A2(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n283), .A2(new_n284), .B1(G150), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n203), .A2(G20), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n281), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n280), .A2(new_n208), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G50), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G50), .B2(new_n290), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n277), .A2(new_n257), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n265), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n279), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT73), .A3(new_n300), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n279), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n304), .A2(new_n265), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n297), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(G169), .C2(new_n311), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n293), .A2(G77), .A3(new_n294), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n291), .A2(new_n273), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n283), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n320));
  INV_X1    g0120(.A(new_n284), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n292), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n318), .A2(KEYINPUT71), .A3(new_n324), .A4(new_n319), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n262), .B1(G244), .B2(new_n264), .ZN(new_n330));
  INV_X1    g0130(.A(G232), .ZN(new_n331));
  INV_X1    g0131(.A(G107), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n271), .A2(new_n331), .B1(new_n332), .B2(new_n269), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n276), .B2(G238), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n334), .B2(new_n257), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(G179), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n329), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(G200), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n327), .A3(new_n328), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  AND4_X1   g0144(.A1(new_n308), .A2(new_n310), .A3(new_n315), .A4(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT74), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n269), .A2(G1698), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n331), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n275), .A2(KEYINPUT74), .A3(G232), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  INV_X1    g0151(.A(G226), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n271), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n257), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n262), .B1(G238), .B2(new_n264), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT13), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n353), .B1(new_n348), .B2(new_n349), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n356), .B(new_n359), .C1(new_n360), .C2(new_n257), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(new_n361), .A3(KEYINPUT75), .ZN(new_n362));
  INV_X1    g0162(.A(new_n355), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT75), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(new_n359), .A4(new_n356), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(G169), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n362), .A2(new_n365), .A3(KEYINPUT14), .A4(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n358), .A2(G179), .A3(new_n361), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n291), .A2(new_n224), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n224), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n321), .B2(new_n273), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n293), .A2(G68), .A3(new_n294), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT11), .B1(new_n377), .B2(new_n292), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n362), .A2(G200), .A3(new_n365), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n358), .A2(new_n361), .A3(G190), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(new_n382), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n345), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n282), .B1(new_n289), .B2(G20), .ZN(new_n389));
  AOI211_X1 g0189(.A(new_n291), .B(new_n292), .C1(new_n389), .C2(KEYINPUT79), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(KEYINPUT79), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n390), .A2(new_n392), .B1(new_n291), .B2(new_n282), .ZN(new_n393));
  INV_X1    g0193(.A(G58), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n224), .ZN(new_n395));
  OAI21_X1  g0195(.A(G20), .B1(new_n395), .B2(new_n201), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n285), .A2(G159), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(KEYINPUT3), .A2(G33), .ZN(new_n401));
  NOR2_X1   g0201(.A1(KEYINPUT3), .A2(G33), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT76), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT76), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n267), .A2(new_n404), .A3(new_n268), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n405), .A3(new_n209), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n401), .A2(new_n402), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT77), .B1(new_n411), .B2(G68), .ZN(new_n412));
  NOR4_X1   g0212(.A1(new_n401), .A2(new_n402), .A3(new_n407), .A4(G20), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n406), .B2(new_n407), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT77), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n414), .A2(new_n415), .A3(new_n224), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n400), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n407), .B1(new_n269), .B2(G20), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n224), .B1(new_n418), .B2(new_n410), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n399), .B1(new_n419), .B2(new_n398), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n292), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT78), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n400), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n411), .A2(KEYINPUT77), .A3(G68), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n415), .B1(new_n414), .B2(new_n224), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT78), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n427), .A2(new_n428), .A3(new_n421), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n393), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n269), .A2(G226), .A3(G1698), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT80), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n275), .A2(KEYINPUT80), .A3(G226), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n269), .A2(G223), .A3(new_n270), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G87), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(KEYINPUT81), .B(new_n263), .C1(new_n436), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT81), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n434), .B2(new_n435), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n257), .ZN(new_n443));
  INV_X1    g0243(.A(new_n262), .ZN(new_n444));
  INV_X1    g0244(.A(new_n264), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n331), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G179), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n442), .A2(new_n257), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n337), .B1(new_n449), .B2(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n430), .A2(new_n431), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n393), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n428), .B1(new_n427), .B2(new_n421), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n417), .A2(KEYINPUT78), .A3(new_n422), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT18), .B1(new_n457), .B2(new_n451), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n340), .A2(KEYINPUT82), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n340), .A2(KEYINPUT82), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n446), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n440), .A2(new_n443), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n303), .B1(new_n449), .B2(new_n446), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n393), .B(new_n467), .C1(new_n423), .C2(new_n429), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n457), .A2(KEYINPUT17), .A3(new_n467), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n459), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n388), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n209), .C1(G33), .C2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n478), .B(new_n292), .C1(new_n209), .C2(G116), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n479), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  XOR2_X1   g0281(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n482));
  AND2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n290), .A2(G116), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n289), .A2(G33), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n281), .A2(new_n290), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n488), .B2(G116), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n275), .A2(G264), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n269), .A2(G257), .A3(new_n270), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n409), .A2(G303), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n263), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT5), .B(G41), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n259), .A2(G1), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n496), .A2(new_n257), .A3(G274), .A4(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n263), .B1(new_n497), .B2(new_n496), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G270), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n490), .A2(new_n501), .A3(G169), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT89), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(KEYINPUT21), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n480), .A2(new_n483), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n337), .B1(new_n507), .B2(new_n489), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n504), .B1(new_n508), .B2(new_n501), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n490), .A2(G179), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n506), .A2(new_n509), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n501), .A2(G200), .ZN(new_n512));
  INV_X1    g0312(.A(new_n490), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n513), .C1(new_n462), .C2(new_n501), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n514), .A2(KEYINPUT90), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(KEYINPUT90), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(G1698), .C1(new_n401), .C2(new_n402), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT85), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n269), .A2(KEYINPUT85), .A3(G244), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n255), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(G1698), .B1(new_n267), .B2(new_n268), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G238), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n257), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n497), .A2(new_n227), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n257), .ZN(new_n529));
  INV_X1    g0329(.A(new_n497), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n258), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n337), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n322), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n290), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n284), .A2(new_n535), .A3(G97), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n226), .B1(new_n351), .B2(new_n209), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n538), .B2(new_n535), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n269), .A2(KEYINPUT86), .A3(new_n209), .A4(G68), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n209), .B(G68), .C1(new_n401), .C2(new_n402), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT86), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n534), .B1(new_n544), .B2(new_n292), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n488), .A2(new_n533), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n531), .ZN(new_n548));
  OAI211_X1 g0348(.A(G238), .B(new_n270), .C1(new_n401), .C2(new_n402), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n255), .B2(new_n523), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n520), .B2(new_n521), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n312), .B(new_n548), .C1(new_n551), .C2(new_n257), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n532), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G190), .B(new_n548), .C1(new_n551), .C2(new_n257), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n487), .A2(new_n226), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n534), .B(new_n557), .C1(new_n544), .C2(new_n292), .ZN(new_n558));
  OAI21_X1  g0358(.A(G200), .B1(new_n527), .B2(new_n531), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n556), .B1(new_n560), .B2(KEYINPUT87), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT87), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n554), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n209), .B(G87), .C1(new_n401), .C2(new_n402), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT91), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT22), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n269), .A2(new_n209), .A3(G87), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n209), .B2(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n332), .A2(KEYINPUT23), .A3(G20), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(new_n524), .B2(new_n209), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n571), .B1(new_n570), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n292), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT25), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n290), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n332), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n488), .A2(G107), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n269), .A2(G250), .A3(new_n270), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G294), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n263), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n499), .A2(G264), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n498), .ZN(new_n592));
  OAI21_X1  g0392(.A(G169), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT92), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n588), .A2(new_n263), .B1(G264), .B2(new_n499), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT92), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(G179), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n584), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n498), .B1(new_n596), .B2(KEYINPUT92), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n589), .A2(KEYINPUT92), .A3(new_n590), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n303), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n591), .A2(G190), .A3(new_n592), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n583), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G250), .B(G1698), .C1(new_n401), .C2(new_n402), .ZN(new_n607));
  OAI211_X1 g0407(.A(G244), .B(new_n270), .C1(new_n401), .C2(new_n402), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT4), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n476), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT4), .B1(new_n525), .B2(G244), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n263), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n496), .A2(new_n497), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(G257), .A3(new_n257), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n614), .A2(new_n498), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n291), .A2(new_n477), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n487), .B2(new_n477), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT7), .B1(new_n409), .B2(new_n209), .ZN(new_n621));
  OAI21_X1  g0421(.A(G107), .B1(new_n621), .B2(new_n413), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT6), .ZN(new_n623));
  AND2_X1   g0423(.A1(G97), .A2(G107), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n623), .B1(new_n624), .B2(new_n537), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n332), .A2(KEYINPUT6), .A3(G97), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(G20), .B1(G77), .B2(new_n285), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n281), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT83), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(KEYINPUT83), .B(new_n281), .C1(new_n622), .C2(new_n628), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n617), .B(new_n620), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT84), .B1(new_n616), .B2(new_n340), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n612), .A2(new_n615), .A3(new_n635), .A4(G190), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n285), .A2(G77), .ZN(new_n638));
  INV_X1    g0438(.A(new_n626), .ZN(new_n639));
  XNOR2_X1  g0439(.A(G97), .B(G107), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n623), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n638), .B1(new_n641), .B2(new_n209), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n332), .B1(new_n418), .B2(new_n410), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n292), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT83), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n629), .A2(new_n630), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n619), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n616), .A2(new_n337), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n612), .A2(new_n615), .A3(new_n312), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n633), .A2(new_n637), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n517), .A2(new_n564), .A3(new_n606), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n475), .A2(new_n653), .ZN(G372));
  INV_X1    g0454(.A(new_n315), .ZN(new_n655));
  INV_X1    g0455(.A(new_n339), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n373), .A2(new_n383), .B1(new_n387), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n470), .A2(new_n471), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n459), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n308), .A2(new_n310), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n647), .A2(new_n650), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n564), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT93), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n647), .B2(new_n650), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n648), .A2(new_n649), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n620), .B1(new_n631), .B2(new_n632), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT93), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n558), .A2(new_n559), .A3(new_n555), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n670), .A2(new_n553), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n662), .A2(new_n666), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n670), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n651), .A2(new_n605), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n598), .A2(new_n593), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n583), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n510), .A2(new_n501), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n502), .A2(new_n505), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n508), .A2(new_n501), .A3(new_n504), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n554), .B1(new_n675), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n661), .B1(new_n475), .B2(new_n685), .ZN(G369));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n289), .A2(new_n209), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n517), .B1(new_n513), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n511), .A2(new_n490), .A3(new_n693), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n687), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n606), .B1(new_n584), .B2(new_n694), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n599), .A2(new_n693), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n681), .A2(new_n693), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n606), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n677), .B2(new_n693), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n702), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n217), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n537), .A2(new_n226), .A3(new_n523), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n708), .A2(new_n289), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n207), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  NAND3_X1  g0512(.A1(new_n564), .A2(new_n662), .A3(new_n663), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n670), .A2(new_n553), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n663), .B2(KEYINPUT93), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n715), .A2(new_n666), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n713), .B1(new_n716), .B2(new_n662), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n599), .A2(new_n511), .ZN(new_n718));
  AOI21_X1  g0518(.A(G200), .B1(new_n595), .B2(new_n597), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n584), .B1(new_n719), .B2(new_n603), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n667), .A2(new_n668), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n647), .A2(new_n617), .A3(new_n634), .A4(new_n636), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n670), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n553), .B1(new_n718), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n694), .B1(new_n717), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n684), .A2(new_n727), .A3(new_n694), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n616), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n527), .A2(new_n531), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n495), .A4(new_n500), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  OR3_X1    g0533(.A1(new_n598), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n595), .A2(new_n597), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n731), .A2(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n616), .A3(new_n501), .A4(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n598), .B2(new_n732), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n693), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n742), .B(new_n743), .C1(new_n653), .C2(new_n693), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n729), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n712), .B1(new_n747), .B2(G1), .ZN(G364));
  NAND3_X1  g0548(.A1(new_n695), .A2(new_n687), .A3(new_n696), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n209), .A2(G13), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n289), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n708), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n697), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n755), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n707), .A2(new_n409), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n523), .B2(new_n707), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n403), .A2(new_n405), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n217), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n207), .A2(new_n259), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n253), .B2(new_n259), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n759), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n215), .A2(new_n255), .A3(KEYINPUT96), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT96), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G13), .B2(G33), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n208), .B1(G20), .B2(new_n337), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n757), .B1(new_n767), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(KEYINPUT97), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n777), .A2(KEYINPUT97), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n303), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G20), .A3(G190), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n409), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G20), .A3(new_n340), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(G329), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n209), .A2(new_n312), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n303), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n209), .B1(new_n784), .B2(G190), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n788), .A2(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n462), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(G326), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n780), .A2(G20), .A3(new_n340), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n787), .B(new_n798), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n796), .A2(G190), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT100), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n808), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(KEYINPUT100), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n462), .A2(new_n789), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G322), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n810), .A2(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT101), .ZN(new_n817));
  INV_X1    g0617(.A(new_n797), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n269), .B1(new_n226), .B2(new_n781), .C1(new_n818), .C2(new_n202), .ZN(new_n819));
  INV_X1    g0619(.A(G159), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n785), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT32), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n794), .A2(new_n477), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n819), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n790), .A2(G77), .B1(new_n821), .B2(new_n822), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n813), .A2(G58), .B1(new_n807), .B2(G68), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n804), .A2(new_n332), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n806), .A2(new_n817), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n778), .B(new_n779), .C1(new_n774), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n695), .A2(new_n696), .A3(new_n773), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n749), .A2(new_n756), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  OAI221_X1 g0634(.A(new_n409), .B1(new_n785), .B2(new_n792), .C1(new_n781), .C2(new_n332), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n818), .A2(new_n782), .B1(new_n791), .B2(new_n523), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(G283), .C2(new_n807), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n824), .B1(new_n813), .B2(G294), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT102), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n803), .A2(G87), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n781), .A2(new_n202), .B1(new_n843), .B2(new_n785), .ZN(new_n844));
  INV_X1    g0644(.A(new_n794), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n844), .B(new_n761), .C1(G58), .C2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n804), .B2(new_n224), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n797), .A2(G137), .B1(new_n790), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  INV_X1    g0650(.A(new_n807), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n848), .B1(new_n849), .B2(new_n814), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT34), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n842), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n774), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n771), .A2(new_n774), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n757), .B1(new_n273), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n329), .A2(new_n693), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n343), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n860), .A2(new_n339), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n339), .A2(new_n693), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n856), .B(new_n858), .C1(new_n863), .C2(new_n772), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n863), .B(KEYINPUT104), .Z(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n685), .B2(new_n693), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n344), .A2(new_n694), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n564), .A2(new_n663), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT26), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n715), .A2(new_n662), .A3(new_n666), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n868), .B1(new_n872), .B2(new_n724), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n755), .B1(new_n874), .B2(new_n745), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n745), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n864), .B1(new_n876), .B2(new_n877), .ZN(G384));
  OR2_X1    g0678(.A1(new_n627), .A2(KEYINPUT35), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n627), .A2(KEYINPUT35), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(G116), .A3(new_n210), .A4(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT36), .Z(new_n882));
  OAI211_X1 g0682(.A(new_n207), .B(G77), .C1(new_n394), .C2(new_n224), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n289), .B(G13), .C1(new_n883), .C2(new_n249), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n867), .B1(new_n673), .B2(new_n683), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT105), .B1(new_n886), .B2(new_n862), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT105), .ZN(new_n888));
  INV_X1    g0688(.A(new_n862), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n873), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n371), .B1(new_n368), .B2(new_n369), .ZN(new_n892));
  OAI211_X1 g0692(.A(KEYINPUT106), .B(new_n387), .C1(new_n892), .C2(new_n382), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n382), .A2(new_n694), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n373), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT106), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(new_n387), .C1(new_n892), .C2(new_n382), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n893), .A2(new_n896), .B1(new_n898), .B2(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n691), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n417), .A2(new_n292), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n425), .A2(new_n426), .ZN(new_n903));
  INV_X1    g0703(.A(new_n398), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT16), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n393), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n453), .A2(new_n458), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n901), .B(new_n906), .C1(new_n907), .C2(new_n658), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n468), .B1(new_n457), .B2(new_n451), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT107), .B(KEYINPUT37), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n457), .B2(new_n691), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n451), .A2(new_n691), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n457), .A2(new_n467), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n909), .A2(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n908), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n906), .A2(new_n901), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n459), .B2(new_n472), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(KEYINPUT38), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n900), .A2(new_n921), .B1(new_n459), .B2(new_n901), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n916), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT109), .B1(new_n918), .B2(new_n919), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT109), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n908), .A2(new_n926), .A3(KEYINPUT38), .A4(new_n915), .ZN(new_n927));
  INV_X1    g0727(.A(new_n910), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n457), .A2(new_n691), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n909), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT108), .B1(new_n909), .B2(new_n911), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n928), .B1(new_n430), .B2(new_n901), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n430), .A2(new_n452), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n468), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n929), .B1(new_n907), .B2(new_n658), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n925), .B(new_n927), .C1(new_n938), .C2(KEYINPUT38), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n924), .B1(new_n939), .B2(new_n923), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n384), .A2(new_n693), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n922), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n726), .A2(new_n728), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n474), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n661), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n942), .B(new_n945), .Z(new_n946));
  AND2_X1   g0746(.A1(new_n744), .A2(new_n863), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n939), .A2(KEYINPUT40), .A3(new_n899), .A4(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n899), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n921), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n474), .A2(new_n744), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n687), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n946), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n289), .B2(new_n752), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n946), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n885), .B1(new_n958), .B2(new_n959), .ZN(G367));
  NOR2_X1   g0760(.A1(new_n558), .A2(new_n694), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT111), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n714), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n554), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n773), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n775), .B1(new_n217), .B2(new_n322), .C1(new_n764), .C2(new_n240), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n755), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n791), .A2(new_n805), .B1(new_n332), .B2(new_n794), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(KEYINPUT112), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n851), .A2(new_n793), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n781), .A2(new_n523), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n818), .A2(new_n792), .B1(new_n971), .B2(KEYINPUT46), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n968), .A2(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n813), .A2(G303), .B1(new_n971), .B2(KEYINPUT46), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n760), .B1(G317), .B2(new_n786), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n477), .C2(new_n802), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n807), .A2(G159), .B1(G68), .B2(new_n845), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n202), .B2(new_n791), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n781), .A2(new_n394), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n409), .B(new_n981), .C1(G137), .C2(new_n786), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G143), .A2(new_n797), .B1(new_n813), .B2(G150), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n273), .C2(new_n802), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n975), .A2(new_n978), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT47), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n967), .B1(new_n986), .B2(new_n774), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n965), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n652), .B1(new_n647), .B2(new_n694), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n663), .A2(new_n693), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n705), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT44), .Z(new_n993));
  NOR2_X1   g0793(.A1(new_n705), .A2(new_n991), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT45), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n993), .A2(new_n701), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n701), .B1(new_n993), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n703), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n698), .A2(new_n699), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n704), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(new_n697), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n746), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n747), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n708), .B(KEYINPUT41), .Z(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n754), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n964), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n991), .A2(new_n704), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT42), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n989), .A2(new_n677), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n693), .B1(new_n1014), .B2(new_n721), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n964), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(KEYINPUT43), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1009), .A3(new_n964), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n701), .A2(new_n991), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1022), .B(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n988), .B1(new_n1008), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT113), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(KEYINPUT113), .B(new_n988), .C1(new_n1008), .C2(new_n1025), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(G387));
  INV_X1    g0831(.A(new_n708), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n1003), .A2(KEYINPUT118), .A3(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n746), .A2(new_n1002), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT119), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT118), .B1(new_n1003), .B2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(KEYINPUT119), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1002), .A2(new_n753), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n698), .A2(new_n699), .A3(new_n773), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n709), .C1(G68), .C2(G77), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT50), .B1(new_n282), .B2(G50), .ZN(new_n1046));
  OR3_X1    g0846(.A1(new_n282), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT115), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1047), .C1(new_n1043), .C2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n763), .B1(new_n1045), .B2(new_n1049), .C1(new_n259), .C2(new_n244), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n758), .A2(new_n709), .B1(new_n332), .B2(new_n707), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n757), .B1(new_n1052), .B2(new_n775), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT116), .Z(new_n1054));
  INV_X1    g0854(.A(new_n781), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(G77), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n760), .C1(new_n850), .C2(new_n785), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n851), .A2(new_n282), .B1(new_n791), .B2(new_n224), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G159), .C2(new_n797), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n794), .A2(new_n322), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n813), .B2(G50), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT117), .Z(new_n1062));
  OAI211_X1 g0862(.A(new_n1059), .B(new_n1062), .C1(new_n477), .C2(new_n804), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n760), .B1(G326), .B2(new_n786), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n781), .A2(new_n793), .B1(new_n794), .B2(new_n805), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n813), .A2(G317), .B1(new_n790), .B2(G303), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n792), .B2(new_n851), .C1(new_n815), .C2(new_n818), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1064), .B1(new_n523), .B2(new_n802), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1063), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1054), .B1(new_n774), .B2(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1040), .A2(new_n1041), .B1(new_n1042), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1038), .A2(new_n1076), .ZN(G393));
  NAND2_X1  g0877(.A1(new_n991), .A2(new_n773), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n775), .B1(new_n477), .B2(new_n217), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n763), .B2(new_n248), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n409), .B1(new_n785), .B2(new_n815), .C1(new_n781), .C2(new_n805), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n790), .A2(G294), .B1(G116), .B2(new_n845), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n782), .B2(new_n851), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n829), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G311), .A2(new_n813), .B1(new_n797), .B2(G317), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n781), .A2(new_n224), .B1(new_n849), .B2(new_n785), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n794), .A2(new_n273), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n761), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT121), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G50), .A2(new_n807), .B1(new_n790), .B2(new_n283), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n840), .B(new_n1089), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G150), .A2(new_n797), .B1(new_n813), .B2(G159), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1092), .A2(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1084), .A2(new_n1086), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n757), .B(new_n1080), .C1(new_n1099), .C2(new_n774), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n998), .A2(new_n754), .B1(new_n1078), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1004), .A2(new_n708), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n998), .A2(new_n1003), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(G390));
  NAND3_X1  g0904(.A1(new_n744), .A2(G330), .A3(new_n863), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n893), .A2(new_n896), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n898), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n894), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n941), .B1(new_n891), .B2(new_n899), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n925), .A2(new_n927), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT38), .B1(new_n936), .B2(new_n937), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n923), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n921), .A2(KEYINPUT39), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n889), .B1(new_n725), .B2(new_n861), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n941), .B1(new_n1116), .B2(new_n899), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n939), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1109), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1109), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n1118), .C1(new_n940), .C2(new_n1110), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n944), .B(new_n661), .C1(new_n475), .C2(new_n745), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1109), .A2(new_n1116), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1108), .B1(new_n865), .B2(new_n745), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n891), .B1(new_n1127), .B2(new_n1109), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1123), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1120), .A2(new_n1122), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT122), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT122), .A4(new_n1129), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1032), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT123), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT123), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1120), .A2(new_n1137), .A3(new_n1122), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1123), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1120), .A2(new_n754), .A3(new_n1122), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n757), .B1(new_n282), .B2(new_n857), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n804), .A2(new_n224), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n409), .B1(new_n785), .B2(new_n793), .C1(new_n781), .C2(new_n226), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1088), .B(new_n1147), .C1(G116), .C2(new_n813), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n797), .A2(G283), .B1(new_n790), .B2(G97), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n332), .C2(new_n851), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n781), .A2(new_n850), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n843), .B2(new_n814), .C1(new_n820), .C2(new_n794), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n409), .B1(new_n786), .B2(G125), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n791), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n797), .A2(G128), .B1(new_n807), .B2(G137), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n202), .C2(new_n802), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1146), .A2(new_n1150), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT124), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n774), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1145), .B1(new_n1162), .B2(new_n1164), .C1(new_n940), .C2(new_n772), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1144), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1143), .A2(new_n1167), .ZN(G378));
  AOI22_X1  g0968(.A1(G97), .A2(new_n807), .B1(new_n790), .B2(new_n533), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n332), .B2(new_n814), .C1(new_n523), .C2(new_n818), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n761), .A2(new_n256), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n802), .A2(new_n394), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1056), .B1(new_n224), .B2(new_n794), .C1(new_n805), .C2(new_n785), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G50), .B1(new_n255), .B2(new_n256), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1174), .A2(KEYINPUT58), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n813), .A2(G128), .B1(new_n790), .B2(G137), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n797), .A2(G125), .B1(new_n807), .B2(G132), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1155), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1055), .A2(new_n1179), .B1(new_n845), .B2(G150), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G33), .B(G41), .C1(new_n786), .C2(G124), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n820), .C2(new_n802), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1176), .B1(KEYINPUT58), .B2(new_n1174), .C1(new_n1182), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n774), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n757), .B1(new_n202), .B2(new_n857), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n660), .A2(new_n315), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n314), .A2(new_n901), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1187), .B(new_n1188), .C1(new_n1193), .C2(new_n772), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1193), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n952), .B2(new_n687), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n948), .A3(G330), .A4(new_n951), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1196), .A2(new_n942), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n942), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1194), .B1(new_n1200), .B2(new_n753), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1140), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT57), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1123), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n708), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1202), .B1(new_n1206), .B2(new_n1209), .ZN(G375));
  OAI221_X1 g1010(.A(new_n409), .B1(new_n785), .B2(new_n782), .C1(new_n781), .C2(new_n477), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1060), .B(new_n1211), .C1(G283), .C2(new_n813), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n797), .A2(G294), .B1(new_n790), .B2(G107), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n523), .C2(new_n851), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G77), .B2(new_n803), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n813), .A2(G137), .B1(new_n807), .B2(new_n1179), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n843), .B2(new_n818), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n790), .A2(G150), .B1(G50), .B2(new_n845), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1055), .A2(G159), .B1(new_n786), .B2(G128), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n760), .A3(new_n1222), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1219), .A2(new_n1220), .A3(new_n1172), .A4(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n774), .B1(new_n1215), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n757), .B1(new_n224), .B2(new_n857), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1108), .B2(new_n771), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1139), .B2(new_n754), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1141), .A2(new_n1007), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(G381));
  AOI21_X1  g1032(.A(new_n1166), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(G390), .A2(G381), .A3(G384), .ZN(new_n1235));
  AND4_X1   g1035(.A1(new_n1030), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G375), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1236), .A2(new_n1237), .A3(KEYINPUT126), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT126), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(new_n1239), .ZN(G407));
  INV_X1    g1040(.A(G213), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G378), .A2(G343), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1244), .B(new_n1245), .ZN(G409));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1241), .A2(G343), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G378), .B(new_n1202), .C1(new_n1206), .C2(new_n1209), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1207), .A2(new_n1200), .A3(new_n1006), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1233), .B1(new_n1250), .B2(new_n1201), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1248), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1231), .A2(KEYINPUT60), .A3(new_n1141), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n708), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1231), .B1(KEYINPUT60), .B2(new_n1141), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1229), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1248), .A2(G2897), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1258), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1247), .B1(new_n1252), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1248), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1268), .B1(new_n1271), .B2(new_n1260), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(G393), .B(G396), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(G390), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1273), .A2(KEYINPUT113), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(G390), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(new_n1026), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1260), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1267), .A2(new_n1272), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1252), .A2(new_n1281), .A3(new_n1278), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1252), .B2(new_n1278), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1282), .A2(new_n1266), .A3(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1280), .B1(new_n1284), .B2(new_n1277), .ZN(G405));
  XOR2_X1   g1085(.A(new_n1276), .B(new_n1026), .Z(new_n1286));
  NAND2_X1  g1086(.A1(G375), .A2(new_n1233), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1249), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1278), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1260), .A3(new_n1249), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1286), .B(new_n1291), .ZN(G402));
endmodule


