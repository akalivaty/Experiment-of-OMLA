//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT78), .ZN(new_n203));
  XOR2_X1   g002(.A(G57gat), .B(G85gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n209), .A2(new_n211), .B1(KEYINPUT2), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT74), .ZN(new_n216));
  XOR2_X1   g015(.A(G155gat), .B(G162gat), .Z(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n215), .B(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n213), .A2(new_n217), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT68), .B(G120gat), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n227), .A2(G120gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n233), .B2(new_n224), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n223), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT75), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245));
  INV_X1    g044(.A(new_n242), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n246), .B1(new_n237), .B2(new_n239), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT5), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n238), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n236), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n253), .A2(new_n246), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n256), .A3(new_n235), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n244), .A2(new_n249), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(KEYINPUT79), .A3(new_n257), .ZN(new_n260));
  OR3_X1    g059(.A1(new_n239), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n248), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(new_n246), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n207), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(new_n246), .A3(new_n253), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT76), .B1(new_n243), .B2(KEYINPUT5), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n247), .A2(new_n245), .A3(new_n248), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n262), .A2(new_n263), .ZN(new_n270));
  INV_X1    g069(.A(new_n207), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n265), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(KEYINPUT6), .B(new_n207), .C1(new_n259), .C2(new_n264), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT26), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT27), .B(G183gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT67), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n284));
  OAI221_X1 g083(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n291), .A2(KEYINPUT26), .A3(new_n279), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n285), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(KEYINPUT23), .B2(new_n279), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n296), .A2(KEYINPUT65), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  NOR2_X1   g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n277), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n300), .B2(new_n277), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(KEYINPUT65), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n297), .A2(new_n298), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n294), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n302), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n295), .B1(new_n294), .B2(new_n305), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT25), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G226gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  OAI22_X1  g112(.A1(new_n311), .A2(KEYINPUT29), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n293), .B2(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT22), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT72), .B(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n323), .A2(new_n318), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n324), .B2(new_n319), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(G218gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(G218gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n317), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n285), .ZN(new_n331));
  INV_X1    g130(.A(new_n292), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n287), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n310), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT29), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n328), .B(new_n316), .C1(new_n335), .C2(new_n315), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n330), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  INV_X1    g140(.A(new_n336), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n328), .B1(new_n314), .B2(new_n316), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n344), .A3(KEYINPUT30), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n336), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n341), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n350));
  AND3_X1   g149(.A1(new_n276), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G228gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(new_n313), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n329), .B1(new_n252), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n326), .A2(new_n354), .A3(new_n327), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n238), .B1(new_n356), .B2(new_n251), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(KEYINPUT83), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n326), .A2(new_n360), .A3(new_n354), .A4(new_n327), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n251), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n355), .B1(new_n362), .B2(new_n223), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n353), .B(new_n358), .C1(new_n363), .C2(KEYINPUT82), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n363), .A2(new_n365), .B1(new_n352), .B2(new_n313), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G22gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n366), .A3(G22gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT81), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT31), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G50gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n370), .B2(KEYINPUT84), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n369), .B(new_n370), .C1(KEYINPUT84), .C2(new_n375), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n333), .A2(KEYINPUT69), .A3(new_n334), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n293), .B2(new_n310), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n383), .A3(new_n236), .ZN(new_n384));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT64), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n333), .A2(new_n334), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n382), .A3(new_n235), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(G15gat), .B(G43gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT33), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(KEYINPUT32), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(KEYINPUT70), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n389), .A2(KEYINPUT32), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n392), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT70), .B1(new_n389), .B2(new_n395), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT34), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n388), .ZN(new_n402));
  INV_X1    g201(.A(new_n386), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(KEYINPUT34), .B(new_n386), .C1(new_n384), .C2(new_n388), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n406), .B(new_n394), .C1(new_n398), .C2(new_n399), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n408), .A2(KEYINPUT87), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT87), .B1(new_n408), .B2(new_n409), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n351), .B(new_n380), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n276), .A2(new_n413), .A3(new_n349), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n408), .A2(new_n377), .A3(new_n409), .A4(new_n378), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n276), .B2(new_n349), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT35), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n412), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n349), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n260), .A2(new_n261), .A3(new_n253), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n242), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n422), .A2(KEYINPUT39), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(KEYINPUT39), .C1(new_n242), .C2(new_n240), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n271), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT40), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT40), .A4(new_n271), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n420), .A2(new_n427), .A3(new_n265), .A4(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n276), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT37), .B1(new_n330), .B2(new_n336), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n341), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n330), .A2(KEYINPUT37), .A3(new_n336), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n432), .A2(KEYINPUT85), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n434), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n433), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n440), .A2(new_n341), .A3(new_n431), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n344), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n380), .B(new_n429), .C1(new_n437), .C2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n379), .B1(new_n414), .B2(new_n416), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n408), .A2(new_n409), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT71), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT36), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT36), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n443), .A2(new_n444), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n419), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G15gat), .B(G22gat), .ZN(new_n453));
  INV_X1    g252(.A(G1gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(KEYINPUT16), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456));
  OAI221_X1 g255(.A(new_n455), .B1(new_n456), .B2(G8gat), .C1(new_n454), .C2(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(G8gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT21), .ZN(new_n461));
  INV_X1    g260(.A(G57gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(G64gat), .ZN(new_n463));
  INV_X1    g262(.A(G64gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(G57gat), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT94), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(G57gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(G64gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT94), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(KEYINPUT9), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G71gat), .A2(G78gat), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(G71gat), .A2(G78gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(KEYINPUT9), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n477), .A2(new_n472), .B1(new_n467), .B2(new_n468), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT95), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n481));
  AOI211_X1 g280(.A(new_n481), .B(new_n478), .C1(new_n471), .C2(new_n475), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n460), .B1(new_n461), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(G183gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n461), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G211gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n487), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G127gat), .B(G155gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(G231gat), .A2(G233gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n490), .B(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G134gat), .B(G162gat), .Z(new_n495));
  AOI21_X1  g294(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g300(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT15), .B(new_n499), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  OR3_X1    g308(.A1(new_n499), .A2(KEYINPUT91), .A3(KEYINPUT15), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n503), .A2(new_n506), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT15), .B1(new_n499), .B2(KEYINPUT91), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT17), .ZN(new_n515));
  XNOR2_X1  g314(.A(G99gat), .B(G106gat), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n516), .A2(KEYINPUT97), .ZN(new_n517));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518));
  INV_X1    g317(.A(G85gat), .ZN(new_n519));
  INV_X1    g318(.A(G92gat), .ZN(new_n520));
  AOI22_X1  g319(.A1(KEYINPUT8), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522));
  OAI22_X1  g321(.A1(new_n519), .A2(new_n520), .B1(new_n522), .B2(KEYINPUT96), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n524), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n516), .A2(KEYINPUT97), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n517), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n526), .A2(KEYINPUT97), .A3(new_n516), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT98), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n530), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n514), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n515), .A2(KEYINPUT98), .A3(new_n530), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT99), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI211_X1 g340(.A(KEYINPUT100), .B(new_n498), .C1(new_n538), .C2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n541), .B2(new_n538), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n538), .A2(new_n541), .A3(new_n498), .ZN(new_n544));
  INV_X1    g343(.A(new_n538), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n545), .B(new_n540), .C1(KEYINPUT100), .C2(new_n498), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n494), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n452), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n515), .A2(new_n460), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n514), .A2(new_n459), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n514), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n460), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT93), .A3(new_n552), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n551), .B(KEYINPUT13), .Z(new_n559));
  OR3_X1    g358(.A1(new_n514), .A2(new_n459), .A3(KEYINPUT93), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n551), .A4(new_n552), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G169gat), .B(G197gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT12), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n561), .A3(new_n569), .A4(new_n562), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT101), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n526), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n516), .ZN(new_n577));
  INV_X1    g376(.A(new_n516), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n526), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n577), .A2(new_n476), .A3(new_n479), .A4(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n483), .B2(new_n530), .ZN(new_n582));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n475), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n469), .B1(new_n467), .B2(new_n468), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n592), .B2(KEYINPUT9), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n481), .B1(new_n593), .B2(new_n478), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n476), .A2(KEYINPUT95), .A3(new_n479), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n535), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n594), .A2(new_n595), .A3(new_n530), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n580), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT102), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n599), .A2(new_n603), .A3(new_n600), .A4(new_n580), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n598), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n583), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n584), .B(new_n588), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n603), .B1(new_n582), .B2(new_n600), .ZN(new_n609));
  INV_X1    g408(.A(new_n604), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n597), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n583), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT103), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n614), .A3(new_n584), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n608), .B1(new_n615), .B2(new_n587), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n549), .A2(new_n574), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n430), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G1gat), .ZN(G1324gat));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n420), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT16), .B(G8gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n624), .A2(KEYINPUT42), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(G8gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(KEYINPUT42), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(G1325gat));
  NOR2_X1   g427(.A1(new_n410), .A2(new_n411), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(G15gat), .B1(new_n618), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n449), .ZN(new_n632));
  INV_X1    g431(.A(new_n450), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n618), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(G15gat), .B2(new_n636), .ZN(G1326gat));
  NAND2_X1  g436(.A1(new_n618), .A2(new_n379), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT43), .B(G22gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1327gat));
  INV_X1    g439(.A(new_n547), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n419), .B2(new_n451), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n574), .A2(new_n617), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n642), .A2(new_n643), .A3(new_n494), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(new_n504), .A3(new_n430), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n452), .A2(new_n547), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n642), .A2(KEYINPUT44), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n650), .A2(new_n643), .A3(new_n494), .A4(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(G29gat), .B1(new_n652), .B2(new_n276), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n653), .ZN(G1328gat));
  OR3_X1    g453(.A1(new_n652), .A2(KEYINPUT106), .A3(new_n349), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT106), .B1(new_n652), .B2(new_n349), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(G36gat), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n644), .A2(new_n505), .A3(new_n420), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT46), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(G1329gat));
  INV_X1    g459(.A(KEYINPUT47), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT107), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n630), .ZN(new_n663));
  INV_X1    g462(.A(G43gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT44), .B1(new_n452), .B2(new_n547), .ZN(new_n666));
  AOI211_X1 g465(.A(new_n649), .B(new_n641), .C1(new_n419), .C2(new_n451), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n668), .A2(new_n643), .A3(new_n635), .A4(new_n494), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n662), .B(new_n665), .C1(new_n669), .C2(new_n664), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n661), .A2(KEYINPUT107), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT108), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n670), .B(new_n672), .ZN(G1330gat));
  OAI21_X1  g472(.A(G50gat), .B1(new_n652), .B2(new_n380), .ZN(new_n674));
  INV_X1    g473(.A(G50gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n644), .A2(new_n675), .A3(new_n379), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT48), .B1(new_n676), .B2(KEYINPUT109), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1331gat));
  NOR3_X1   g478(.A1(new_n549), .A2(new_n573), .A3(new_n616), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n430), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT110), .B(G57gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1332gat));
  INV_X1    g482(.A(new_n680), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n349), .ZN(new_n685));
  NOR2_X1   g484(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n686));
  AND2_X1   g485(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n685), .B2(new_n686), .ZN(G1333gat));
  INV_X1    g488(.A(G71gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n680), .B2(new_n635), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n573), .A2(new_n616), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n452), .A2(new_n630), .A3(new_n548), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT111), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n379), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT112), .B(G78gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1335gat));
  NAND3_X1  g498(.A1(new_n668), .A2(new_n494), .A3(new_n692), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(new_n519), .A3(new_n276), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n642), .A2(new_n574), .A3(new_n494), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT51), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT51), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n642), .A2(new_n704), .A3(new_n574), .A4(new_n494), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n617), .A3(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(new_n276), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n701), .B1(new_n519), .B2(new_n707), .ZN(G1336gat));
  OAI21_X1  g507(.A(new_n520), .B1(new_n706), .B2(new_n349), .ZN(new_n709));
  AND4_X1   g508(.A1(new_n494), .A2(new_n650), .A3(new_n651), .A4(new_n692), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(G92gat), .A3(new_n420), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT52), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n709), .A2(new_n711), .A3(KEYINPUT52), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1337gat));
  OAI21_X1  g515(.A(G99gat), .B1(new_n700), .B2(new_n634), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n706), .A2(G99gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n629), .ZN(G1338gat));
  OAI21_X1  g518(.A(G106gat), .B1(new_n700), .B2(new_n380), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT53), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n617), .A3(new_n379), .A4(new_n705), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n720), .B(new_n721), .C1(G106gat), .C2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(G106gat), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n710), .B2(new_n379), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n722), .A2(G106gat), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT53), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(G1339gat));
  NAND2_X1  g527(.A1(new_n613), .A2(new_n614), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n588), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n605), .A2(new_n606), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n583), .B(new_n598), .C1(new_n602), .C2(new_n604), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT113), .B1(new_n734), .B2(KEYINPUT54), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737));
  NOR4_X1   g536(.A1(new_n732), .A2(new_n733), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n731), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n731), .B(KEYINPUT55), .C1(new_n735), .C2(new_n738), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n573), .A3(new_n607), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n568), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n572), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n617), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n547), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n741), .A2(new_n607), .A3(new_n742), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n748), .A2(KEYINPUT115), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(new_n544), .A3(new_n543), .A4(new_n546), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n494), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n494), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n758), .A2(new_n574), .A3(new_n616), .A4(new_n641), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT116), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n420), .A2(new_n276), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n630), .A2(new_n380), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n573), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G113gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n415), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n764), .A2(new_n773), .A3(new_n765), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(new_n227), .A3(new_n573), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(G1340gat));
  NAND3_X1  g576(.A1(new_n769), .A2(new_n617), .A3(new_n770), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G120gat), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n616), .A2(new_n226), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n774), .B2(new_n780), .ZN(G1341gat));
  AOI21_X1  g580(.A(G127gat), .B1(new_n775), .B2(new_n758), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n769), .A2(new_n770), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n758), .A2(G127gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(G1342gat));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n547), .A3(new_n770), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G134gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n774), .A2(new_n641), .ZN(new_n788));
  INV_X1    g587(.A(G134gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT56), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n790), .B2(KEYINPUT56), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n788), .A2(KEYINPUT118), .A3(new_n794), .A4(new_n789), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n787), .A2(new_n791), .A3(new_n793), .A4(new_n795), .ZN(G1343gat));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n761), .A2(new_n797), .A3(new_n379), .A4(new_n763), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT119), .B1(new_n748), .B2(new_n617), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n747), .A2(new_n616), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n547), .B1(new_n802), .B2(new_n743), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n494), .B1(new_n803), .B2(new_n756), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n759), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n379), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT57), .ZN(new_n807));
  NOR4_X1   g606(.A1(new_n632), .A2(new_n633), .A3(new_n276), .A4(new_n420), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n798), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n798), .A2(new_n807), .A3(KEYINPUT120), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n208), .B1(new_n813), .B2(new_n573), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n634), .A2(new_n379), .ZN(new_n815));
  NOR4_X1   g614(.A1(new_n766), .A2(G141gat), .A3(new_n574), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT58), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(KEYINPUT58), .ZN(new_n818));
  OAI21_X1  g617(.A(G141gat), .B1(new_n809), .B2(new_n574), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1344gat));
  NOR4_X1   g620(.A1(new_n766), .A2(G148gat), .A3(new_n616), .A4(new_n815), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT121), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n761), .A2(KEYINPUT57), .A3(new_n379), .A4(new_n763), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n826), .A3(new_n797), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n380), .B1(new_n804), .B2(new_n759), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT122), .B1(new_n828), .B2(KEYINPUT57), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n617), .A3(new_n808), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n210), .B1(new_n831), .B2(KEYINPUT123), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n830), .A2(new_n833), .A3(new_n617), .A4(new_n808), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n824), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n616), .B1(new_n811), .B2(new_n812), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n836), .A2(KEYINPUT59), .A3(new_n210), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n823), .B1(new_n835), .B2(new_n837), .ZN(G1345gat));
  NOR2_X1   g637(.A1(new_n766), .A2(new_n815), .ZN(new_n839));
  AOI21_X1  g638(.A(G155gat), .B1(new_n839), .B2(new_n758), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n494), .B1(new_n811), .B2(new_n812), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g641(.A(G162gat), .B1(new_n839), .B2(new_n547), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n641), .B1(new_n811), .B2(new_n812), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g644(.A1(new_n430), .A2(new_n349), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n630), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT125), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(KEYINPUT125), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n764), .A2(new_n380), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G169gat), .B1(new_n850), .B2(new_n574), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n764), .A2(new_n276), .A3(new_n773), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(G169gat), .A3(new_n349), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n855), .A2(new_n856), .A3(new_n573), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n855), .B2(new_n573), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(G1348gat));
  NOR3_X1   g658(.A1(new_n850), .A2(new_n290), .A3(new_n616), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n854), .A2(new_n349), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n617), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n862), .B2(new_n290), .ZN(G1349gat));
  NOR2_X1   g662(.A1(new_n494), .A2(new_n282), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G183gat), .B1(new_n850), .B2(new_n494), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(KEYINPUT127), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT60), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n865), .A2(KEYINPUT127), .A3(new_n866), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n850), .B2(new_n641), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT61), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n861), .A2(new_n286), .A3(new_n547), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1351gat));
  NAND2_X1  g674(.A1(new_n764), .A2(new_n276), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n349), .A3(new_n815), .ZN(new_n877));
  INV_X1    g676(.A(G197gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n573), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n634), .A2(new_n846), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n830), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(new_n573), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n879), .B1(new_n883), .B2(new_n878), .ZN(G1352gat));
  INV_X1    g683(.A(G204gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n877), .A2(new_n885), .A3(new_n617), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(KEYINPUT62), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n830), .A2(new_n617), .A3(new_n881), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G204gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(KEYINPUT62), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(G1353gat));
  NAND3_X1  g690(.A1(new_n877), .A2(new_n319), .A3(new_n758), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n830), .A2(new_n758), .A3(new_n881), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT63), .B1(new_n893), .B2(G211gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1354gat));
  AOI21_X1  g695(.A(G218gat), .B1(new_n877), .B2(new_n547), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n641), .A2(new_n321), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n882), .B2(new_n898), .ZN(G1355gat));
endmodule


