

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U556 ( .A(G2104), .B(KEYINPUT66), .Z(n523) );
  XNOR2_X2 U557 ( .A(n531), .B(n530), .ZN(n772) );
  XOR2_X2 U558 ( .A(KEYINPUT65), .B(n568), .Z(n661) );
  AND2_X1 U559 ( .A1(n548), .A2(n543), .ZN(n542) );
  NOR2_X1 U560 ( .A1(n803), .A2(n802), .ZN(n805) );
  NOR2_X2 U561 ( .A1(n611), .A2(n610), .ZN(n1018) );
  NOR2_X1 U562 ( .A1(G1966), .A2(n794), .ZN(n774) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n721) );
  NOR2_X1 U564 ( .A1(n720), .A2(n719), .ZN(n722) );
  OR2_X1 U565 ( .A1(n731), .A2(n715), .ZN(n716) );
  OR2_X1 U566 ( .A1(n728), .A2(n1006), .ZN(n727) );
  XNOR2_X1 U567 ( .A(n746), .B(n534), .ZN(n533) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n534) );
  XNOR2_X1 U569 ( .A(n536), .B(KEYINPUT31), .ZN(n535) );
  NOR2_X2 U570 ( .A1(n823), .A2(n825), .ZN(n731) );
  OR2_X1 U571 ( .A1(G164), .A2(G1384), .ZN(n823) );
  XNOR2_X1 U572 ( .A(G164), .B(G2078), .ZN(n968) );
  AND2_X1 U573 ( .A1(n606), .A2(n605), .ZN(n609) );
  XNOR2_X1 U574 ( .A(n607), .B(KEYINPUT13), .ZN(n608) );
  XNOR2_X1 U575 ( .A(KEYINPUT67), .B(KEYINPUT23), .ZN(n552) );
  INV_X1 U576 ( .A(n854), .ZN(n540) );
  NAND2_X1 U577 ( .A1(n528), .A2(n544), .ZN(n543) );
  NAND2_X1 U578 ( .A1(n854), .A2(n545), .ZN(n544) );
  NAND2_X1 U579 ( .A1(n547), .A2(n546), .ZN(n545) );
  INV_X1 U580 ( .A(KEYINPUT96), .ZN(n738) );
  NOR2_X1 U581 ( .A1(n774), .A2(n752), .ZN(n754) );
  INV_X1 U582 ( .A(KEYINPUT97), .ZN(n530) );
  INV_X1 U583 ( .A(n551), .ZN(n547) );
  INV_X1 U584 ( .A(n855), .ZN(n546) );
  NAND2_X1 U585 ( .A1(n523), .A2(n526), .ZN(n697) );
  XNOR2_X1 U586 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U587 ( .A(n557), .B(n556), .ZN(n711) );
  XNOR2_X1 U588 ( .A(n553), .B(n552), .ZN(n555) );
  NAND2_X1 U589 ( .A1(n541), .A2(n539), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n540), .A2(n855), .ZN(n539) );
  XNOR2_X1 U591 ( .A(n705), .B(n704), .ZN(n706) );
  AND2_X1 U592 ( .A1(n523), .A2(G2105), .ZN(n524) );
  OR2_X1 U593 ( .A1(G301), .A2(n756), .ZN(n525) );
  AND2_X1 U594 ( .A1(G2105), .A2(G126), .ZN(n526) );
  NAND2_X1 U595 ( .A1(G301), .A2(n756), .ZN(n527) );
  OR2_X1 U596 ( .A1(n854), .A2(n855), .ZN(n528) );
  NOR2_X1 U597 ( .A1(n791), .A2(n794), .ZN(n529) );
  NOR2_X2 U598 ( .A1(n707), .A2(n706), .ZN(G164) );
  XNOR2_X1 U599 ( .A(n925), .B(G164), .ZN(n926) );
  NAND2_X1 U600 ( .A1(n535), .A2(n532), .ZN(n531) );
  NAND2_X1 U601 ( .A1(n533), .A2(n525), .ZN(n532) );
  NAND2_X1 U602 ( .A1(n537), .A2(n527), .ZN(n536) );
  INV_X1 U603 ( .A(n757), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n542), .A2(n538), .ZN(G329) );
  INV_X1 U605 ( .A(n550), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n548) );
  AND2_X1 U607 ( .A1(n551), .A2(n855), .ZN(n549) );
  XNOR2_X1 U608 ( .A(n805), .B(n804), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n716), .B(KEYINPUT94), .ZN(n717) );
  BUF_X1 U610 ( .A(n731), .Z(n747) );
  INV_X1 U611 ( .A(n731), .ZN(n750) );
  AND2_X1 U612 ( .A1(n841), .A2(n840), .ZN(n551) );
  INV_X1 U613 ( .A(KEYINPUT27), .ZN(n732) );
  XNOR2_X1 U614 ( .A(n733), .B(n732), .ZN(n734) );
  INV_X1 U615 ( .A(KEYINPUT93), .ZN(n736) );
  XNOR2_X1 U616 ( .A(n737), .B(n736), .ZN(n742) );
  INV_X1 U617 ( .A(KEYINPUT30), .ZN(n753) );
  INV_X1 U618 ( .A(KEYINPUT32), .ZN(n768) );
  INV_X1 U619 ( .A(KEYINPUT102), .ZN(n800) );
  NOR2_X1 U620 ( .A1(n523), .A2(G2105), .ZN(n636) );
  INV_X1 U621 ( .A(KEYINPUT104), .ZN(n804) );
  INV_X1 U622 ( .A(KEYINPUT75), .ZN(n607) );
  NOR2_X1 U623 ( .A1(G651), .A2(n649), .ZN(n668) );
  INV_X1 U624 ( .A(KEYINPUT84), .ZN(n704) );
  NAND2_X1 U625 ( .A1(G101), .A2(n636), .ZN(n553) );
  NAND2_X1 U626 ( .A1(G125), .A2(n524), .ZN(n554) );
  NAND2_X1 U627 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U628 ( .A(KEYINPUT68), .ZN(n556) );
  NAND2_X1 U629 ( .A1(G2104), .A2(G2105), .ZN(n558) );
  XNOR2_X2 U630 ( .A(n558), .B(KEYINPUT69), .ZN(n915) );
  NAND2_X1 U631 ( .A1(G113), .A2(n915), .ZN(n563) );
  NOR2_X1 U632 ( .A1(G2105), .A2(G2104), .ZN(n559) );
  XNOR2_X1 U633 ( .A(n559), .B(KEYINPUT70), .ZN(n561) );
  XNOR2_X1 U634 ( .A(KEYINPUT71), .B(KEYINPUT17), .ZN(n560) );
  XNOR2_X1 U635 ( .A(n561), .B(n560), .ZN(n703) );
  NAND2_X1 U636 ( .A1(G137), .A2(n703), .ZN(n562) );
  AND2_X1 U637 ( .A1(n563), .A2(n562), .ZN(n709) );
  AND2_X1 U638 ( .A1(n711), .A2(n709), .ZN(G160) );
  INV_X1 U639 ( .A(G651), .ZN(n567) );
  NOR2_X1 U640 ( .A1(G543), .A2(n567), .ZN(n564) );
  XOR2_X1 U641 ( .A(KEYINPUT1), .B(n564), .Z(n665) );
  NAND2_X1 U642 ( .A1(G60), .A2(n665), .ZN(n566) );
  XOR2_X1 U643 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  NAND2_X1 U644 ( .A1(G47), .A2(n668), .ZN(n565) );
  NAND2_X1 U645 ( .A1(n566), .A2(n565), .ZN(n572) );
  NOR2_X2 U646 ( .A1(n649), .A2(n567), .ZN(n660) );
  NAND2_X1 U647 ( .A1(G72), .A2(n660), .ZN(n570) );
  NOR2_X1 U648 ( .A1(G651), .A2(G543), .ZN(n568) );
  NAND2_X1 U649 ( .A1(G85), .A2(n661), .ZN(n569) );
  NAND2_X1 U650 ( .A1(n570), .A2(n569), .ZN(n571) );
  OR2_X1 U651 ( .A1(n572), .A2(n571), .ZN(G290) );
  AND2_X1 U652 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U653 ( .A(G108), .ZN(G238) );
  INV_X1 U654 ( .A(G120), .ZN(G236) );
  INV_X1 U655 ( .A(G57), .ZN(G237) );
  INV_X1 U656 ( .A(G132), .ZN(G219) );
  INV_X1 U657 ( .A(G82), .ZN(G220) );
  NAND2_X1 U658 ( .A1(G64), .A2(n665), .ZN(n574) );
  NAND2_X1 U659 ( .A1(G52), .A2(n668), .ZN(n573) );
  NAND2_X1 U660 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U661 ( .A(KEYINPUT72), .B(n575), .ZN(n580) );
  NAND2_X1 U662 ( .A1(G77), .A2(n660), .ZN(n577) );
  NAND2_X1 U663 ( .A1(G90), .A2(n661), .ZN(n576) );
  NAND2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U665 ( .A(KEYINPUT9), .B(n578), .Z(n579) );
  NOR2_X1 U666 ( .A1(n580), .A2(n579), .ZN(G171) );
  NAND2_X1 U667 ( .A1(G62), .A2(n665), .ZN(n582) );
  NAND2_X1 U668 ( .A1(G50), .A2(n668), .ZN(n581) );
  NAND2_X1 U669 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U670 ( .A(KEYINPUT80), .B(n583), .Z(n587) );
  NAND2_X1 U671 ( .A1(G75), .A2(n660), .ZN(n585) );
  NAND2_X1 U672 ( .A1(G88), .A2(n661), .ZN(n584) );
  AND2_X1 U673 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U674 ( .A1(n587), .A2(n586), .ZN(G303) );
  NAND2_X1 U675 ( .A1(n661), .A2(G89), .ZN(n588) );
  XNOR2_X1 U676 ( .A(n588), .B(KEYINPUT4), .ZN(n590) );
  NAND2_X1 U677 ( .A1(G76), .A2(n660), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U679 ( .A(n591), .B(KEYINPUT5), .ZN(n596) );
  NAND2_X1 U680 ( .A1(G63), .A2(n665), .ZN(n593) );
  NAND2_X1 U681 ( .A1(G51), .A2(n668), .ZN(n592) );
  NAND2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U683 ( .A(KEYINPUT6), .B(n594), .Z(n595) );
  NAND2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U685 ( .A(n597), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U686 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U687 ( .A1(G7), .A2(G661), .ZN(n598) );
  XNOR2_X1 U688 ( .A(n598), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U689 ( .A(G567), .ZN(n692) );
  NOR2_X1 U690 ( .A1(n692), .A2(G223), .ZN(n599) );
  XNOR2_X1 U691 ( .A(n599), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U692 ( .A1(n665), .A2(G56), .ZN(n600) );
  XNOR2_X1 U693 ( .A(n600), .B(KEYINPUT14), .ZN(n602) );
  NAND2_X1 U694 ( .A1(G43), .A2(n668), .ZN(n601) );
  NAND2_X1 U695 ( .A1(n602), .A2(n601), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n661), .A2(G81), .ZN(n603) );
  XNOR2_X1 U697 ( .A(KEYINPUT12), .B(n603), .ZN(n606) );
  NAND2_X1 U698 ( .A1(n660), .A2(G68), .ZN(n604) );
  XNOR2_X1 U699 ( .A(n604), .B(KEYINPUT74), .ZN(n605) );
  NAND2_X1 U700 ( .A1(n1018), .A2(G860), .ZN(G153) );
  INV_X1 U701 ( .A(G171), .ZN(G301) );
  NAND2_X1 U702 ( .A1(G79), .A2(n660), .ZN(n613) );
  NAND2_X1 U703 ( .A1(G92), .A2(n661), .ZN(n612) );
  NAND2_X1 U704 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U705 ( .A1(G66), .A2(n665), .ZN(n615) );
  NAND2_X1 U706 ( .A1(G54), .A2(n668), .ZN(n614) );
  NAND2_X1 U707 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U708 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U709 ( .A(n618), .B(KEYINPUT15), .ZN(n1006) );
  INV_X1 U710 ( .A(G868), .ZN(n679) );
  NAND2_X1 U711 ( .A1(n1006), .A2(n679), .ZN(n619) );
  XNOR2_X1 U712 ( .A(n619), .B(KEYINPUT76), .ZN(n621) );
  NAND2_X1 U713 ( .A1(G868), .A2(G301), .ZN(n620) );
  NAND2_X1 U714 ( .A1(n621), .A2(n620), .ZN(G284) );
  NAND2_X1 U715 ( .A1(G78), .A2(n660), .ZN(n623) );
  NAND2_X1 U716 ( .A1(G91), .A2(n661), .ZN(n622) );
  NAND2_X1 U717 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U718 ( .A1(G65), .A2(n665), .ZN(n625) );
  NAND2_X1 U719 ( .A1(G53), .A2(n668), .ZN(n624) );
  NAND2_X1 U720 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U721 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U722 ( .A(n628), .B(KEYINPUT73), .ZN(G299) );
  NAND2_X1 U723 ( .A1(G286), .A2(G868), .ZN(n630) );
  NAND2_X1 U724 ( .A1(G299), .A2(n679), .ZN(n629) );
  NAND2_X1 U725 ( .A1(n630), .A2(n629), .ZN(G297) );
  INV_X1 U726 ( .A(G860), .ZN(n865) );
  NAND2_X1 U727 ( .A1(n865), .A2(G559), .ZN(n631) );
  INV_X1 U728 ( .A(n1006), .ZN(n930) );
  NAND2_X1 U729 ( .A1(n631), .A2(n930), .ZN(n632) );
  XNOR2_X1 U730 ( .A(n632), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U731 ( .A1(n930), .A2(G868), .ZN(n633) );
  NOR2_X1 U732 ( .A1(G559), .A2(n633), .ZN(n635) );
  AND2_X1 U733 ( .A1(n679), .A2(n1018), .ZN(n634) );
  NOR2_X1 U734 ( .A1(n635), .A2(n634), .ZN(G282) );
  BUF_X2 U735 ( .A(n636), .Z(n918) );
  NAND2_X1 U736 ( .A1(n918), .A2(G99), .ZN(n638) );
  BUF_X1 U737 ( .A(n703), .Z(n919) );
  NAND2_X1 U738 ( .A1(G135), .A2(n919), .ZN(n637) );
  NAND2_X1 U739 ( .A1(n638), .A2(n637), .ZN(n643) );
  NAND2_X1 U740 ( .A1(n524), .A2(G123), .ZN(n639) );
  XNOR2_X1 U741 ( .A(n639), .B(KEYINPUT18), .ZN(n641) );
  NAND2_X1 U742 ( .A1(G111), .A2(n915), .ZN(n640) );
  NAND2_X1 U743 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U744 ( .A1(n643), .A2(n642), .ZN(n953) );
  XNOR2_X1 U745 ( .A(n953), .B(G2096), .ZN(n645) );
  INV_X1 U746 ( .A(G2100), .ZN(n644) );
  NAND2_X1 U747 ( .A1(n645), .A2(n644), .ZN(G156) );
  NAND2_X1 U748 ( .A1(G49), .A2(n668), .ZN(n647) );
  NAND2_X1 U749 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U750 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U751 ( .A1(n665), .A2(n648), .ZN(n651) );
  NAND2_X1 U752 ( .A1(n649), .A2(G87), .ZN(n650) );
  NAND2_X1 U753 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U754 ( .A1(G61), .A2(n665), .ZN(n653) );
  NAND2_X1 U755 ( .A1(G48), .A2(n668), .ZN(n652) );
  NAND2_X1 U756 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U757 ( .A1(n660), .A2(G73), .ZN(n654) );
  XOR2_X1 U758 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U759 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U760 ( .A1(n661), .A2(G86), .ZN(n657) );
  NAND2_X1 U761 ( .A1(n658), .A2(n657), .ZN(G305) );
  NAND2_X1 U762 ( .A1(G559), .A2(n930), .ZN(n659) );
  XNOR2_X1 U763 ( .A(n659), .B(n1018), .ZN(n864) );
  NAND2_X1 U764 ( .A1(G80), .A2(n660), .ZN(n663) );
  NAND2_X1 U765 ( .A1(G93), .A2(n661), .ZN(n662) );
  NAND2_X1 U766 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U767 ( .A(n664), .B(KEYINPUT77), .ZN(n667) );
  NAND2_X1 U768 ( .A1(G67), .A2(n665), .ZN(n666) );
  NAND2_X1 U769 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U770 ( .A1(n668), .A2(G55), .ZN(n669) );
  XOR2_X1 U771 ( .A(KEYINPUT78), .B(n669), .Z(n670) );
  NOR2_X1 U772 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U773 ( .A(KEYINPUT79), .B(n672), .ZN(n866) );
  XNOR2_X1 U774 ( .A(G303), .B(n866), .ZN(n677) );
  XNOR2_X1 U775 ( .A(KEYINPUT19), .B(G299), .ZN(n673) );
  XNOR2_X1 U776 ( .A(n673), .B(G288), .ZN(n674) );
  XNOR2_X1 U777 ( .A(n674), .B(G290), .ZN(n675) );
  XNOR2_X1 U778 ( .A(n675), .B(G305), .ZN(n676) );
  XNOR2_X1 U779 ( .A(n677), .B(n676), .ZN(n929) );
  XNOR2_X1 U780 ( .A(n864), .B(n929), .ZN(n678) );
  NAND2_X1 U781 ( .A1(n678), .A2(G868), .ZN(n681) );
  NAND2_X1 U782 ( .A1(n679), .A2(n866), .ZN(n680) );
  NAND2_X1 U783 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U784 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U785 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U786 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U787 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U788 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U789 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U790 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U791 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U792 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U793 ( .A1(G96), .A2(n688), .ZN(n861) );
  NAND2_X1 U794 ( .A1(G2106), .A2(n861), .ZN(n689) );
  XNOR2_X1 U795 ( .A(n689), .B(KEYINPUT81), .ZN(n694) );
  NOR2_X1 U796 ( .A1(G236), .A2(G238), .ZN(n690) );
  NAND2_X1 U797 ( .A1(G69), .A2(n690), .ZN(n691) );
  NOR2_X1 U798 ( .A1(G237), .A2(n691), .ZN(n863) );
  NOR2_X1 U799 ( .A1(n692), .A2(n863), .ZN(n693) );
  NOR2_X1 U800 ( .A1(n694), .A2(n693), .ZN(G319) );
  INV_X1 U801 ( .A(G319), .ZN(n696) );
  NAND2_X1 U802 ( .A1(G483), .A2(G661), .ZN(n695) );
  NOR2_X1 U803 ( .A1(n696), .A2(n695), .ZN(n860) );
  NAND2_X1 U804 ( .A1(n860), .A2(G36), .ZN(G176) );
  INV_X1 U805 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U806 ( .A(n697), .B(KEYINPUT82), .ZN(n699) );
  NAND2_X1 U807 ( .A1(G114), .A2(n915), .ZN(n698) );
  NAND2_X1 U808 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U809 ( .A(n700), .B(KEYINPUT83), .ZN(n702) );
  NAND2_X1 U810 ( .A1(G102), .A2(n918), .ZN(n701) );
  NAND2_X1 U811 ( .A1(n702), .A2(n701), .ZN(n707) );
  NAND2_X1 U812 ( .A1(n703), .A2(G138), .ZN(n705) );
  NOR2_X1 U813 ( .A1(G1981), .A2(G305), .ZN(n708) );
  XNOR2_X1 U814 ( .A(KEYINPUT24), .B(n708), .ZN(n714) );
  AND2_X1 U815 ( .A1(G40), .A2(n709), .ZN(n710) );
  NAND2_X1 U816 ( .A1(n711), .A2(n710), .ZN(n825) );
  NAND2_X1 U817 ( .A1(n750), .A2(G8), .ZN(n712) );
  XOR2_X2 U818 ( .A(KEYINPUT91), .B(n712), .Z(n794) );
  INV_X1 U819 ( .A(n794), .ZN(n713) );
  NAND2_X1 U820 ( .A1(n714), .A2(n713), .ZN(n785) );
  INV_X1 U821 ( .A(G1341), .ZN(n715) );
  NAND2_X1 U822 ( .A1(n717), .A2(n1018), .ZN(n720) );
  NAND2_X1 U823 ( .A1(G1996), .A2(n731), .ZN(n718) );
  XOR2_X1 U824 ( .A(KEYINPUT26), .B(n718), .Z(n719) );
  XNOR2_X1 U825 ( .A(n722), .B(n721), .ZN(n728) );
  INV_X1 U826 ( .A(G1348), .ZN(n1029) );
  NOR2_X1 U827 ( .A1(n747), .A2(n1029), .ZN(n723) );
  XNOR2_X1 U828 ( .A(n723), .B(KEYINPUT95), .ZN(n725) );
  NAND2_X1 U829 ( .A1(n747), .A2(G2067), .ZN(n724) );
  NAND2_X1 U830 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U831 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U832 ( .A1(n728), .A2(n1006), .ZN(n729) );
  NAND2_X1 U833 ( .A1(n730), .A2(n729), .ZN(n741) );
  NAND2_X1 U834 ( .A1(G1956), .A2(n750), .ZN(n735) );
  NAND2_X1 U835 ( .A1(n731), .A2(G2072), .ZN(n733) );
  NAND2_X1 U836 ( .A1(n735), .A2(n734), .ZN(n737) );
  NOR2_X1 U837 ( .A1(G299), .A2(n742), .ZN(n739) );
  XNOR2_X1 U838 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U839 ( .A1(n741), .A2(n740), .ZN(n745) );
  NAND2_X1 U840 ( .A1(G299), .A2(n742), .ZN(n743) );
  XNOR2_X1 U841 ( .A(n743), .B(KEYINPUT28), .ZN(n744) );
  NAND2_X1 U842 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U843 ( .A1(G1961), .A2(n750), .ZN(n749) );
  XOR2_X1 U844 ( .A(G2078), .B(KEYINPUT25), .Z(n985) );
  NAND2_X1 U845 ( .A1(n747), .A2(n985), .ZN(n748) );
  NAND2_X1 U846 ( .A1(n749), .A2(n748), .ZN(n756) );
  NOR2_X1 U847 ( .A1(G2084), .A2(n750), .ZN(n751) );
  XOR2_X1 U848 ( .A(KEYINPUT92), .B(n751), .Z(n770) );
  NAND2_X1 U849 ( .A1(G8), .A2(n770), .ZN(n752) );
  XNOR2_X1 U850 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U851 ( .A1(G168), .A2(n755), .ZN(n757) );
  AND2_X1 U852 ( .A1(G286), .A2(G8), .ZN(n758) );
  NAND2_X1 U853 ( .A1(n772), .A2(n758), .ZN(n767) );
  INV_X1 U854 ( .A(G8), .ZN(n765) );
  NOR2_X1 U855 ( .A1(G2090), .A2(n750), .ZN(n759) );
  XNOR2_X1 U856 ( .A(n759), .B(KEYINPUT98), .ZN(n761) );
  NOR2_X1 U857 ( .A1(n794), .A2(G1971), .ZN(n760) );
  NOR2_X1 U858 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U859 ( .A1(n762), .A2(G303), .ZN(n763) );
  XOR2_X1 U860 ( .A(KEYINPUT99), .B(n763), .Z(n764) );
  OR2_X1 U861 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U862 ( .A1(n767), .A2(n766), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n769), .B(n768), .ZN(n778) );
  INV_X1 U864 ( .A(n770), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n771), .A2(G8), .ZN(n776) );
  INV_X1 U866 ( .A(n772), .ZN(n773) );
  NOR2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n779), .B(KEYINPUT100), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G8), .A2(G166), .ZN(n780) );
  NOR2_X1 U872 ( .A1(G2090), .A2(n780), .ZN(n781) );
  XNOR2_X1 U873 ( .A(KEYINPUT103), .B(n781), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n789), .A2(n782), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n783), .A2(n794), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n803) );
  NOR2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n792) );
  NOR2_X1 U878 ( .A1(G1971), .A2(G303), .ZN(n786) );
  NOR2_X1 U879 ( .A1(n792), .A2(n786), .ZN(n1003) );
  INV_X1 U880 ( .A(KEYINPUT33), .ZN(n787) );
  AND2_X1 U881 ( .A1(n1003), .A2(n787), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G288), .A2(G1976), .ZN(n790) );
  XOR2_X1 U884 ( .A(KEYINPUT101), .B(n790), .Z(n1002) );
  INV_X1 U885 ( .A(n1002), .ZN(n791) );
  NOR2_X1 U886 ( .A1(KEYINPUT33), .A2(n529), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n792), .A2(KEYINPUT33), .ZN(n793) );
  NOR2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U890 ( .A(G1981), .B(G305), .Z(n1014) );
  AND2_X1 U891 ( .A1(n797), .A2(n1014), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n801) );
  XNOR2_X1 U893 ( .A(n801), .B(n800), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G129), .A2(n524), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G141), .A2(n919), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n918), .A2(G105), .ZN(n808) );
  XOR2_X1 U898 ( .A(KEYINPUT38), .B(n808), .Z(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n915), .A2(G117), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n912) );
  NAND2_X1 U902 ( .A1(G1996), .A2(n912), .ZN(n822) );
  NAND2_X1 U903 ( .A1(n918), .A2(G95), .ZN(n814) );
  NAND2_X1 U904 ( .A1(G131), .A2(n919), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT88), .B(n815), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G107), .A2(n915), .ZN(n816) );
  XNOR2_X1 U908 ( .A(KEYINPUT87), .B(n816), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U910 ( .A1(n524), .A2(G119), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n897) );
  NAND2_X1 U912 ( .A1(G1991), .A2(n897), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n963) );
  INV_X1 U914 ( .A(n823), .ZN(n824) );
  NOR2_X1 U915 ( .A1(n824), .A2(n825), .ZN(n852) );
  NAND2_X1 U916 ( .A1(n963), .A2(n852), .ZN(n826) );
  XNOR2_X1 U917 ( .A(n826), .B(KEYINPUT89), .ZN(n844) );
  INV_X1 U918 ( .A(n844), .ZN(n838) );
  NAND2_X1 U919 ( .A1(n918), .A2(G104), .ZN(n827) );
  XOR2_X1 U920 ( .A(KEYINPUT85), .B(n827), .Z(n829) );
  NAND2_X1 U921 ( .A1(G140), .A2(n919), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(KEYINPUT34), .B(n830), .ZN(n835) );
  NAND2_X1 U924 ( .A1(G128), .A2(n524), .ZN(n832) );
  NAND2_X1 U925 ( .A1(G116), .A2(n915), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U927 ( .A(n833), .B(KEYINPUT35), .Z(n834) );
  NOR2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U929 ( .A(KEYINPUT36), .B(n836), .Z(n837) );
  XOR2_X1 U930 ( .A(KEYINPUT86), .B(n837), .Z(n898) );
  XNOR2_X1 U931 ( .A(G2067), .B(KEYINPUT37), .ZN(n850) );
  NOR2_X1 U932 ( .A1(n898), .A2(n850), .ZN(n964) );
  NAND2_X1 U933 ( .A1(n852), .A2(n964), .ZN(n848) );
  NAND2_X1 U934 ( .A1(n838), .A2(n848), .ZN(n839) );
  XOR2_X1 U935 ( .A(KEYINPUT90), .B(n839), .Z(n841) );
  XNOR2_X1 U936 ( .A(G1986), .B(G290), .ZN(n1005) );
  NAND2_X1 U937 ( .A1(n1005), .A2(n852), .ZN(n840) );
  NOR2_X1 U938 ( .A1(G1996), .A2(n912), .ZN(n958) );
  NOR2_X1 U939 ( .A1(G1986), .A2(G290), .ZN(n842) );
  NOR2_X1 U940 ( .A1(G1991), .A2(n897), .ZN(n954) );
  NOR2_X1 U941 ( .A1(n842), .A2(n954), .ZN(n843) );
  NOR2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U943 ( .A1(n958), .A2(n845), .ZN(n846) );
  XOR2_X1 U944 ( .A(n846), .B(KEYINPUT105), .Z(n847) );
  XNOR2_X1 U945 ( .A(n847), .B(KEYINPUT39), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n851) );
  NAND2_X1 U947 ( .A1(n898), .A2(n850), .ZN(n955) );
  NAND2_X1 U948 ( .A1(n851), .A2(n955), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U950 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n855) );
  INV_X1 U951 ( .A(G223), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n856), .A2(G2106), .ZN(n857) );
  XOR2_X1 U953 ( .A(KEYINPUT109), .B(n857), .Z(G217) );
  AND2_X1 U954 ( .A1(G15), .A2(G2), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G661), .A2(n858), .ZN(G259) );
  NAND2_X1 U956 ( .A1(G3), .A2(G1), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(G188) );
  INV_X1 U959 ( .A(G96), .ZN(G221) );
  INV_X1 U960 ( .A(n861), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(G261) );
  INV_X1 U962 ( .A(G261), .ZN(G325) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n867) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(G145) );
  XNOR2_X1 U965 ( .A(G1991), .B(G2474), .ZN(n877) );
  XOR2_X1 U966 ( .A(G1956), .B(G1961), .Z(n869) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1986), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U969 ( .A(G1976), .B(G1981), .Z(n871) );
  XNOR2_X1 U970 ( .A(G1966), .B(G1971), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U972 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(G229) );
  XOR2_X1 U976 ( .A(G2100), .B(G2096), .Z(n879) );
  XNOR2_X1 U977 ( .A(KEYINPUT42), .B(G2678), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U979 ( .A(KEYINPUT43), .B(G2090), .Z(n881) );
  XNOR2_X1 U980 ( .A(G2067), .B(G2072), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U983 ( .A(G2078), .B(G2084), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(G227) );
  NAND2_X1 U985 ( .A1(G112), .A2(n915), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G100), .A2(n918), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n894) );
  NAND2_X1 U988 ( .A1(G136), .A2(n919), .ZN(n888) );
  XNOR2_X1 U989 ( .A(KEYINPUT111), .B(n888), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n524), .A2(G124), .ZN(n889) );
  XOR2_X1 U991 ( .A(KEYINPUT44), .B(n889), .Z(n890) );
  NOR2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(KEYINPUT112), .B(n892), .Z(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(G162) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n896) );
  XNOR2_X1 U996 ( .A(n953), .B(KEYINPUT113), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n897), .B(G162), .ZN(n900) );
  XNOR2_X1 U999 ( .A(G160), .B(n898), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n914) );
  NAND2_X1 U1002 ( .A1(G127), .A2(n524), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(G115), .A2(n915), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n905), .B(KEYINPUT47), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(n918), .A2(G103), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(G139), .A2(n919), .ZN(n906) );
  NAND2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1009 ( .A(KEYINPUT114), .B(n908), .Z(n909) );
  NAND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n911), .B(KEYINPUT115), .ZN(n967) );
  XNOR2_X1 U1012 ( .A(n912), .B(n967), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n927) );
  NAND2_X1 U1014 ( .A1(G130), .A2(n524), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(G118), .A2(n915), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n924) );
  NAND2_X1 U1017 ( .A1(n918), .A2(G106), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(G142), .A2(n919), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1020 ( .A(KEYINPUT45), .B(n922), .Z(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n928), .ZN(G395) );
  XOR2_X1 U1024 ( .A(n929), .B(G286), .Z(n932) );
  XNOR2_X1 U1025 ( .A(G171), .B(n930), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(n932), .B(n931), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(n933), .B(n1018), .ZN(n934) );
  NOR2_X1 U1028 ( .A1(G37), .A2(n934), .ZN(G397) );
  XNOR2_X1 U1029 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(G229), .A2(G227), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(n936), .B(n935), .ZN(n949) );
  XNOR2_X1 U1032 ( .A(KEYINPUT108), .B(G2438), .ZN(n946) );
  XOR2_X1 U1033 ( .A(G2435), .B(G2454), .Z(n938) );
  XNOR2_X1 U1034 ( .A(G2446), .B(KEYINPUT107), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n938), .B(n937), .ZN(n942) );
  XOR2_X1 U1036 ( .A(G2451), .B(G2427), .Z(n940) );
  XNOR2_X1 U1037 ( .A(G1348), .B(G1341), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(n940), .B(n939), .ZN(n941) );
  XOR2_X1 U1039 ( .A(n942), .B(n941), .Z(n944) );
  XNOR2_X1 U1040 ( .A(G2443), .B(G2430), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(n944), .B(n943), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(n946), .B(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n947), .A2(G14), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(G319), .A2(n952), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(G395), .A2(G397), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(G225) );
  INV_X1 U1048 ( .A(G225), .ZN(G308) );
  INV_X1 U1049 ( .A(G69), .ZN(G235) );
  INV_X1 U1050 ( .A(n952), .ZN(G401) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G162), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n957), .B(KEYINPUT117), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT51), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n975) );
  XNOR2_X1 U1058 ( .A(G160), .B(G2084), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(G2072), .B(n967), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n968), .B(KEYINPUT118), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n971), .B(KEYINPUT50), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT52), .B(n976), .ZN(n977) );
  XOR2_X1 U1068 ( .A(KEYINPUT119), .B(n977), .Z(n978) );
  NOR2_X1 U1069 ( .A1(KEYINPUT55), .A2(n978), .ZN(n979) );
  XOR2_X1 U1070 ( .A(KEYINPUT120), .B(n979), .Z(n980) );
  NAND2_X1 U1071 ( .A1(G29), .A2(n980), .ZN(n1058) );
  XOR2_X1 U1072 ( .A(G34), .B(KEYINPUT123), .Z(n982) );
  XNOR2_X1 U1073 ( .A(G2084), .B(KEYINPUT54), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n982), .B(n981), .ZN(n999) );
  XNOR2_X1 U1075 ( .A(G2090), .B(G35), .ZN(n996) );
  XNOR2_X1 U1076 ( .A(G2067), .B(G26), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G32), .B(G1996), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n985), .B(G27), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G33), .B(G2072), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(KEYINPUT121), .B(n990), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n991), .A2(G28), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(G25), .B(G1991), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(KEYINPUT53), .B(n994), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1089 ( .A(KEYINPUT122), .B(n997), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1091 ( .A(KEYINPUT55), .B(n1000), .Z(n1001) );
  NOR2_X1 U1092 ( .A1(G29), .A2(n1001), .ZN(n1056) );
  XNOR2_X1 U1093 ( .A(G16), .B(KEYINPUT56), .ZN(n1026) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1024) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G1348), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT125), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G171), .B(G1961), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(G1971), .A2(G303), .ZN(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(G1956), .B(G299), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1022) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G168), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(n1016), .B(KEYINPUT57), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT124), .B(n1017), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(n1018), .B(G1341), .ZN(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1052) );
  INV_X1 U1113 ( .A(G16), .ZN(n1050) );
  XNOR2_X1 U1114 ( .A(G1966), .B(G21), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(G5), .B(G1961), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1039) );
  XNOR2_X1 U1117 ( .A(G4), .B(KEYINPUT59), .ZN(n1030) );
  XNOR2_X1 U1118 ( .A(n1030), .B(n1029), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(G20), .B(G1956), .ZN(n1031) );
  NOR2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1036) );
  XNOR2_X1 U1121 ( .A(G1341), .B(G19), .ZN(n1034) );
  XNOR2_X1 U1122 ( .A(G1981), .B(G6), .ZN(n1033) );
  NOR2_X1 U1123 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1124 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1125 ( .A(KEYINPUT60), .B(n1037), .Z(n1038) );
  NAND2_X1 U1126 ( .A1(n1039), .A2(n1038), .ZN(n1047) );
  XNOR2_X1 U1127 ( .A(G1986), .B(G24), .ZN(n1041) );
  XNOR2_X1 U1128 ( .A(G1971), .B(G22), .ZN(n1040) );
  NOR2_X1 U1129 ( .A1(n1041), .A2(n1040), .ZN(n1044) );
  XOR2_X1 U1130 ( .A(G1976), .B(KEYINPUT126), .Z(n1042) );
  XNOR2_X1 U1131 ( .A(G23), .B(n1042), .ZN(n1043) );
  NAND2_X1 U1132 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1133 ( .A(KEYINPUT58), .B(n1045), .ZN(n1046) );
  NOR2_X1 U1134 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XNOR2_X1 U1135 ( .A(KEYINPUT61), .B(n1048), .ZN(n1049) );
  NAND2_X1 U1136 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  NAND2_X1 U1137 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  XNOR2_X1 U1138 ( .A(KEYINPUT127), .B(n1053), .ZN(n1054) );
  NAND2_X1 U1139 ( .A1(n1054), .A2(G11), .ZN(n1055) );
  NOR2_X1 U1140 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
  NAND2_X1 U1141 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  XOR2_X1 U1142 ( .A(KEYINPUT62), .B(n1059), .Z(G311) );
  INV_X1 U1143 ( .A(G311), .ZN(G150) );
endmodule

