//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n566, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT69), .Z(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT70), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(new_n462), .A3(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(new_n470), .B1(KEYINPUT3), .B2(new_n460), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n467), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n471), .A2(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT72), .Z(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n459), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n460), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT73), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n480), .A2(G136), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(new_n468), .A2(new_n470), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(G126), .A3(new_n461), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n459), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n459), .A2(G102), .A3(G2104), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n459), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n488), .A2(new_n459), .A3(new_n461), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n491), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT75), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT74), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT74), .A2(G651), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n500), .B(KEYINPUT6), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT74), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT75), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n501), .A2(new_n502), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n511), .A2(G50), .B1(G75), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n511), .A2(G88), .B1(G62), .B2(new_n512), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(new_n510), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n521), .B1(new_n512), .B2(new_n504), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n514), .B1(new_n522), .B2(new_n503), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n511), .A2(G89), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n517), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G168));
  AOI21_X1  g108(.A(new_n518), .B1(new_n522), .B2(new_n503), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G90), .ZN(new_n535));
  INV_X1    g110(.A(new_n512), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT77), .B(G52), .Z(new_n539));
  AOI21_X1  g114(.A(new_n538), .B1(new_n525), .B2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(new_n525), .A2(G43), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT78), .B(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n518), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n534), .A2(new_n542), .B1(new_n512), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT79), .Z(G176));
  XOR2_X1   g127(.A(KEYINPUT80), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(G188));
  AOI22_X1  g131(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n506), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n534), .B2(G91), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n523), .A2(KEYINPUT9), .A3(G53), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n532), .B(new_n566), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n523), .A2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n534), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND3_X1  g147(.A1(new_n511), .A2(G86), .A3(new_n517), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n517), .A2(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n536), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT82), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n525), .A2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT83), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(new_n512), .B1(G85), .B2(new_n534), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(new_n525), .A2(G54), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n511), .A2(G92), .A3(new_n517), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n506), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(G171), .ZN(G321));
  XOR2_X1   g174(.A(G321), .B(KEYINPUT84), .Z(G284));
  NAND2_X1  g175(.A1(G299), .A2(new_n597), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n532), .B(KEYINPUT81), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n597), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n597), .ZN(G280));
  AND3_X1   g179(.A1(new_n591), .A2(new_n595), .A3(new_n593), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n547), .A2(new_n597), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n606), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT85), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n610), .B2(new_n597), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g187(.A1(new_n476), .A2(G123), .B1(G135), .B2(new_n480), .ZN(new_n613));
  NOR2_X1   g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT13), .Z(new_n621));
  NOR2_X1   g196(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n622));
  AND2_X1   g197(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n617), .B(new_n624), .C1(new_n622), .C2(new_n621), .ZN(G156));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  OAI21_X1  g203(.A(KEYINPUT14), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT88), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT89), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(G14), .ZN(G401));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n642), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n644), .A2(new_n645), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT18), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n649), .B(new_n652), .Z(G227));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n665), .C1(new_n663), .C2(new_n662), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n666), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT90), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G19), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n548), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G1341), .Z(new_n677));
  INV_X1    g252(.A(KEYINPUT23), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(G20), .ZN(new_n679));
  AOI22_X1  g254(.A1(G299), .A2(G16), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G1956), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(G171), .A2(G16), .ZN(new_n684));
  OR2_X1    g259(.A1(G5), .A2(G16), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(G1961), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n463), .A3(G127), .ZN(new_n687));
  INV_X1    g262(.A(G115), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n460), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n480), .A2(G139), .B1(G2105), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT25), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G33), .B(new_n693), .S(G29), .Z(new_n694));
  NOR2_X1   g269(.A1(KEYINPUT24), .A2(G34), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(KEYINPUT24), .A2(G34), .ZN(new_n697));
  AOI21_X1  g272(.A(G29), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI211_X1 g277(.A(new_n700), .B(new_n702), .C1(G160), .C2(G29), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n694), .A2(G2072), .B1(new_n703), .B2(G2084), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT26), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n476), .B2(G129), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n480), .A2(G141), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT97), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n707), .A2(KEYINPUT97), .A3(new_n708), .A4(new_n709), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(G29), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT27), .B(G1996), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G32), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n683), .A2(new_n686), .A3(new_n704), .A4(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n694), .A2(G2072), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(G27), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n717), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2078), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G26), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(KEYINPUT28), .ZN(new_n728));
  INV_X1    g303(.A(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G140), .ZN(new_n730));
  NOR2_X1   g305(.A1(G104), .A2(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT93), .Z(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n733));
  OAI22_X1  g308(.A1(new_n479), .A2(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n476), .B2(G128), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n729), .B1(new_n736), .B2(new_n717), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n728), .B1(new_n737), .B2(KEYINPUT28), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT95), .B(G2067), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT30), .B(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  NAND2_X1  g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n741), .A2(new_n717), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n616), .B2(new_n717), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT98), .Z(new_n746));
  NAND3_X1  g321(.A1(new_n725), .A2(new_n740), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n674), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n605), .B2(new_n674), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n716), .B1(new_n714), .B2(new_n718), .ZN(new_n752));
  AOI21_X1  g327(.A(G1961), .B1(new_n684), .B2(new_n685), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n703), .A2(G2084), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT99), .A4(new_n754), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n747), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n674), .B1(new_n581), .B2(new_n583), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT32), .B(G1981), .Z(new_n762));
  NOR2_X1   g337(.A1(G6), .A2(G16), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G22), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT91), .B1(new_n765), .B2(G16), .ZN(new_n766));
  OR3_X1    g341(.A1(new_n765), .A2(KEYINPUT91), .A3(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(G166), .C2(new_n674), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(G1971), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n762), .B1(new_n761), .B2(new_n763), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(G1971), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n764), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G288), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G16), .B2(G23), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT33), .B(G1976), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  OR3_X1    g352(.A1(new_n772), .A2(KEYINPUT34), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT34), .B1(new_n772), .B2(new_n777), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n674), .A2(G24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n589), .B2(new_n674), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n476), .A2(G119), .B1(G131), .B2(new_n480), .ZN(new_n784));
  NOR2_X1   g359(.A1(G95), .A2(G2105), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G25), .B(new_n787), .S(G29), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT35), .B(G1991), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n783), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n780), .A2(KEYINPUT92), .A3(KEYINPUT36), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n792), .A2(new_n778), .A3(new_n779), .ZN(new_n794));
  NAND2_X1  g369(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n795));
  OR2_X1    g370(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AND4_X1   g372(.A1(new_n677), .A2(new_n760), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n674), .A2(G21), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G168), .B2(new_n674), .ZN(new_n800));
  INV_X1    g375(.A(G1966), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n717), .A2(G35), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n717), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2090), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n798), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(G311));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT101), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n798), .A2(new_n811), .A3(new_n802), .A4(new_n807), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(G150));
  NAND2_X1  g388(.A1(new_n525), .A2(G55), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(new_n536), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n534), .A2(G93), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n548), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT103), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n820), .B1(new_n822), .B2(new_n547), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n596), .A2(new_n606), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT39), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n823), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT104), .B(G860), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT105), .Z(new_n831));
  INV_X1    g406(.A(new_n822), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n829), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(G145));
  XNOR2_X1  g411(.A(new_n787), .B(new_n710), .ZN(new_n837));
  INV_X1    g412(.A(new_n736), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n693), .A2(new_n711), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G164), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n616), .B(new_n473), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n486), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n480), .A2(G142), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT107), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n476), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n620), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n845), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n843), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n842), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g434(.A(G166), .B(G288), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(G305), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n589), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT42), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n610), .B(new_n823), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n596), .B(G299), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT41), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n865), .B2(new_n864), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT108), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n863), .A2(new_n868), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n597), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n870), .A2(new_n872), .B1(new_n597), .B2(new_n822), .ZN(G295));
  AOI22_X1  g448(.A1(new_n870), .A2(new_n872), .B1(new_n597), .B2(new_n822), .ZN(G331));
  NAND2_X1  g449(.A1(new_n822), .A2(new_n547), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n819), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n532), .A2(G171), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(G286), .B2(G171), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n602), .A2(G301), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n823), .B1(new_n880), .B2(new_n877), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n879), .A2(new_n881), .A3(new_n866), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n865), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  OAI211_X1 g458(.A(KEYINPUT109), .B(new_n862), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n861), .A2(new_n589), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n861), .A2(new_n589), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT109), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n879), .A2(new_n881), .A3(new_n866), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n879), .A2(new_n881), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n865), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n884), .A2(new_n890), .A3(new_n857), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n882), .A2(new_n883), .A3(new_n862), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n862), .B1(new_n882), .B2(new_n883), .ZN(new_n895));
  AND4_X1   g470(.A1(KEYINPUT43), .A2(new_n894), .A3(new_n857), .A4(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT44), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n891), .A2(KEYINPUT43), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n894), .A2(new_n892), .A3(new_n857), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n897), .A2(new_n902), .ZN(G397));
  INV_X1    g478(.A(G1384), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n491), .B2(new_n498), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(G40), .B(new_n467), .C1(new_n472), .C2(G2105), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G1996), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT46), .Z(new_n912));
  XNOR2_X1  g487(.A(new_n736), .B(G2067), .ZN(new_n913));
  INV_X1    g488(.A(new_n710), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT47), .ZN(new_n917));
  INV_X1    g492(.A(new_n909), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n710), .A2(G1996), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n712), .A2(new_n713), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n910), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n922), .A2(new_n789), .A3(new_n787), .ZN(new_n923));
  INV_X1    g498(.A(G2067), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n736), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n918), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(G290), .A2(G1986), .A3(new_n918), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT48), .ZN(new_n928));
  INV_X1    g503(.A(new_n922), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n787), .B(new_n789), .Z(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n931), .B2(new_n909), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n917), .A2(new_n926), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(KEYINPUT45), .B(new_n904), .C1(new_n491), .C2(new_n498), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n907), .ZN(new_n937));
  INV_X1    g512(.A(G2078), .ZN(new_n938));
  INV_X1    g513(.A(new_n908), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n905), .A2(new_n935), .A3(new_n906), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT53), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n905), .A2(KEYINPUT50), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n489), .A2(new_n490), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G2105), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n495), .A2(new_n497), .ZN(new_n949));
  AOI21_X1  g524(.A(G1384), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n908), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n905), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n946), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1961), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n907), .A2(new_n934), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n908), .B(KEYINPUT122), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n942), .A2(G2078), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(KEYINPUT123), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT123), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n908), .B(KEYINPUT122), .Z(new_n963));
  NAND3_X1  g538(.A1(new_n907), .A2(new_n934), .A3(new_n960), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n943), .A2(new_n956), .A3(new_n961), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G171), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND4_X1   g544(.A1(new_n907), .A2(new_n939), .A3(new_n934), .A4(new_n960), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n954), .B2(new_n955), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n943), .A3(G301), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(KEYINPUT54), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(KEYINPUT125), .A3(G171), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n976));
  INV_X1    g551(.A(G1971), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(G2090), .B2(new_n954), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT55), .B(G8), .C1(new_n515), .C2(new_n519), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(G166), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n979), .A2(G8), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n573), .A2(new_n574), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n573), .B2(new_n574), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(new_n577), .ZN(new_n991));
  INV_X1    g566(.A(G1981), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT115), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n580), .A2(new_n992), .ZN(new_n994));
  INV_X1    g569(.A(new_n990), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n573), .A2(new_n574), .A3(new_n988), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n578), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(G1981), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n994), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n905), .A2(new_n908), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n983), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n993), .A2(new_n999), .A3(KEYINPUT49), .A4(new_n994), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n939), .B1(new_n905), .B2(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(new_n944), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1008), .A2(new_n1009), .A3(G2090), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n977), .B2(new_n976), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1007), .B1(new_n1011), .B2(new_n983), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1004), .B1(new_n1013), .B2(G288), .ZN(new_n1014));
  NAND2_X1  g589(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OR3_X1    g591(.A1(new_n773), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AND4_X1   g594(.A1(new_n987), .A2(new_n1006), .A3(new_n1012), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n801), .B1(new_n957), .B2(new_n908), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n954), .B2(G2084), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n532), .A2(G8), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n1024), .C1(KEYINPUT120), .C2(KEYINPUT51), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT51), .B1(new_n1024), .B2(KEYINPUT120), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(G8), .C1(new_n1022), .C2(new_n532), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1025), .B(new_n1027), .C1(G168), .C2(new_n1023), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n975), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT56), .B(G2072), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n682), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT117), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1035), .A3(new_n1032), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n562), .A2(new_n563), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n559), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  NAND2_X1  g616(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1042));
  NAND3_X1  g617(.A1(G299), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1034), .A2(new_n1036), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n954), .A2(new_n750), .B1(new_n924), .B2(new_n1003), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n596), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1044), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n1032), .A3(new_n1031), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1046), .A2(KEYINPUT60), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1046), .A2(KEYINPUT60), .A3(new_n596), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n596), .B1(new_n1046), .B2(KEYINPUT60), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT61), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1048), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1033), .A2(new_n1044), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n937), .A2(new_n910), .A3(new_n939), .A4(new_n940), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n905), .B2(new_n908), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n547), .B(new_n1059), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n548), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1054), .A2(new_n1058), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1055), .B1(new_n1057), .B2(KEYINPUT119), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1049), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1069), .A2(new_n1045), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1050), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n971), .A2(new_n943), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(G171), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n966), .A2(G171), .ZN(new_n1077));
  AOI211_X1 g652(.A(KEYINPUT121), .B(G301), .C1(new_n971), .C2(new_n943), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT124), .B1(new_n1079), .B2(KEYINPUT54), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1076), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1081), .B(new_n1082), .C1(new_n1085), .C2(new_n1077), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1029), .A2(new_n1073), .A3(new_n1080), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT126), .ZN(new_n1088));
  INV_X1    g663(.A(new_n954), .ZN(new_n1089));
  INV_X1    g664(.A(G2090), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1089), .A2(new_n1090), .B1(new_n976), .B2(new_n977), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1007), .B1(new_n1091), .B2(new_n983), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1023), .A2(G286), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(new_n1006), .A3(new_n1093), .A4(new_n1019), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1094), .A2(KEYINPUT63), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1006), .A2(new_n1019), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1012), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1096), .B1(new_n1098), .B2(new_n987), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1004), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1006), .A2(new_n1013), .A3(new_n773), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(new_n994), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1095), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1087), .A2(new_n1088), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1088), .B1(new_n1087), .B2(new_n1103), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1107));
  AND4_X1   g682(.A1(new_n1085), .A2(new_n1106), .A3(new_n1020), .A4(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1104), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n931), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n589), .B(G1986), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n918), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n933), .B1(new_n1109), .B2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g688(.A(G227), .ZN(new_n1115));
  NAND2_X1  g689(.A1(new_n1115), .A2(G319), .ZN(new_n1116));
  OR2_X1    g690(.A1(new_n1116), .A2(KEYINPUT127), .ZN(new_n1117));
  AND2_X1   g691(.A1(new_n858), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g692(.A(G229), .ZN(new_n1119));
  AOI21_X1  g693(.A(G401), .B1(KEYINPUT127), .B2(new_n1116), .ZN(new_n1120));
  NAND4_X1  g694(.A1(new_n900), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(G225));
  INV_X1    g695(.A(G225), .ZN(G308));
endmodule


