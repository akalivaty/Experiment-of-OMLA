//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT70), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n205), .C1(new_n203), .C2(KEYINPUT70), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(KEYINPUT28), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n218), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(KEYINPUT28), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n217), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(KEYINPUT24), .Z(new_n226));
  NOR2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n220), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT25), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n233), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n235), .B(new_n236), .C1(new_n226), .C2(new_n227), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n224), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT71), .ZN(new_n239));
  AND2_X1   g038(.A1(G226gat), .A2(G233gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(KEYINPUT29), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n213), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n238), .A2(KEYINPUT71), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n238), .A2(KEYINPUT71), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n242), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n224), .A2(new_n234), .A3(new_n237), .A4(new_n240), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n247), .A2(new_n213), .A3(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT72), .B(G64gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G92gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  NOR2_X1   g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT73), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n250), .A2(new_n256), .A3(KEYINPUT30), .A4(new_n254), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT30), .B(new_n254), .C1(new_n244), .C2(new_n249), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT73), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n255), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n250), .A2(new_n254), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT30), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G148gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G141gat), .ZN(new_n269));
  INV_X1    g068(.A(G141gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G148gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275));
  INV_X1    g074(.A(G155gat), .ZN(new_n276));
  INV_X1    g075(.A(G162gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(KEYINPUT2), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n269), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n269), .B2(new_n271), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT75), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n278), .A2(new_n288), .A3(new_n275), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n279), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n293));
  OAI21_X1  g092(.A(G120gat), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G120gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G113gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G113gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n299), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n287), .A2(new_n289), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n270), .A2(G148gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n268), .A2(G141gat), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT74), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n269), .A2(new_n271), .A3(new_n281), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n308), .A2(new_n313), .A3(new_n280), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n314), .A2(new_n279), .B1(new_n305), .B2(new_n300), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n267), .B1(new_n307), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT5), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n291), .A2(new_n306), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT1), .B1(new_n294), .B2(new_n296), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n304), .B1(new_n320), .B2(new_n299), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(new_n314), .A3(new_n279), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n266), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT78), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n325), .A3(KEYINPUT77), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n291), .A2(new_n306), .A3(KEYINPUT4), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n278), .A2(new_n275), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n272), .B2(new_n273), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n311), .A2(new_n312), .B1(KEYINPUT2), .B2(new_n275), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n308), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n332), .B2(new_n321), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n266), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(new_n279), .C1(new_n284), .C2(new_n290), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n306), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n335), .A2(KEYINPUT76), .A3(new_n306), .A4(new_n337), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n334), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n326), .A2(KEYINPUT5), .A3(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G1gat), .B(G29gat), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G85gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n318), .A2(new_n325), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n340), .A2(new_n341), .ZN(new_n350));
  INV_X1    g149(.A(new_n334), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n343), .A2(new_n347), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT6), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n347), .B1(new_n343), .B2(new_n353), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT6), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n354), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n265), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n361));
  INV_X1    g160(.A(G22gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n337), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n213), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT79), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n367), .B(new_n213), .C1(new_n337), .C2(new_n363), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n210), .A2(new_n203), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n210), .B2(new_n203), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n336), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n291), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n366), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT80), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n364), .A2(new_n365), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n367), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n364), .A2(KEYINPUT79), .A3(new_n365), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n372), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n375), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n211), .B2(new_n212), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n291), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n376), .A3(new_n378), .A4(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n362), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n390), .ZN(new_n392));
  AOI211_X1 g191(.A(G22gat), .B(new_n392), .C1(new_n377), .C2(new_n383), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n361), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n374), .A2(KEYINPUT80), .A3(new_n376), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n382), .B1(new_n381), .B2(new_n375), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G22gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n384), .A2(new_n362), .A3(new_n390), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(KEYINPUT82), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT31), .B(G50gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n394), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n238), .A2(new_n321), .ZN(new_n406));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n407), .B(KEYINPUT64), .Z(new_n408));
  NAND4_X1  g207(.A1(new_n224), .A2(new_n234), .A3(new_n237), .A4(new_n306), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT32), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n410), .B(KEYINPUT32), .C1(new_n412), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT68), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n409), .ZN(new_n422));
  INV_X1    g221(.A(new_n408), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT34), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(KEYINPUT67), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n422), .B2(new_n423), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n421), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n422), .A2(new_n423), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n426), .B(KEYINPUT68), .C1(new_n432), .C2(new_n428), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n420), .A2(new_n430), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n420), .A2(new_n430), .A3(new_n433), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n427), .A2(new_n429), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT69), .B1(new_n420), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n398), .A2(KEYINPUT82), .A3(new_n399), .A4(new_n403), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n405), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT86), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n405), .A2(new_n443), .A3(new_n440), .A4(new_n439), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(KEYINPUT35), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(KEYINPUT36), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n420), .A2(new_n437), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n420), .A2(new_n437), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n405), .A2(new_n440), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n360), .B1(new_n445), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n453), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n452), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n343), .A2(new_n353), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n343), .A2(KEYINPUT84), .A3(new_n353), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n347), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n357), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT37), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n244), .B2(new_n249), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n241), .A2(new_n213), .A3(new_n243), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n247), .A2(new_n248), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n466), .B(KEYINPUT37), .C1(new_n467), .C2(new_n213), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  INV_X1    g268(.A(new_n254), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n465), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n463), .A2(new_n355), .A3(new_n261), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT85), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n250), .A2(new_n464), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n465), .A2(new_n470), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT38), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n462), .A2(new_n357), .B1(KEYINPUT6), .B2(new_n354), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n261), .A4(new_n471), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n327), .ZN(new_n481));
  INV_X1    g280(.A(new_n333), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n266), .B1(new_n350), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT39), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n347), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n307), .A2(new_n315), .A3(new_n267), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n488), .B2(new_n485), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n489), .A2(new_n490), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n264), .A3(new_n494), .A4(new_n462), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n457), .B1(new_n480), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n264), .A2(new_n477), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n453), .A2(new_n449), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT35), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n455), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501));
  XOR2_X1   g300(.A(G15gat), .B(G22gat), .Z(new_n502));
  INV_X1    g301(.A(G1gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(G1gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n510), .A3(G8gat), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n504), .B(new_n509), .C1(new_n505), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G43gat), .B(G50gat), .Z(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT87), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT14), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n521), .B(new_n524), .C1(new_n519), .C2(new_n520), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n517), .A2(new_n518), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n520), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n501), .B1(new_n516), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n514), .B(KEYINPUT89), .ZN(new_n532));
  INV_X1    g331(.A(new_n530), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT91), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n530), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n511), .A2(new_n513), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n527), .A2(new_n542), .A3(new_n529), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n527), .B2(new_n529), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(new_n535), .A3(new_n538), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT11), .B(G169gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n545), .A2(new_n535), .A3(KEYINPUT18), .A4(new_n538), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n540), .A2(new_n548), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n554), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n561), .A3(new_n554), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n548), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n553), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n557), .A2(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n202), .B1(new_n500), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n480), .A2(new_n495), .ZN(new_n567));
  INV_X1    g366(.A(new_n457), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n499), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n445), .A2(new_n454), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n360), .ZN(new_n572));
  INV_X1    g371(.A(new_n565), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n532), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT97), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n587), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n578), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT96), .ZN(new_n598));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  NAND3_X1  g399(.A1(new_n590), .A2(new_n594), .A3(new_n578), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n600), .ZN(new_n603));
  INV_X1    g402(.A(new_n601), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(new_n595), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT7), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n608), .B(KEYINPUT98), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G99gat), .B(G106gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT99), .B(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n616), .A2(new_n617), .B1(KEYINPUT8), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n611), .A2(new_n614), .A3(new_n615), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT101), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n611), .A2(new_n614), .A3(new_n619), .ZN(new_n624));
  INV_X1    g423(.A(new_n615), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n620), .A2(new_n621), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n621), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n623), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n544), .B2(new_n543), .ZN(new_n632));
  NAND3_X1  g431(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n632), .B(new_n633), .C1(new_n631), .C2(new_n533), .ZN(new_n634));
  XOR2_X1   g433(.A(G190gat), .B(G218gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G134gat), .B(G162gat), .Z(new_n637));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n636), .B(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n607), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n585), .A2(KEYINPUT10), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n585), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n631), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n622), .A2(new_n583), .A3(new_n626), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n622), .A2(KEYINPUT102), .A3(new_n583), .A4(new_n626), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n644), .B1(new_n652), .B2(KEYINPUT10), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n655), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(G176gat), .B(G204gat), .Z(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n657), .A2(KEYINPUT104), .A3(new_n658), .A4(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n566), .A2(new_n574), .A3(new_n642), .A4(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n359), .A2(KEYINPUT105), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n359), .A2(KEYINPUT105), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n503), .ZN(G1324gat));
  NOR2_X1   g475(.A1(new_n671), .A2(new_n265), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n512), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n679), .B(G8gat), .C1(new_n671), .C2(new_n265), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT106), .B(KEYINPUT16), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G8gat), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n677), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n677), .B2(new_n685), .ZN(new_n687));
  OAI22_X1  g486(.A1(new_n680), .A2(new_n682), .B1(new_n686), .B2(new_n687), .ZN(G1325gat));
  INV_X1    g487(.A(new_n671), .ZN(new_n689));
  INV_X1    g488(.A(new_n449), .ZN(new_n690));
  AOI21_X1  g489(.A(G15gat), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n452), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT108), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n689), .B2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n671), .A2(new_n456), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  OAI21_X1  g497(.A(KEYINPUT44), .B1(new_n500), .B2(new_n640), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n569), .A2(new_n570), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n700), .B(new_n641), .C1(new_n701), .C2(new_n455), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n565), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n674), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n606), .B(KEYINPUT109), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n669), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G29gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT45), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n566), .A2(new_n574), .A3(new_n607), .A4(new_n670), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n640), .ZN(new_n711));
  INV_X1    g510(.A(G29gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n704), .ZN(new_n713));
  MUX2_X1   g512(.A(KEYINPUT45), .B(new_n709), .S(new_n713), .Z(G1328gat));
  INV_X1    g513(.A(new_n711), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n265), .A2(G36gat), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n703), .A2(new_n706), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n718), .B2(new_n265), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT46), .B1(new_n715), .B2(new_n716), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(G1329gat));
  NAND4_X1  g520(.A1(new_n703), .A2(G43gat), .A3(new_n692), .A4(new_n706), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n710), .A2(new_n640), .A3(new_n449), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(G43gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n724), .B(new_n726), .ZN(G1330gat));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n728), .A3(new_n453), .ZN(new_n729));
  OAI21_X1  g528(.A(G50gat), .B1(new_n718), .B2(new_n456), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n729), .B2(new_n730), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1331gat));
  NAND3_X1  g533(.A1(new_n606), .A2(new_n640), .A3(new_n565), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n670), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT111), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n572), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n572), .A2(new_n737), .A3(KEYINPUT112), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n704), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n745));
  INV_X1    g544(.A(G64gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n264), .B(KEYINPUT113), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n740), .A2(new_n741), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n751), .A2(KEYINPUT114), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(KEYINPUT114), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n745), .A2(new_n746), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1333gat));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n690), .ZN(new_n758));
  INV_X1    g557(.A(G71gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n742), .A2(G71gat), .A3(new_n692), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT50), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n764), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n742), .A2(new_n453), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n699), .A2(new_n702), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n573), .A2(new_n606), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n669), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n769), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g573(.A(KEYINPUT115), .B(new_n772), .C1(new_n699), .C2(new_n702), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n704), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n616), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n572), .A2(new_n641), .A3(new_n771), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT51), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n572), .A2(new_n780), .A3(new_n641), .A4(new_n771), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n669), .A3(new_n704), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n777), .B1(new_n616), .B2(new_n783), .ZN(G1336gat));
  NOR2_X1   g583(.A1(new_n749), .A2(G92gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n779), .A2(new_n669), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n787));
  AOI211_X1 g586(.A(new_n749), .B(new_n772), .C1(new_n699), .C2(new_n702), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n617), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n702), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n700), .B1(new_n572), .B2(new_n641), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n773), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G92gat), .B1(new_n794), .B2(new_n749), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n795), .A2(KEYINPUT117), .A3(new_n786), .A4(new_n787), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  INV_X1    g597(.A(new_n786), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n264), .B1(new_n774), .B2(new_n775), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(G92gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(G1337gat));
  NOR2_X1   g601(.A1(new_n774), .A2(new_n775), .ZN(new_n803));
  OAI21_X1  g602(.A(G99gat), .B1(new_n803), .B2(new_n452), .ZN(new_n804));
  INV_X1    g603(.A(G99gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n782), .A2(new_n805), .A3(new_n669), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n449), .B2(new_n806), .ZN(G1338gat));
  NOR2_X1   g606(.A1(new_n456), .A2(G106gat), .ZN(new_n808));
  AND4_X1   g607(.A1(new_n669), .A2(new_n779), .A3(new_n781), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n794), .B2(new_n456), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n453), .B1(new_n774), .B2(new_n775), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n813), .B2(G106gat), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(new_n705), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n644), .B(new_n655), .C1(new_n652), .C2(KEYINPUT10), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n653), .A2(new_n656), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n662), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n657), .A2(KEYINPUT118), .A3(KEYINPUT54), .A4(new_n818), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n821), .A2(new_n824), .A3(KEYINPUT55), .A4(new_n825), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n828), .A2(new_n573), .A3(new_n668), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n558), .A2(new_n557), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n536), .A2(new_n539), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n538), .B1(new_n545), .B2(new_n535), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n552), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n669), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n641), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n829), .A2(new_n668), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n834), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n640), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n838), .A2(new_n828), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n817), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n735), .A2(new_n669), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n674), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n442), .A2(new_n444), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(new_n749), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(new_n573), .C1(new_n293), .C2(new_n292), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n498), .A3(new_n749), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n565), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1340gat));
  NAND3_X1  g651(.A1(new_n848), .A2(new_n295), .A3(new_n669), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n850), .B2(new_n670), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1341gat));
  INV_X1    g654(.A(G127gat), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n850), .A2(new_n856), .A3(new_n817), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n848), .A2(new_n606), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n856), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n640), .A2(new_n264), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n847), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT56), .Z(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n850), .B2(new_n640), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1343gat));
  XOR2_X1   g664(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n866));
  NAND2_X1  g665(.A1(new_n826), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n573), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n835), .B1(new_n868), .B2(new_n837), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n640), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n838), .A2(new_n828), .A3(new_n840), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n606), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n453), .B1(new_n872), .B2(new_n843), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n704), .A2(new_n749), .A3(new_n452), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n456), .B1(new_n842), .B2(new_n844), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n874), .A2(new_n573), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT121), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n875), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n882), .A2(new_n883), .A3(new_n573), .A4(new_n879), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(G141gat), .A3(new_n884), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n454), .B(new_n674), .C1(new_n842), .C2(new_n844), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n749), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n270), .A3(new_n573), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n880), .A2(G141gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(G1344gat));
  NAND3_X1  g694(.A1(new_n888), .A2(new_n268), .A3(new_n669), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n882), .A2(new_n879), .ZN(new_n897));
  AOI211_X1 g696(.A(KEYINPUT59), .B(new_n268), .C1(new_n897), .C2(new_n669), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n839), .B1(new_n668), .B2(new_n663), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n565), .B1(new_n826), .B2(new_n866), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n838), .B2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n900), .B(new_n871), .C1(new_n903), .C2(new_n641), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n607), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n900), .B1(new_n870), .B2(new_n871), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n844), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n878), .A3(new_n453), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n842), .A2(new_n844), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n456), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n908), .A2(new_n669), .A3(new_n876), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n899), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n896), .B1(new_n898), .B2(new_n912), .ZN(G1345gat));
  AOI21_X1  g712(.A(G155gat), .B1(new_n888), .B2(new_n606), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n817), .A2(new_n276), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n897), .B2(new_n915), .ZN(G1346gat));
  NAND3_X1  g715(.A1(new_n886), .A2(new_n277), .A3(new_n861), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n882), .A2(new_n641), .A3(new_n879), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n277), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n917), .C1(new_n918), .C2(new_n277), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1347gat));
  AOI21_X1  g722(.A(new_n704), .B1(new_n842), .B2(new_n844), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(new_n846), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n750), .ZN(new_n926));
  INV_X1    g725(.A(G169gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(new_n573), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n264), .A3(new_n498), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n565), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n926), .B2(new_n669), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n929), .A2(new_n670), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(G176gat), .B2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n926), .A2(new_n606), .A3(new_n214), .ZN(new_n935));
  AND2_X1   g734(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n929), .B2(new_n817), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n936), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n926), .A2(new_n215), .A3(new_n641), .ZN(new_n941));
  OAI21_X1  g740(.A(G190gat), .B1(new_n929), .B2(new_n640), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  NAND2_X1  g744(.A1(new_n674), .A2(new_n452), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n264), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n908), .A2(new_n910), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(G197gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n565), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n946), .A2(new_n749), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n877), .A2(new_n573), .A3(new_n953), .ZN(new_n954));
  AOI22_X1  g753(.A1(new_n950), .A2(new_n952), .B1(new_n951), .B2(new_n954), .ZN(G1352gat));
  NAND4_X1  g754(.A1(new_n908), .A2(new_n669), .A3(new_n910), .A4(new_n949), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G204gat), .ZN(new_n957));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n877), .A2(new_n958), .A3(new_n669), .A4(new_n953), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n957), .A2(KEYINPUT126), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1353gat));
  NAND4_X1  g765(.A1(new_n877), .A2(new_n207), .A3(new_n606), .A4(new_n953), .ZN(new_n967));
  INV_X1    g766(.A(new_n948), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n908), .A2(new_n968), .A3(new_n606), .A4(new_n910), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  NOR2_X1   g771(.A1(new_n640), .A2(new_n208), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT127), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n877), .A2(new_n641), .A3(new_n953), .ZN(new_n975));
  AOI22_X1  g774(.A1(new_n950), .A2(new_n974), .B1(new_n208), .B2(new_n975), .ZN(G1355gat));
endmodule


