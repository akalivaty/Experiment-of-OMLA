//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n462), .A2(G2105), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT68), .Z(G160));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT70), .Z(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(G136), .B2(new_n471), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n468), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n478), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n460), .B2(new_n461), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n461), .C2(new_n460), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT71), .A2(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(G2105), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n485), .A2(G126), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n514), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n509), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n511), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n524), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  AOI22_X1  g103(.A1(new_n517), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n520), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n534));
  AND3_X1   g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n517), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n512), .A2(KEYINPUT73), .A3(new_n514), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(G543), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n537), .B1(new_n543), .B2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  AOI22_X1  g121(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n511), .B1(new_n522), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n541), .B(KEYINPUT74), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n549), .B1(new_n550), .B2(G52), .ZN(G171));
  NAND2_X1  g126(.A1(new_n550), .A2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n532), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n512), .A2(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n555), .A2(G651), .B1(G81), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n532), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(G91), .B2(new_n556), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n539), .A2(G53), .A3(G543), .A4(new_n540), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n509), .B1(new_n517), .B2(new_n538), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n572), .A2(new_n573), .A3(G53), .A4(new_n540), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n571), .B1(new_n570), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n568), .B1(new_n575), .B2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G52), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n543), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT77), .B1(new_n579), .B2(new_n549), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n581));
  NAND2_X1  g156(.A1(G171), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G301));
  NAND4_X1  g159(.A1(new_n539), .A2(G49), .A3(G543), .A4(new_n540), .ZN(new_n585));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n519), .A2(new_n586), .A3(new_n520), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n556), .A2(G87), .B1(G651), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n532), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G48), .B2(new_n515), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n556), .A2(G86), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n596), .A2(new_n511), .B1(new_n522), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n543), .B2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(new_n550), .A2(G54), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n522), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n532), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n605), .A2(new_n606), .B1(G651), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n583), .B2(G868), .ZN(G284));
  XNOR2_X1  g188(.A(G284), .B(KEYINPUT78), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(G286), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(G299), .B(KEYINPUT79), .Z(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(G297));
  AOI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(G280));
  AND2_X1   g194(.A1(new_n602), .A2(new_n610), .ZN(new_n620));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n624), .A2(KEYINPUT80), .A3(new_n615), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT80), .B1(new_n624), .B2(new_n615), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n625), .B(new_n626), .C1(G868), .C2(new_n559), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n471), .A2(G135), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n630), .A2(KEYINPUT82), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(KEYINPUT82), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G111), .B2(new_n468), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n629), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n488), .B2(G123), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT83), .Z(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT84), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n649), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(KEYINPUT17), .ZN(new_n670));
  INV_X1    g245(.A(new_n665), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n664), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT87), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n664), .A2(new_n666), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n664), .A2(new_n670), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n669), .B(new_n673), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G4), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n620), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT93), .B(G1348), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G19), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT94), .Z(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n559), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1341), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(G21), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G168), .B2(new_n702), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1966), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT24), .B(G34), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT97), .ZN(new_n714));
  INV_X1    g289(.A(G160), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2084), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G35), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G162), .B2(G29), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT29), .B(G2090), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(G164), .A2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G27), .B2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(G28), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n712), .B1(new_n726), .B2(G28), .ZN(new_n728));
  AND2_X1   g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n723), .B2(new_n724), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n712), .A2(G32), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n488), .A2(G129), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n735), .B(new_n737), .C1(G141), .C2(new_n471), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n712), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT27), .B(G1996), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n721), .A2(new_n725), .A3(new_n732), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n741), .A2(new_n743), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n719), .A2(new_n720), .B1(new_n636), .B2(new_n712), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AND4_X1   g323(.A1(new_n701), .A2(new_n710), .A3(new_n717), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n702), .A2(G20), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT23), .ZN(new_n751));
  INV_X1    g326(.A(G299), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n702), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT99), .Z(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT98), .B(G1956), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G33), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT95), .Z(new_n759));
  NAND3_X1  g334(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n479), .A2(new_n468), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n479), .A2(G127), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n468), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n759), .B1(new_n770), .B2(new_n712), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2072), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n702), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n702), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G1961), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(G1961), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n712), .A2(G26), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT28), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n471), .A2(G140), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n468), .A2(G116), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  INV_X1    g357(.A(G128), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n780), .B1(new_n781), .B2(new_n782), .C1(new_n487), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n779), .B1(new_n784), .B2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n773), .A2(new_n776), .A3(new_n777), .A4(new_n787), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n749), .A2(new_n757), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n755), .A2(new_n756), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n712), .A2(G25), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n471), .A2(G131), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n468), .A2(G107), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n795));
  INV_X1    g370(.A(G119), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n793), .B1(new_n794), .B2(new_n795), .C1(new_n487), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT88), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n792), .B1(new_n799), .B2(new_n712), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT35), .B(G1991), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT89), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n800), .A2(new_n803), .ZN(new_n805));
  INV_X1    g380(.A(G1986), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n598), .B1(new_n550), .B2(G47), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n702), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n702), .B2(G24), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n806), .B2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n702), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n702), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G1971), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(G1971), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n702), .A2(G6), .ZN(new_n818));
  INV_X1    g393(.A(G305), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n702), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT32), .B(G1981), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n815), .B1(new_n814), .B2(new_n816), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G23), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n826));
  NAND2_X1  g401(.A1(G288), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT90), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n825), .B1(new_n830), .B2(G16), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT33), .B(G1976), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n823), .A2(new_n824), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT34), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n811), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(KEYINPUT92), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n840), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n791), .B1(new_n842), .B2(new_n843), .ZN(G311));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n790), .B(new_n789), .C1(new_n845), .C2(new_n841), .ZN(G150));
  NAND2_X1  g421(.A1(new_n620), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(new_n511), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n556), .A2(G93), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n850), .B(new_n851), .C1(new_n543), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n558), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n851), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n550), .B2(G55), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n552), .A3(new_n557), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n848), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  AOI21_X1  g435(.A(G860), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n853), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n797), .B(KEYINPUT101), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n639), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n488), .A2(G130), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  INV_X1    g444(.A(G118), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(G2105), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n471), .B2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n867), .A2(new_n874), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n739), .B(new_n784), .ZN(new_n879));
  INV_X1    g454(.A(new_n497), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n496), .B1(new_n479), .B2(new_n493), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n503), .A2(new_n505), .ZN(new_n883));
  INV_X1    g458(.A(G126), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n480), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT100), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n498), .A2(new_n506), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n879), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n769), .ZN(new_n891));
  INV_X1    g466(.A(new_n889), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n879), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n770), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n877), .A2(new_n878), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n875), .A2(new_n876), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n891), .B(new_n894), .C1(new_n897), .C2(KEYINPUT102), .ZN(new_n898));
  XNOR2_X1  g473(.A(G160), .B(new_n490), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n636), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n897), .B2(new_n895), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n895), .B2(new_n897), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g481(.A1(new_n752), .A2(new_n620), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n611), .A2(G299), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n908), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n858), .B(new_n623), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n624), .B(new_n858), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(G290), .A2(G166), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n807), .A2(G303), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n830), .A2(G305), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n829), .A2(new_n819), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n926), .A3(new_n929), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n934), .A2(KEYINPUT104), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n916), .A2(new_n922), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n924), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n935), .B1(new_n924), .B2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g516(.A(new_n940), .B1(G868), .B2(new_n856), .ZN(G331));
  INV_X1    g517(.A(new_n858), .ZN(new_n943));
  AOI21_X1  g518(.A(G286), .B1(new_n580), .B2(new_n582), .ZN(new_n944));
  NOR2_X1   g519(.A1(G168), .A2(G171), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n583), .A2(G168), .ZN(new_n947));
  INV_X1    g522(.A(new_n945), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n858), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n909), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n858), .A3(new_n948), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n919), .A4(new_n920), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n933), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n954), .A2(new_n902), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n953), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n933), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT105), .B1(new_n931), .B2(new_n932), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT43), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n954), .A2(new_n902), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n958), .A2(new_n959), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n910), .B(new_n913), .C1(new_n946), .C2(new_n949), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n953), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n955), .B2(new_n960), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n962), .A2(new_n965), .A3(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n593), .A2(KEYINPUT111), .A3(new_n974), .A4(new_n594), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n591), .B1(new_n519), .B2(new_n520), .ZN(new_n976));
  INV_X1    g551(.A(new_n590), .ZN(new_n977));
  OAI21_X1  g552(.A(G651), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n515), .A2(G48), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n594), .A2(new_n978), .A3(new_n979), .A4(new_n974), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n975), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT112), .B(G86), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n978), .B(new_n979), .C1(new_n522), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G1981), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(KEYINPUT49), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  INV_X1    g563(.A(G137), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n469), .B1(new_n764), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n479), .A2(G125), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n468), .B1(new_n991), .B2(new_n465), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT106), .B(G40), .Z(new_n993));
  NOR3_X1   g568(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n498), .B2(new_n506), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n988), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n987), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n975), .A2(new_n982), .B1(new_n985), .B2(G1981), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT113), .B1(new_n998), .B2(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n983), .A2(new_n986), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n997), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n827), .A2(G1976), .A3(new_n828), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n996), .A3(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1005), .A2(new_n996), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT114), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1003), .A2(new_n999), .ZN(new_n1013));
  INV_X1    g588(.A(new_n997), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1011), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT55), .Z(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n886), .A2(new_n888), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT107), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n886), .A2(new_n1026), .A3(new_n888), .A4(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n994), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1971), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n993), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n467), .A2(new_n472), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n882), .B2(new_n885), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT109), .B(G2090), .Z(new_n1037));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n995), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n995), .B2(new_n1039), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1036), .B(new_n1037), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(G8), .B(new_n1021), .C1(new_n1031), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1029), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1042), .B1(new_n1047), .B2(G1971), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1048), .A2(KEYINPUT110), .A3(G8), .A4(new_n1021), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1019), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1004), .A2(G1976), .A3(G288), .ZN(new_n1051));
  INV_X1    g626(.A(new_n983), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n996), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1037), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n995), .A2(new_n1039), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1036), .A2(new_n1057), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1047), .A2(G1971), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1021), .B1(new_n1059), .B2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2084), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1036), .B(new_n1063), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1064));
  INV_X1    g639(.A(G1966), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n507), .A2(new_n1023), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1029), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(G8), .A3(G168), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT115), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1055), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1021), .B1(new_n1048), .B2(G8), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n1072), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1055), .A2(new_n1019), .A3(new_n1070), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1054), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n724), .A2(KEYINPUT53), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1029), .A2(new_n1066), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1057), .A2(KEYINPUT108), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n995), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1961), .B1(new_n1082), .B2(new_n1036), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1047), .A2(new_n724), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1079), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1086), .A2(G301), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1068), .A2(G8), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G168), .A2(new_n988), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(KEYINPUT51), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1064), .A2(KEYINPUT122), .A3(new_n1067), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT122), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(G286), .ZN(new_n1094));
  NAND2_X1  g669(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1087), .B1(new_n1098), .B2(KEYINPUT62), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1055), .A2(new_n1062), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT124), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1055), .A2(new_n1102), .A3(new_n1062), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1096), .A2(new_n1104), .A3(new_n1097), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1099), .A2(new_n1101), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT45), .B1(new_n892), .B2(new_n1034), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G40), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT123), .B1(new_n473), .B2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n473), .A2(KEYINPUT123), .A3(new_n1110), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(new_n1078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1109), .A2(new_n1028), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1083), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1107), .A2(new_n1114), .A3(G301), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1086), .B2(G301), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1117), .A2(new_n1118), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1107), .A2(new_n1115), .A3(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G171), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT125), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1123), .A3(G171), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1118), .B1(new_n1086), .B2(G301), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1101), .A2(new_n1119), .A3(new_n1126), .A4(new_n1103), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT116), .B(G1956), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1047), .A2(new_n1129), .B1(new_n1058), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT57), .B(new_n568), .C1(new_n575), .C2(new_n576), .ZN(new_n1132));
  INV_X1    g707(.A(new_n568), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n570), .B2(new_n574), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT117), .B1(new_n1134), .B2(KEYINPUT57), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n570), .A2(new_n574), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1136), .B(new_n1137), .C1(new_n1138), .C2(new_n1133), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1132), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1131), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1047), .A2(new_n1129), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1058), .A2(new_n1130), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1142), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1128), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n994), .B1(new_n995), .B2(new_n1039), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n994), .A2(new_n995), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1147), .A2(G1348), .B1(G2067), .B2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1149), .A2(KEYINPUT60), .A3(new_n611), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n620), .ZN(new_n1151));
  OAI221_X1 g726(.A(new_n611), .B1(G2067), .B2(new_n1148), .C1(new_n1147), .C2(G1348), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1150), .B1(new_n1153), .B2(KEYINPUT60), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1140), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1132), .A2(new_n1135), .A3(KEYINPUT118), .A4(new_n1139), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1131), .A2(new_n1140), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(KEYINPUT61), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(G1996), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1047), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT58), .B(G1341), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n994), .B2(new_n995), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n559), .B(new_n1163), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1047), .B2(new_n1164), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1162), .B(KEYINPUT59), .C1(new_n1169), .C2(new_n558), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1145), .A2(new_n1154), .A3(new_n1161), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1159), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT119), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1159), .B(KEYINPUT119), .C1(new_n1144), .C2(new_n1151), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1172), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1077), .B(new_n1106), .C1(new_n1127), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1108), .A2(new_n994), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(G1996), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n739), .B(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n784), .B(new_n786), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n797), .B(new_n803), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(G290), .A2(G1986), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n807), .A2(new_n806), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1180), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1178), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1179), .B1(new_n740), .B2(new_n1183), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT46), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(new_n1192), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT47), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n799), .A2(new_n803), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1202));
  OAI22_X1  g777(.A1(new_n1201), .A2(new_n1202), .B1(G2067), .B2(new_n784), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1180), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1179), .A2(new_n1187), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT127), .Z(new_n1207));
  INV_X1    g782(.A(KEYINPUT48), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1185), .A2(new_n1180), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AND4_X1   g787(.A1(new_n1200), .A2(new_n1204), .A3(new_n1205), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1190), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g789(.A1(new_n679), .A2(G319), .A3(new_n661), .ZN(new_n1216));
  NOR2_X1   g790(.A1(G229), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g791(.A(new_n905), .B(new_n1217), .C1(new_n970), .C2(new_n971), .ZN(G225));
  INV_X1    g792(.A(G225), .ZN(G308));
endmodule


