//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n197), .A3(KEYINPUT70), .A4(new_n195), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(G110), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n195), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT24), .B(G110), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(G146), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  AOI211_X1 g027(.A(new_n213), .B(new_n210), .C1(KEYINPUT16), .C2(new_n207), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n202), .B(new_n206), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G125), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n209), .A2(G140), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT73), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT73), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n213), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n208), .A2(G146), .A3(new_n211), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT71), .B(G110), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n198), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n228), .A2(KEYINPUT72), .B1(new_n204), .B2(new_n205), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT72), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n198), .B2(new_n227), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n191), .B1(new_n216), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(KEYINPUT72), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n204), .A2(new_n205), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n225), .A3(new_n224), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n215), .A3(new_n190), .ZN(new_n238));
  INV_X1    g052(.A(G902), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n233), .A2(new_n238), .A3(KEYINPUT25), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G217), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(G234), .B2(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n233), .A2(new_n238), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n249), .A2(G902), .A3(new_n246), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n213), .A2(G143), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n213), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n253), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G137), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT11), .B1(new_n264), .B2(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(G134), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT65), .A2(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT65), .A2(G137), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT11), .A2(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G131), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n267), .B2(new_n271), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n263), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(G143), .B2(new_n213), .ZN(new_n277));
  OAI22_X1  g091(.A1(new_n277), .A2(new_n196), .B1(new_n256), .B2(new_n257), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n260), .A2(new_n261), .A3(new_n276), .A4(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n281));
  AOI21_X1  g095(.A(G134), .B1(new_n268), .B2(new_n269), .ZN(new_n282));
  INV_X1    g096(.A(new_n266), .ZN(new_n283));
  OAI21_X1  g097(.A(G131), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n275), .A2(KEYINPUT30), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n193), .A2(G116), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G113), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT2), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G113), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n294), .ZN(new_n296));
  XNOR2_X1  g110(.A(G116), .B(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n286), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT66), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n262), .A2(new_n259), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n253), .B1(new_n260), .B2(new_n261), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n258), .A2(KEYINPUT64), .A3(new_n259), .A4(new_n262), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n306), .B(new_n307), .C1(new_n273), .C2(new_n274), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n285), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT30), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI211_X1 g125(.A(KEYINPUT66), .B(KEYINPUT30), .C1(new_n308), .C2(new_n285), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n301), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n299), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n275), .A2(new_n314), .A3(new_n285), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT27), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n316), .A2(KEYINPUT68), .A3(new_n322), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n314), .B1(new_n308), .B2(new_n285), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n275), .A2(new_n314), .A3(new_n285), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT28), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n315), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n330), .B(KEYINPUT28), .C1(new_n327), .C2(new_n328), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n335), .B2(new_n321), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n325), .A2(new_n326), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n314), .B1(new_n275), .B2(new_n285), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT28), .B1(new_n328), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n315), .A2(new_n331), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT69), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G472), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n333), .A2(new_n322), .A3(new_n334), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT31), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n267), .A2(new_n271), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G131), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n352), .A2(new_n281), .B1(new_n263), .B2(new_n303), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n267), .A2(new_n271), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n354), .A2(new_n272), .B1(new_n278), .B2(new_n279), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n353), .A2(new_n307), .B1(new_n355), .B2(new_n284), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT66), .B1(new_n356), .B2(KEYINPUT30), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n309), .A2(new_n302), .A3(new_n310), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n300), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n328), .A2(new_n322), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n350), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n313), .A2(KEYINPUT31), .A3(new_n360), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n349), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G472), .A2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT32), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n333), .A2(new_n322), .A3(new_n334), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n313), .A2(KEYINPUT31), .A3(new_n360), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT31), .B1(new_n313), .B2(new_n360), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT32), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n365), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n252), .B1(new_n348), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n376));
  INV_X1    g190(.A(new_n279), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT1), .B1(new_n255), .B2(G146), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n378), .A2(G128), .B1(new_n260), .B2(new_n261), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G104), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n383), .B2(G107), .ZN(new_n386));
  AOI21_X1  g200(.A(G101), .B1(new_n383), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n381), .A3(G104), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n376), .B1(new_n380), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT10), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n383), .A2(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n386), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G101), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT74), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(KEYINPUT74), .A3(G101), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n390), .A2(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n402), .A3(G101), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n263), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n385), .A2(new_n390), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n280), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n376), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n393), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n273), .A2(new_n274), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n393), .A2(new_n405), .A3(new_n411), .A4(new_n409), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G140), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n188), .A2(G227), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n391), .A2(new_n279), .A3(new_n278), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n352), .A2(new_n281), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n422), .A2(new_n423), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n421), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n421), .B2(new_n424), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n418), .B1(new_n429), .B2(new_n414), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n239), .B1(new_n419), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(G469), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n421), .A2(new_n424), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n425), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n421), .A2(new_n424), .A3(new_n426), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n414), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n417), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT77), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n418), .B1(new_n413), .B2(new_n414), .ZN(new_n443));
  AND4_X1   g257(.A1(new_n414), .A2(new_n435), .A3(new_n436), .A4(new_n418), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n441), .B(new_n239), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n433), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT9), .B(G234), .ZN(new_n447));
  OAI21_X1  g261(.A(G221), .B1(new_n447), .B2(G902), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n299), .A2(new_n403), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n401), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n288), .A2(G119), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT5), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n291), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n298), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT78), .B1(new_n460), .B2(new_n391), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n457), .A2(new_n458), .B1(new_n297), .B2(new_n296), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT78), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n406), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n452), .B1(new_n454), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n401), .A2(new_n299), .A3(new_n403), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n467), .A2(new_n451), .A3(new_n461), .A4(new_n464), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT6), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT79), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT79), .A4(KEYINPUT6), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n466), .A2(KEYINPUT6), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n280), .B2(G125), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n278), .A2(KEYINPUT80), .A3(new_n209), .A4(new_n279), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n258), .A2(G125), .A3(new_n259), .A4(new_n262), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n188), .A2(G224), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n454), .A2(new_n465), .A3(new_n452), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n451), .B(KEYINPUT8), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n406), .A2(new_n462), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n459), .A2(new_n298), .B1(new_n390), .B2(new_n385), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT81), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n406), .A2(new_n462), .A3(KEYINPUT81), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n481), .A2(KEYINPUT7), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n476), .B2(new_n479), .ZN(new_n493));
  INV_X1    g307(.A(new_n479), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n494), .A2(KEYINPUT7), .A3(new_n481), .A4(new_n475), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n484), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n491), .A2(new_n493), .A3(new_n495), .A4(KEYINPUT82), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n483), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n483), .B2(new_n500), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n450), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n449), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n317), .A2(G143), .A3(G214), .ZN(new_n506));
  AOI21_X1  g320(.A(G143), .B1(new_n317), .B2(G214), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n317), .A2(G214), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n255), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n317), .A2(G143), .A3(G214), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n272), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n208), .A2(new_n211), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n213), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n511), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT17), .A3(G131), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n514), .A2(new_n516), .A3(new_n225), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n220), .A2(G146), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n224), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(KEYINPUT83), .A3(KEYINPUT18), .A4(G131), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n506), .A2(new_n507), .ZN(new_n523));
  NAND3_X1  g337(.A1(KEYINPUT83), .A2(KEYINPUT18), .A3(G131), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n383), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n519), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT19), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n222), .A2(new_n530), .A3(new_n223), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT84), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n220), .A2(new_n532), .A3(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT84), .B1(new_n207), .B2(new_n530), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n531), .A2(new_n213), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n210), .B1(new_n207), .B2(KEYINPUT16), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n508), .A2(new_n512), .B1(new_n536), .B2(G146), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n528), .B1(new_n538), .B2(new_n526), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT85), .B1(new_n529), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G475), .A2(G902), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n519), .A2(new_n526), .A3(new_n528), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n224), .A2(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n522), .A2(new_n544), .B1(new_n535), .B2(new_n537), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n542), .B(new_n543), .C1(new_n545), .C2(new_n528), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT20), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n529), .A2(new_n539), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n541), .B1(new_n550), .B2(KEYINPUT20), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n550), .B2(new_n541), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n528), .B1(new_n519), .B2(new_n526), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n239), .B1(new_n529), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n188), .A2(G952), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(G234), .B2(G237), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT21), .B(G898), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT88), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n239), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n255), .A2(G128), .ZN(new_n567));
  OAI21_X1  g381(.A(G134), .B1(new_n567), .B2(KEYINPUT13), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n255), .A2(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n196), .A2(G143), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT13), .A4(G134), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(KEYINPUT87), .A2(G122), .ZN(new_n575));
  NAND2_X1  g389(.A1(KEYINPUT87), .A2(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G116), .ZN(new_n578));
  INV_X1    g392(.A(G122), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G116), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n381), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n288), .B1(new_n575), .B2(new_n576), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n583), .A2(G107), .A3(new_n580), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n574), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n571), .B(G134), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(new_n381), .A3(new_n581), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT14), .B1(new_n579), .B2(G116), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT14), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n288), .A3(G122), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G107), .B1(new_n583), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n447), .A2(new_n245), .A3(G953), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n585), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n585), .B2(new_n593), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n239), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G478), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(KEYINPUT15), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n585), .A2(new_n593), .ZN(new_n601));
  INV_X1    g415(.A(new_n594), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n585), .A2(new_n593), .A3(new_n594), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n599), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n239), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n559), .A2(new_n566), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n375), .A2(new_n505), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  INV_X1    g425(.A(new_n566), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n450), .B(new_n612), .C1(new_n502), .C2(new_n503), .ZN(new_n613));
  NAND2_X1  g427(.A1(G478), .A2(G902), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n597), .B2(G478), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n605), .A2(KEYINPUT33), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n603), .B2(new_n604), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n615), .B1(new_n619), .B2(G478), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n559), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n449), .A2(new_n252), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n362), .A2(new_n363), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n624), .B2(new_n368), .ZN(new_n625));
  INV_X1    g439(.A(G472), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n364), .A2(new_n366), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n622), .A2(new_n623), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT89), .Z(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  INV_X1    g447(.A(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n547), .B(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT90), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n557), .A2(new_n638), .A3(G475), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n636), .A2(new_n608), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n613), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n623), .A3(new_n629), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  OAI22_X1  g459(.A1(new_n216), .A2(new_n232), .B1(KEYINPUT36), .B2(new_n191), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n246), .A2(G902), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n237), .A2(new_n215), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n244), .B2(new_n246), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n505), .A2(new_n609), .A3(new_n629), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n344), .A2(new_n345), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n239), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT68), .B1(new_n316), .B2(new_n322), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n324), .B(new_n321), .C1(new_n313), .C2(new_n315), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n657), .B1(new_n660), .B2(new_n336), .ZN(new_n661));
  AOI211_X1 g475(.A(KEYINPUT32), .B(new_n366), .C1(new_n624), .C2(new_n368), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n372), .B1(new_n371), .B2(new_n365), .ZN(new_n663));
  OAI22_X1  g477(.A1(new_n661), .A2(new_n626), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n561), .B1(new_n565), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n636), .A2(new_n640), .A3(new_n608), .A4(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n651), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n664), .A2(new_n505), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  INV_X1    g485(.A(new_n449), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n666), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n503), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n483), .A2(new_n500), .A3(new_n501), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n322), .B1(new_n313), .B2(new_n315), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n328), .A2(new_n338), .ZN(new_n683));
  AOI21_X1  g497(.A(G902), .B1(new_n683), .B2(new_n322), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n662), .B2(new_n663), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n608), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n555), .B2(new_n558), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n450), .A3(new_n651), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n681), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT92), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT92), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n676), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n255), .ZN(G45));
  AOI21_X1  g512(.A(new_n553), .B1(new_n547), .B2(KEYINPUT20), .ZN(new_n699));
  INV_X1    g513(.A(new_n558), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n620), .B(new_n667), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n651), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n664), .A2(new_n505), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  OAI21_X1  g518(.A(new_n239), .B1(new_n443), .B2(new_n444), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n448), .A3(new_n445), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT93), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n709), .A3(new_n448), .A4(new_n445), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n375), .A2(new_n622), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT94), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n712), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n642), .A2(new_n664), .A3(new_n251), .A4(new_n711), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NOR2_X1   g531(.A1(new_n504), .A2(new_n707), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n664), .A2(new_n718), .A3(new_n609), .A4(new_n652), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  INV_X1    g534(.A(KEYINPUT96), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n708), .A2(new_n612), .A3(new_n710), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n339), .A2(new_n340), .ZN(new_n723));
  OAI22_X1  g537(.A1(new_n369), .A2(new_n370), .B1(new_n321), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n365), .B(KEYINPUT95), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n251), .B(new_n726), .C1(new_n625), .C2(new_n626), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n690), .B(new_n450), .C1(new_n502), .C2(new_n503), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n721), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n722), .A2(new_n727), .A3(new_n729), .A4(KEYINPUT96), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n579), .ZN(G24));
  INV_X1    g548(.A(KEYINPUT97), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n559), .A2(new_n735), .A3(new_n620), .A4(new_n667), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n701), .A2(KEYINPUT97), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n726), .B(new_n652), .C1(new_n625), .C2(new_n626), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n718), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n677), .A2(new_n450), .A3(new_n678), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n448), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n437), .A2(KEYINPUT98), .A3(new_n417), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT98), .B1(new_n437), .B2(new_n417), .ZN(new_n748));
  OAI211_X1 g562(.A(G469), .B(new_n439), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n441), .A2(new_n239), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n445), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT99), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT99), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(new_n754), .A3(new_n445), .A4(new_n751), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n746), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n375), .A2(new_n745), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n743), .B1(new_n757), .B2(new_n738), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n664), .A2(new_n745), .A3(new_n251), .A4(new_n756), .ZN(new_n759));
  INV_X1    g573(.A(new_n738), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT100), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n758), .A2(new_n761), .A3(KEYINPUT100), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n272), .ZN(G33));
  INV_X1    g581(.A(new_n668), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n375), .A2(new_n768), .A3(new_n745), .A4(new_n756), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NOR2_X1   g584(.A1(new_n629), .A2(new_n651), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n699), .A2(new_n700), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT101), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(KEYINPUT43), .A3(new_n620), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n775));
  INV_X1    g589(.A(new_n620), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n559), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n774), .A2(KEYINPUT102), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT102), .B1(new_n774), .B2(new_n777), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT44), .B(new_n771), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(KEYINPUT103), .A3(new_n745), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n438), .B2(new_n439), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n441), .ZN(new_n783));
  OAI211_X1 g597(.A(KEYINPUT45), .B(new_n439), .C1(new_n747), .C2(new_n748), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n750), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT46), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n445), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n448), .B(new_n673), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n771), .B1(new_n778), .B2(new_n779), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n781), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT103), .B1(new_n780), .B2(new_n745), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  OAI21_X1  g609(.A(new_n448), .B1(new_n786), .B2(new_n787), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n664), .A2(new_n251), .A3(new_n701), .A4(new_n744), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n217), .ZN(G42));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n802));
  INV_X1    g616(.A(new_n798), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n706), .A2(new_n746), .A3(new_n445), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n561), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n806), .B(new_n727), .C1(new_n774), .C2(new_n777), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(new_n745), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n802), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n739), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n806), .B1(new_n774), .B2(new_n777), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n744), .A2(new_n707), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT112), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n251), .A2(new_n688), .A3(new_n561), .A4(new_n812), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n772), .A3(new_n776), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n450), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n681), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n707), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n807), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(KEYINPUT110), .A2(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n823), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n807), .A2(new_n820), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n818), .A2(KEYINPUT113), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n815), .A2(new_n828), .A3(new_n817), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT114), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n811), .A2(new_n812), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n812), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n739), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n817), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT113), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n824), .A2(new_n826), .ZN(new_n838));
  AND4_X1   g652(.A1(KEYINPUT114), .A2(new_n837), .A3(new_n829), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n809), .B1(new_n830), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT115), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n816), .A2(new_n559), .A3(new_n620), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n560), .B(KEYINPUT116), .Z(new_n843));
  AND2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n807), .A2(new_n821), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n833), .A2(new_n834), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT48), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n375), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n847), .B1(new_n846), .B2(new_n375), .ZN(new_n850));
  OAI221_X1 g664(.A(new_n844), .B1(new_n504), .B2(new_n845), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n803), .A2(KEYINPUT109), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n803), .A2(KEYINPUT109), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n804), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n808), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n818), .B1(new_n838), .B2(KEYINPUT111), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n855), .B(new_n856), .C1(KEYINPUT111), .C2(new_n838), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n851), .B1(new_n857), .B2(new_n802), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n859), .B(new_n809), .C1(new_n830), .C2(new_n839), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n841), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n610), .B(new_n719), .C1(new_n731), .C2(new_n732), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n600), .A2(new_n607), .A3(new_n667), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n637), .A3(new_n639), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n635), .A2(new_n651), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n865), .A2(new_n448), .A3(new_n446), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n740), .A2(new_n756), .B1(new_n664), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n769), .B1(new_n867), .B2(new_n744), .ZN(new_n868));
  INV_X1    g682(.A(new_n613), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n772), .A2(new_n620), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n772), .B2(new_n689), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n623), .A2(new_n869), .A3(new_n629), .A4(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n712), .A2(new_n716), .A3(new_n653), .A4(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n862), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n764), .A3(new_n875), .A4(new_n765), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n664), .B(new_n505), .C1(new_n669), .C2(new_n702), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n651), .A2(new_n667), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT105), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n730), .A2(new_n756), .A3(new_n880), .A4(new_n687), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n877), .A2(new_n741), .A3(new_n881), .A4(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT106), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n877), .A2(new_n741), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT106), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT52), .A4(new_n881), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n741), .A3(new_n881), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT107), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n883), .B(new_n886), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT108), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n887), .A2(new_n889), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT107), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n882), .B(new_n885), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT108), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n876), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n882), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n874), .A2(new_n764), .A3(new_n765), .A4(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n874), .A2(KEYINPUT53), .A3(new_n762), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n894), .B2(new_n900), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n903), .A2(new_n875), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT54), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n861), .A2(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n706), .A2(new_n445), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT49), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n776), .A2(new_n819), .A3(new_n746), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n773), .A2(new_n251), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT104), .Z(new_n917));
  OR2_X1    g731(.A1(new_n913), .A2(KEYINPUT49), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n681), .A3(new_n688), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n912), .A2(new_n919), .ZN(G75));
  INV_X1    g734(.A(new_n907), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n892), .A2(new_n893), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT108), .B1(new_n898), .B2(new_n899), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n903), .A2(new_n875), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n239), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(G210), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n482), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT55), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n188), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT56), .B1(new_n927), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n926), .A2(KEYINPUT117), .A3(G210), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n935), .B1(new_n939), .B2(new_n930), .ZN(G51));
  XNOR2_X1  g754(.A(new_n750), .B(KEYINPUT57), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n905), .B1(new_n924), .B2(new_n925), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n910), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n443), .B2(new_n444), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n926), .A2(new_n784), .A3(new_n783), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(G54));
  NAND2_X1  g760(.A1(new_n540), .A2(new_n546), .ZN(new_n947));
  INV_X1    g761(.A(new_n926), .ZN(new_n948));
  NAND2_X1  g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n934), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n948), .A2(new_n947), .A3(new_n949), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G60));
  INV_X1    g767(.A(new_n619), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n614), .B(KEYINPUT59), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n910), .B2(new_n942), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(KEYINPUT118), .A3(new_n934), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT118), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n924), .A2(new_n905), .A3(new_n925), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT54), .B1(new_n908), .B2(new_n909), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(new_n933), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n955), .B1(new_n906), .B2(new_n910), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n619), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n959), .A2(new_n964), .A3(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT119), .Z(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT60), .Z(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n908), .B2(new_n909), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n933), .B1(new_n971), .B2(new_n249), .ZN(new_n972));
  INV_X1    g786(.A(new_n970), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n924), .B2(new_n925), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n646), .A2(new_n649), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT120), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n975), .B(new_n970), .C1(new_n908), .C2(new_n909), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT120), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT61), .B(new_n972), .C1(new_n976), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(G66));
  INV_X1    g798(.A(G224), .ZN(new_n985));
  OAI21_X1  g799(.A(G953), .B1(new_n564), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n862), .A2(new_n873), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n928), .B1(G898), .B2(new_n188), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G69));
  OAI21_X1  g804(.A(new_n286), .B1(new_n311), .B2(new_n312), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(G900), .A2(G953), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n375), .A2(new_n730), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n884), .B(new_n769), .C1(new_n788), .C2(new_n996), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n766), .A2(new_n800), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n794), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(KEYINPUT124), .B(new_n995), .C1(new_n999), .C2(G953), .ZN(new_n1003));
  INV_X1    g817(.A(new_n800), .ZN(new_n1004));
  INV_X1    g818(.A(new_n674), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1005), .A2(new_n375), .A3(new_n745), .A4(new_n871), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1004), .B(new_n1006), .C1(new_n792), .C2(new_n793), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n694), .A2(new_n1008), .A3(new_n696), .A4(new_n884), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT121), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(KEYINPUT121), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n884), .ZN(new_n1013));
  OAI21_X1  g827(.A(KEYINPUT62), .B1(new_n697), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT122), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(KEYINPUT122), .B(KEYINPUT62), .C1(new_n697), .C2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(G953), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1002), .B(new_n1003), .C1(new_n1019), .C2(new_n993), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(KEYINPUT123), .Z(new_n1023));
  OAI211_X1 g837(.A(new_n1000), .B(new_n1023), .C1(new_n1019), .C2(new_n993), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1024), .ZN(G72));
  NAND3_X1  g839(.A1(new_n1012), .A2(new_n987), .A3(new_n1018), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT63), .Z(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT125), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(KEYINPUT126), .B1(new_n1030), .B2(new_n682), .ZN(new_n1031));
  INV_X1    g845(.A(new_n987), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1029), .B1(new_n999), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n1033), .A2(new_n315), .A3(new_n313), .A4(new_n322), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n901), .A2(new_n904), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n660), .B1(new_n359), .B2(new_n361), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1035), .A2(new_n1028), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1034), .A2(new_n1037), .A3(new_n934), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  INV_X1    g853(.A(new_n682), .ZN(new_n1040));
  AOI211_X1 g854(.A(new_n1039), .B(new_n1040), .C1(new_n1026), .C2(new_n1029), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1031), .A2(new_n1038), .A3(new_n1041), .ZN(G57));
endmodule


