

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U324 ( .A(n419), .B(KEYINPUT119), .ZN(n420) );
  XNOR2_X1 U325 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U326 ( .A(n396), .B(KEYINPUT48), .ZN(n537) );
  XNOR2_X1 U327 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U328 ( .A(n458), .B(n457), .ZN(n566) );
  XOR2_X1 U329 ( .A(KEYINPUT28), .B(n471), .Z(n543) );
  XOR2_X1 U330 ( .A(G29GAT), .B(KEYINPUT8), .Z(n291) );
  XNOR2_X1 U331 ( .A(n468), .B(KEYINPUT98), .ZN(n469) );
  XNOR2_X1 U332 ( .A(n470), .B(n469), .ZN(n475) );
  XNOR2_X1 U333 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n392) );
  XNOR2_X1 U334 ( .A(n349), .B(KEYINPUT71), .ZN(n350) );
  XNOR2_X1 U335 ( .A(n397), .B(n350), .ZN(n354) );
  XNOR2_X1 U336 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G8GAT), .Z(n398) );
  NOR2_X1 U338 ( .A1(n526), .A2(n422), .ZN(n423) );
  XNOR2_X1 U339 ( .A(n375), .B(n374), .ZN(n377) );
  XNOR2_X1 U340 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U341 ( .A(n537), .ZN(n539) );
  XNOR2_X1 U342 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U343 ( .A(n411), .B(n410), .ZN(n447) );
  XNOR2_X1 U344 ( .A(n329), .B(n328), .ZN(n563) );
  OR2_X1 U345 ( .A1(n582), .A2(n572), .ZN(n573) );
  INV_X1 U346 ( .A(G29GAT), .ZN(n487) );
  XNOR2_X1 U347 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n461) );
  XNOR2_X1 U348 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U349 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  XNOR2_X1 U350 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  INV_X1 U351 ( .A(KEYINPUT122), .ZN(n458) );
  XOR2_X1 U352 ( .A(G148GAT), .B(G85GAT), .Z(n293) );
  XNOR2_X1 U353 ( .A(G1GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U354 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U355 ( .A(G57GAT), .B(G155GAT), .Z(n295) );
  XNOR2_X1 U356 ( .A(G127GAT), .B(KEYINPUT6), .ZN(n294) );
  XNOR2_X1 U357 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U358 ( .A(n297), .B(n296), .Z(n305) );
  XOR2_X1 U359 ( .A(KEYINPUT88), .B(KEYINPUT2), .Z(n299) );
  XNOR2_X1 U360 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n298) );
  XNOR2_X1 U361 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U362 ( .A(G141GAT), .B(n300), .Z(n429) );
  XOR2_X1 U363 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n302) );
  XNOR2_X1 U364 ( .A(KEYINPUT1), .B(KEYINPUT92), .ZN(n301) );
  XNOR2_X1 U365 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U366 ( .A(n429), .B(n303), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n312) );
  XOR2_X1 U368 ( .A(G120GAT), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n446) );
  XOR2_X1 U371 ( .A(G162GAT), .B(n446), .Z(n309) );
  NAND2_X1 U372 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U373 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U374 ( .A(G29GAT), .B(n310), .Z(n311) );
  XOR2_X1 U375 ( .A(n312), .B(n311), .Z(n477) );
  INV_X1 U376 ( .A(n477), .ZN(n526) );
  XNOR2_X1 U377 ( .A(KEYINPUT7), .B(KEYINPUT67), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n291), .B(n313), .ZN(n378) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(G162GAT), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n314), .B(KEYINPUT72), .ZN(n428) );
  XNOR2_X1 U381 ( .A(n378), .B(n428), .ZN(n319) );
  XOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT74), .Z(n316) );
  NAND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U384 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U385 ( .A(n317), .B(KEYINPUT73), .Z(n318) );
  XNOR2_X1 U386 ( .A(n319), .B(n318), .ZN(n323) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .ZN(n361) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(n361), .ZN(n321) );
  XOR2_X1 U389 ( .A(G43GAT), .B(G134GAT), .Z(n444) );
  XNOR2_X1 U390 ( .A(n444), .B(G92GAT), .ZN(n320) );
  XNOR2_X1 U391 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U392 ( .A(n323), .B(n322), .Z(n329) );
  XOR2_X1 U393 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n325) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(KEYINPUT11), .ZN(n324) );
  XNOR2_X1 U395 ( .A(n325), .B(n324), .ZN(n327) );
  XNOR2_X1 U396 ( .A(G190GAT), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U397 ( .A(KEYINPUT36), .B(n563), .ZN(n583) );
  XOR2_X1 U398 ( .A(KEYINPUT77), .B(G78GAT), .Z(n331) );
  XNOR2_X1 U399 ( .A(G183GAT), .B(G64GAT), .ZN(n330) );
  XNOR2_X1 U400 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U401 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n333) );
  XNOR2_X1 U402 ( .A(KEYINPUT76), .B(KEYINPUT12), .ZN(n332) );
  XNOR2_X1 U403 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n335), .B(n334), .ZN(n346) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G57GAT), .ZN(n336) );
  XNOR2_X1 U406 ( .A(n336), .B(KEYINPUT13), .ZN(n358) );
  XOR2_X1 U407 ( .A(n358), .B(KEYINPUT14), .Z(n338) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U409 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U410 ( .A(G22GAT), .B(G155GAT), .Z(n435) );
  XOR2_X1 U411 ( .A(n435), .B(G211GAT), .Z(n340) );
  XOR2_X1 U412 ( .A(G15GAT), .B(G127GAT), .Z(n449) );
  XNOR2_X1 U413 ( .A(G8GAT), .B(n449), .ZN(n339) );
  XNOR2_X1 U414 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U415 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n367) );
  INV_X1 U417 ( .A(n367), .ZN(n343) );
  XOR2_X1 U418 ( .A(n344), .B(n343), .Z(n345) );
  XNOR2_X1 U419 ( .A(n346), .B(n345), .ZN(n579) );
  NOR2_X1 U420 ( .A1(n583), .A2(n579), .ZN(n347) );
  XNOR2_X1 U421 ( .A(n347), .B(KEYINPUT45), .ZN(n365) );
  XNOR2_X1 U422 ( .A(G92GAT), .B(G64GAT), .ZN(n348) );
  XNOR2_X1 U423 ( .A(n348), .B(G204GAT), .ZN(n397) );
  AND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XOR2_X1 U425 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n352) );
  XNOR2_X1 U426 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n351) );
  XNOR2_X1 U427 ( .A(n352), .B(n351), .ZN(n353) );
  NAND2_X1 U428 ( .A1(n354), .A2(n353), .ZN(n356) );
  OR2_X1 U429 ( .A1(n354), .A2(n353), .ZN(n355) );
  NAND2_X1 U430 ( .A1(n356), .A2(n355), .ZN(n360) );
  XNOR2_X1 U431 ( .A(G148GAT), .B(G106GAT), .ZN(n357) );
  XNOR2_X1 U432 ( .A(n357), .B(G78GAT), .ZN(n426) );
  XOR2_X1 U433 ( .A(n358), .B(n426), .Z(n359) );
  XNOR2_X1 U434 ( .A(n360), .B(n359), .ZN(n364) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(G120GAT), .ZN(n362) );
  XOR2_X1 U436 ( .A(n362), .B(n361), .Z(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n576) );
  NAND2_X1 U438 ( .A1(n365), .A2(n576), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n366), .B(KEYINPUT115), .ZN(n385) );
  XOR2_X1 U440 ( .A(G43GAT), .B(G50GAT), .Z(n369) );
  XOR2_X1 U441 ( .A(n398), .B(n367), .Z(n368) );
  XNOR2_X1 U442 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U443 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n371) );
  XNOR2_X1 U444 ( .A(G22GAT), .B(G15GAT), .ZN(n370) );
  XOR2_X1 U445 ( .A(n371), .B(n370), .Z(n373) );
  NAND2_X1 U446 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  INV_X1 U447 ( .A(KEYINPUT66), .ZN(n376) );
  XNOR2_X1 U448 ( .A(n377), .B(n376), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n378), .B(KEYINPUT69), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U451 ( .A(G197GAT), .B(G141GAT), .Z(n382) );
  XNOR2_X1 U452 ( .A(G169GAT), .B(G113GAT), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n572) );
  NAND2_X1 U455 ( .A1(n385), .A2(n572), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n386), .B(KEYINPUT116), .ZN(n395) );
  XOR2_X1 U457 ( .A(n576), .B(KEYINPUT41), .Z(n557) );
  NOR2_X1 U458 ( .A1(n572), .A2(n557), .ZN(n388) );
  XNOR2_X1 U459 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n387) );
  XNOR2_X1 U460 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U461 ( .A(KEYINPUT111), .B(n579), .ZN(n548) );
  NOR2_X1 U462 ( .A1(n389), .A2(n548), .ZN(n390) );
  XNOR2_X1 U463 ( .A(n390), .B(KEYINPUT113), .ZN(n391) );
  INV_X1 U464 ( .A(n563), .ZN(n551) );
  NOR2_X1 U465 ( .A1(n391), .A2(n551), .ZN(n393) );
  XNOR2_X1 U466 ( .A(n393), .B(n392), .ZN(n394) );
  NAND2_X1 U467 ( .A1(n395), .A2(n394), .ZN(n396) );
  XOR2_X1 U468 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U471 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n402) );
  XNOR2_X1 U472 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U474 ( .A(n404), .B(n403), .Z(n418) );
  XOR2_X1 U475 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n406) );
  XNOR2_X1 U476 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n407), .B(KEYINPUT19), .ZN(n411) );
  XOR2_X1 U479 ( .A(G190GAT), .B(G183GAT), .Z(n409) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G176GAT), .ZN(n408) );
  XOR2_X1 U481 ( .A(KEYINPUT84), .B(KEYINPUT21), .Z(n413) );
  XNOR2_X1 U482 ( .A(G218GAT), .B(KEYINPUT86), .ZN(n412) );
  XNOR2_X1 U483 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U484 ( .A(n414), .B(KEYINPUT85), .Z(n416) );
  XNOR2_X1 U485 ( .A(G197GAT), .B(G211GAT), .ZN(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n439) );
  XNOR2_X1 U487 ( .A(n447), .B(n439), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n528) );
  NAND2_X1 U489 ( .A1(n537), .A2(n528), .ZN(n421) );
  XOR2_X1 U490 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n419) );
  XNOR2_X1 U491 ( .A(n423), .B(KEYINPUT64), .ZN(n570) );
  XOR2_X1 U492 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n425) );
  XNOR2_X1 U493 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n424) );
  XNOR2_X1 U494 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U495 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n441) );
  XOR2_X1 U498 ( .A(KEYINPUT89), .B(KEYINPUT83), .Z(n433) );
  XNOR2_X1 U499 ( .A(G204GAT), .B(KEYINPUT91), .ZN(n432) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U501 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U502 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U504 ( .A(n439), .B(n438), .Z(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n471) );
  NAND2_X1 U506 ( .A1(n570), .A2(n471), .ZN(n443) );
  XOR2_X1 U507 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n442) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n456) );
  NAND2_X1 U509 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n445), .B(n444), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n447), .B(n446), .ZN(n451) );
  XNOR2_X1 U512 ( .A(KEYINPUT20), .B(KEYINPUT79), .ZN(n448) );
  XNOR2_X1 U513 ( .A(G99GAT), .B(G71GAT), .ZN(n452) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X2 U515 ( .A(n455), .B(n454), .ZN(n540) );
  NAND2_X1 U516 ( .A1(n456), .A2(n540), .ZN(n457) );
  NAND2_X1 U517 ( .A1(n566), .A2(n548), .ZN(n460) );
  XNOR2_X1 U518 ( .A(KEYINPUT124), .B(G183GAT), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n460), .B(n459), .ZN(G1350GAT) );
  NAND2_X1 U520 ( .A1(n566), .A2(n551), .ZN(n462) );
  INV_X1 U521 ( .A(n543), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n528), .B(KEYINPUT27), .ZN(n473) );
  NAND2_X1 U523 ( .A1(n526), .A2(n473), .ZN(n538) );
  XNOR2_X1 U524 ( .A(KEYINPUT82), .B(n540), .ZN(n463) );
  NOR2_X1 U525 ( .A1(n538), .A2(n463), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n481) );
  INV_X1 U527 ( .A(KEYINPUT99), .ZN(n479) );
  NAND2_X1 U528 ( .A1(n528), .A2(n540), .ZN(n466) );
  XOR2_X1 U529 ( .A(KEYINPUT97), .B(n466), .Z(n467) );
  NAND2_X1 U530 ( .A1(n471), .A2(n467), .ZN(n470) );
  INV_X1 U531 ( .A(KEYINPUT25), .ZN(n468) );
  NOR2_X1 U532 ( .A1(n471), .A2(n540), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT26), .ZN(n569) );
  NAND2_X1 U534 ( .A1(n473), .A2(n569), .ZN(n474) );
  NAND2_X1 U535 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(KEYINPUT100), .ZN(n496) );
  NAND2_X1 U540 ( .A1(n496), .A2(n579), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n583), .A2(n483), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n484), .ZN(n525) );
  INV_X1 U543 ( .A(n572), .ZN(n567) );
  NAND2_X1 U544 ( .A1(n567), .A2(n576), .ZN(n498) );
  NOR2_X1 U545 ( .A1(n525), .A2(n498), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n512) );
  NAND2_X1 U548 ( .A1(n512), .A2(n526), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n488) );
  INV_X1 U550 ( .A(n557), .ZN(n545) );
  NAND2_X1 U551 ( .A1(n545), .A2(n566), .ZN(n494) );
  XOR2_X1 U552 ( .A(G176GAT), .B(KEYINPUT57), .Z(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1349GAT) );
  NOR2_X1 U556 ( .A1(n551), .A2(n579), .ZN(n495) );
  XNOR2_X1 U557 ( .A(KEYINPUT16), .B(n495), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n497), .A2(n496), .ZN(n516) );
  NOR2_X1 U559 ( .A1(n498), .A2(n516), .ZN(n499) );
  XOR2_X1 U560 ( .A(KEYINPUT101), .B(n499), .Z(n506) );
  NAND2_X1 U561 ( .A1(n526), .A2(n506), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U564 ( .A1(n506), .A2(n528), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT102), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G8GAT), .B(n503), .ZN(G1325GAT) );
  XOR2_X1 U567 ( .A(G15GAT), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U568 ( .A1(n506), .A2(n540), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NAND2_X1 U570 ( .A1(n543), .A2(n506), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n507), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U572 ( .A1(n512), .A2(n528), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n510) );
  NAND2_X1 U575 ( .A1(n512), .A2(n540), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G43GAT), .B(n511), .ZN(G1330GAT) );
  XNOR2_X1 U578 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n543), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1331GAT) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  NOR2_X1 U582 ( .A1(n557), .A2(n567), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(KEYINPUT107), .ZN(n524) );
  NOR2_X1 U584 ( .A1(n516), .A2(n524), .ZN(n521) );
  NAND2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n528), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n540), .A2(n521), .ZN(n520) );
  XNOR2_X1 U590 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U592 ( .A1(n521), .A2(n543), .ZN(n522) );
  XNOR2_X1 U593 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NOR2_X1 U594 ( .A1(n525), .A2(n524), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n533), .A2(n526), .ZN(n527) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n528), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n529), .B(KEYINPUT108), .ZN(n530) );
  XNOR2_X1 U599 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  XOR2_X1 U600 ( .A(G99GAT), .B(KEYINPUT109), .Z(n532) );
  NAND2_X1 U601 ( .A1(n533), .A2(n540), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U604 ( .A1(n533), .A2(n543), .ZN(n534) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U606 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  NOR2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n555), .A2(n540), .ZN(n541) );
  XOR2_X1 U609 ( .A(KEYINPUT117), .B(n541), .Z(n542) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n552), .A2(n567), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U614 ( .A1(n552), .A2(n545), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  NAND2_X1 U616 ( .A1(n552), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(KEYINPUT50), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1343GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n569), .ZN(n562) );
  NOR2_X1 U623 ( .A1(n572), .A2(n562), .ZN(n556) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n556), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n557), .A2(n562), .ZN(n559) );
  XNOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n579), .A2(n562), .ZN(n561) );
  XOR2_X1 U630 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT118), .B(n564), .Z(n565) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(n565), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(n571), .Z(n582) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  OR2_X1 U642 ( .A1(n582), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT126), .ZN(n581) );
  OR2_X1 U645 ( .A1(n579), .A2(n582), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

