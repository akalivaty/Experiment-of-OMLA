//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT94), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT68), .A2(G953), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT68), .A2(G953), .ZN(new_n192));
  OAI211_X1 g006(.A(G214), .B(new_n190), .C1(new_n191), .C2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT86), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT68), .B(G953), .ZN(new_n196));
  INV_X1    g010(.A(new_n194), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n196), .A2(G214), .A3(new_n190), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT87), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT18), .A3(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT87), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G125), .B(G140), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n205), .B(KEYINPUT88), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(new_n206), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n202), .A2(KEYINPUT87), .A3(KEYINPUT18), .A4(G131), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n195), .A2(new_n198), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G125), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n216), .A2(KEYINPUT16), .A3(G140), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n205), .B2(KEYINPUT16), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT19), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n208), .B2(new_n220), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n215), .B(new_n219), .C1(G146), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT89), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(G113), .B(G122), .Z(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT90), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n211), .A2(new_n223), .A3(KEYINPUT89), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n218), .B(new_n206), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(new_n212), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n233), .B(KEYINPUT91), .C1(new_n234), .C2(new_n212), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n212), .A2(new_n234), .A3(new_n214), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT92), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT92), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n212), .A2(new_n241), .A3(new_n234), .A4(new_n214), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n237), .A2(new_n238), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n230), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(new_n211), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n232), .A2(KEYINPUT93), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT93), .B1(new_n232), .B2(new_n245), .ZN(new_n247));
  OAI211_X1 g061(.A(KEYINPUT20), .B(new_n189), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n232), .A2(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n189), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G902), .ZN(new_n253));
  INV_X1    g067(.A(new_n245), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n244), .B1(new_n243), .B2(new_n211), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G475), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n248), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G122), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G107), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G128), .B(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G128), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n267), .B(G134), .C1(KEYINPUT13), .C2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n265), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n264), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n266), .B(new_n271), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT95), .B1(new_n262), .B2(KEYINPUT14), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n262), .A2(KEYINPUT14), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT14), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n261), .A4(G122), .ZN(new_n280));
  AND4_X1   g094(.A1(new_n260), .A2(new_n276), .A3(new_n277), .A4(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n274), .B(new_n275), .C1(new_n281), .C2(new_n264), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT9), .B(G234), .Z(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(G217), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n273), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n253), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n294));
  INV_X1    g108(.A(G478), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(KEYINPUT97), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n292), .B(KEYINPUT97), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI211_X1 g115(.A(new_n253), .B(new_n196), .C1(G234), .C2(G237), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT21), .B(G898), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G952), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(KEYINPUT98), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT98), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n285), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G234), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n190), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n312), .B(KEYINPUT99), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n258), .A2(new_n301), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(G469), .A2(G902), .ZN(new_n316));
  INV_X1    g130(.A(G469), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n206), .A2(G143), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n268), .A2(G146), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .A4(G128), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G128), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT1), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(new_n318), .A3(new_n319), .A4(KEYINPUT78), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n318), .A2(new_n319), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n318), .B2(KEYINPUT1), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n323), .B(new_n326), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n229), .A2(G107), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n229), .A2(G107), .ZN(new_n332));
  OAI21_X1  g146(.A(G101), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n264), .A3(G104), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .A4(new_n330), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n329), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n338), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n268), .A2(G146), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT64), .B1(new_n206), .B2(G143), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT64), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n268), .A3(G146), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n341), .B(new_n321), .C1(new_n346), .C2(new_n328), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(KEYINPUT79), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT11), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n271), .B2(G137), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n271), .A2(G137), .ZN(new_n351));
  INV_X1    g165(.A(G137), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT11), .A3(G134), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G131), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n350), .A2(new_n353), .A3(new_n213), .A4(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n321), .B1(new_n346), .B2(new_n328), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n339), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n348), .A2(new_n362), .A3(KEYINPUT12), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT12), .B1(new_n348), .B2(new_n362), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n334), .A2(new_n336), .A3(new_n330), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G101), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT77), .B1(new_n367), .B2(KEYINPUT4), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .A4(G101), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n344), .B1(new_n268), .B2(G146), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n206), .A2(KEYINPUT64), .A3(G143), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n318), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT0), .A2(G128), .ZN(new_n376));
  OR2_X1    g190(.A1(KEYINPUT0), .A2(G128), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n318), .A2(new_n319), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n379), .A2(new_n376), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n367), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n367), .A2(new_n384), .A3(KEYINPUT4), .A4(new_n338), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n372), .A2(new_n381), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n340), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n339), .A2(new_n359), .A3(KEYINPUT10), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n386), .A2(new_n358), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n196), .A2(G227), .ZN(new_n391));
  XNOR2_X1  g205(.A(G110), .B(G140), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n365), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n357), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n397), .B2(new_n390), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n317), .B(new_n253), .C1(new_n395), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(KEYINPUT80), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n401), .A3(new_n393), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n390), .B1(new_n363), .B2(new_n364), .ZN(new_n404));
  INV_X1    g218(.A(new_n393), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n316), .B(new_n399), .C1(new_n407), .C2(new_n317), .ZN(new_n408));
  INV_X1    g222(.A(G221), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n284), .B2(new_n253), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n315), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n219), .A2(new_n207), .ZN(new_n415));
  INV_X1    g229(.A(G119), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G128), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT73), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(new_n416), .B2(G128), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT74), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI22_X1  g237(.A1(new_n324), .A2(G119), .B1(KEYINPUT73), .B2(KEYINPUT23), .ZN(new_n424));
  INV_X1    g238(.A(new_n422), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n418), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(KEYINPUT23), .B2(new_n418), .ZN(new_n429));
  INV_X1    g243(.A(G110), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT24), .B(G110), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(G119), .B(G128), .Z(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n415), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n233), .ZN(new_n438));
  OAI221_X1 g252(.A(new_n438), .B1(new_n434), .B2(new_n433), .C1(new_n429), .C2(new_n430), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n196), .A2(G221), .A3(G234), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT22), .Z(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(new_n352), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(G137), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n429), .A2(new_n430), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n433), .A2(new_n434), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n445), .A2(new_n233), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n447), .B2(new_n436), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT25), .B1(new_n449), .B2(G902), .ZN(new_n450));
  INV_X1    g264(.A(new_n286), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(G234), .B2(new_n253), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT25), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n443), .A2(new_n448), .A3(new_n453), .A4(new_n253), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n449), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n452), .A2(G902), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n457), .B(KEYINPUT75), .Z(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n357), .A2(new_n378), .A3(new_n380), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT67), .ZN(new_n463));
  XOR2_X1   g277(.A(G116), .B(G119), .Z(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT2), .B(G113), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n465), .ZN(new_n467));
  XNOR2_X1  g281(.A(G116), .B(G119), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT67), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n470), .B2(new_n465), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(KEYINPUT66), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n466), .A2(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT65), .B1(new_n271), .B2(G137), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n352), .A3(G134), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n476), .A3(new_n351), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G131), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n359), .A2(new_n356), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n462), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT28), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n462), .A2(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n469), .A2(new_n466), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n471), .A2(new_n472), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n462), .A2(new_n473), .A3(new_n479), .A4(KEYINPUT28), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G101), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n196), .A2(G210), .A3(new_n190), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n490), .B(new_n337), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n492), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n480), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n483), .A2(KEYINPUT30), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n462), .A2(new_n504), .A3(new_n479), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n502), .B1(new_n506), .B2(new_n486), .ZN(new_n507));
  INV_X1    g321(.A(new_n497), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT31), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n462), .A2(new_n504), .A3(new_n479), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n504), .B1(new_n462), .B2(new_n479), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n486), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(KEYINPUT31), .A3(new_n508), .A4(new_n480), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n501), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(G472), .A2(G902), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(KEYINPUT32), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT32), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n508), .A3(new_n480), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n500), .B1(new_n521), .B2(new_n513), .ZN(new_n522));
  INV_X1    g336(.A(new_n516), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n517), .A2(new_n524), .A3(KEYINPUT70), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n515), .A2(new_n516), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n518), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n507), .A2(new_n508), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n489), .A2(new_n499), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n487), .A2(KEYINPUT71), .A3(new_n480), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n483), .A2(new_n535), .A3(new_n486), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(KEYINPUT28), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT29), .A3(new_n482), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n497), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G472), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n461), .B1(new_n529), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n383), .A2(new_n385), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n542), .A2(KEYINPUT81), .A3(new_n486), .A4(new_n372), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT5), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n416), .A3(G116), .ZN(new_n545));
  OAI211_X1 g359(.A(G113), .B(new_n545), .C1(new_n464), .C2(new_n544), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n484), .A2(new_n339), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n372), .A2(new_n486), .A3(new_n383), .A4(new_n385), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT81), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  XOR2_X1   g365(.A(G110), .B(G122), .Z(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n552), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n543), .A2(new_n550), .A3(new_n554), .A4(new_n547), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n553), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n553), .A2(KEYINPUT6), .A3(new_n555), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT6), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n558), .A3(new_n552), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT82), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n556), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n359), .A2(G125), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n381), .B2(new_n216), .ZN(new_n564));
  INV_X1    g378(.A(G224), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(G953), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n564), .B(new_n566), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G210), .B1(G237), .B2(G902), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT84), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n552), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n484), .A2(new_n546), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n341), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n575), .B2(new_n547), .ZN(new_n576));
  INV_X1    g390(.A(new_n564), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT7), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT83), .B1(new_n566), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n381), .A2(new_n216), .ZN(new_n581));
  OAI221_X1 g395(.A(new_n564), .B1(new_n578), .B2(new_n566), .C1(new_n581), .C2(KEYINPUT83), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n555), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n253), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n569), .A2(new_n572), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n553), .A2(KEYINPUT6), .A3(new_n555), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n560), .A3(new_n559), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n567), .B1(new_n588), .B2(new_n556), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n571), .B1(new_n589), .B2(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G214), .B1(G237), .B2(G902), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT85), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT85), .ZN(new_n594));
  INV_X1    g408(.A(new_n592), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n594), .B(new_n595), .C1(new_n586), .C2(new_n590), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n414), .B(new_n541), .C1(new_n593), .C2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n455), .A2(new_n460), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n411), .A3(new_n408), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n522), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n526), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n599), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n603), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n413), .A2(KEYINPUT100), .A3(new_n600), .A4(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n569), .A2(new_n570), .A3(new_n585), .ZN(new_n608));
  INV_X1    g422(.A(new_n570), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n589), .B2(new_n584), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n595), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n313), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT101), .B(KEYINPUT33), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n291), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n290), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n290), .A2(new_n617), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(KEYINPUT33), .A3(new_n288), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n291), .A2(KEYINPUT102), .A3(new_n613), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n616), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n622), .A2(new_n623), .A3(G478), .A4(new_n253), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n292), .A2(new_n295), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n616), .A2(new_n620), .A3(G478), .A4(new_n621), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT104), .B1(new_n626), .B2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n258), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n607), .A2(new_n612), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n248), .A2(new_n257), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT93), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n249), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n232), .A2(new_n245), .A3(KEYINPUT93), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT20), .B1(new_n638), .B2(new_n189), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n634), .A2(new_n639), .A3(new_n300), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n607), .A2(new_n612), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND2_X1  g457(.A1(new_n437), .A2(new_n439), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n459), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n455), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n414), .B(new_n650), .C1(new_n593), .C2(new_n596), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(new_n603), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT37), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n430), .ZN(G12));
  XNOR2_X1  g468(.A(new_n311), .B(KEYINPUT105), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n302), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n634), .A2(new_n639), .A3(new_n300), .A4(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n412), .B1(new_n529), .B2(new_n540), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n611), .A4(new_n650), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n657), .B(KEYINPUT39), .Z(new_n662));
  AND2_X1   g476(.A1(new_n413), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  INV_X1    g478(.A(G472), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n534), .A2(new_n499), .A3(new_n536), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n519), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n665), .B1(new_n669), .B2(new_n253), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n525), .B2(new_n528), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n650), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n591), .B(KEYINPUT38), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n258), .A2(new_n592), .A3(new_n301), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n664), .A2(new_n672), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  INV_X1    g490(.A(new_n657), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n258), .A2(new_n628), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n659), .A2(new_n611), .A3(new_n650), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  NAND2_X1  g494(.A1(new_n529), .A2(new_n540), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n395), .A2(new_n398), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G469), .B1(new_n683), .B2(G902), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n684), .A2(new_n411), .A3(new_n399), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n681), .A2(new_n600), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n612), .A2(new_n630), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n313), .A3(new_n611), .A4(new_n640), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  NAND2_X1  g505(.A1(new_n608), .A2(new_n610), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n692), .A2(new_n592), .A3(new_n650), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n681), .A3(new_n315), .A4(new_n685), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT107), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  AND2_X1   g510(.A1(new_n674), .A2(new_n692), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n537), .A2(new_n482), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n521), .A2(new_n513), .B1(new_n698), .B2(new_n499), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(new_n523), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n515), .A2(new_n253), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT108), .B1(new_n701), .B2(G472), .ZN(new_n702));
  OAI211_X1 g516(.A(KEYINPUT108), .B(G472), .C1(new_n522), .C2(G902), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n700), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n461), .A3(new_n314), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n697), .A2(new_n685), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  NAND3_X1  g522(.A1(new_n258), .A2(new_n628), .A3(new_n677), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n705), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n611), .A3(new_n650), .A4(new_n685), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  AND3_X1   g526(.A1(new_n586), .A2(new_n590), .A3(new_n592), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n412), .A2(KEYINPUT109), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n408), .A2(new_n715), .A3(new_n411), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n713), .A2(new_n541), .A3(new_n678), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n408), .A2(new_n715), .A3(new_n411), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n715), .B1(new_n408), .B2(new_n411), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n586), .A2(new_n590), .A3(new_n592), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n540), .A2(new_n524), .A3(new_n517), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(new_n600), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n678), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n720), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND4_X1  g544(.A1(new_n658), .A2(new_n713), .A3(new_n541), .A4(new_n717), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n725), .A2(new_n733), .A3(new_n541), .A4(new_n658), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  XNOR2_X1  g550(.A(new_n407), .B(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n316), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n740), .B(G469), .C1(new_n737), .C2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n399), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n411), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n662), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(KEYINPUT111), .Z(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n713), .ZN(new_n747));
  INV_X1    g561(.A(new_n258), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n628), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(KEYINPUT43), .A3(new_n628), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n603), .A3(new_n650), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT44), .Z(new_n755));
  OR2_X1    g569(.A1(new_n747), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  NOR2_X1   g571(.A1(new_n709), .A2(new_n600), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n724), .A2(new_n681), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n758), .B(new_n759), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  NAND2_X1  g578(.A1(new_n713), .A2(new_n685), .ZN(new_n765));
  INV_X1    g579(.A(new_n671), .ZN(new_n766));
  OR4_X1    g580(.A1(new_n461), .A2(new_n765), .A3(new_n311), .A4(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n258), .A3(new_n628), .ZN(new_n768));
  INV_X1    g582(.A(new_n765), .ZN(new_n769));
  INV_X1    g583(.A(new_n650), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n705), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n753), .A2(new_n655), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT118), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(KEYINPUT118), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n769), .B(new_n771), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n773), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(KEYINPUT120), .A3(new_n769), .A4(new_n771), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n768), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n705), .A2(new_n461), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n685), .B(new_n784), .C1(new_n774), .C2(new_n775), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n673), .A2(new_n592), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n784), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n779), .B2(new_n773), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(KEYINPUT50), .A3(new_n685), .A4(new_n786), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n713), .ZN(new_n793));
  INV_X1    g607(.A(new_n762), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(KEYINPUT119), .A3(new_n760), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n684), .A2(new_n399), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT112), .Z(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n411), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT119), .B1(new_n794), .B2(new_n760), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n782), .B(new_n792), .C1(new_n793), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n308), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n761), .A2(new_n762), .A3(new_n798), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n793), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n804), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n782), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g624(.A(KEYINPUT121), .B(new_n768), .C1(new_n778), .C2(new_n781), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n792), .B(new_n808), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n780), .A2(new_n727), .A3(new_n769), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT48), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n805), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n711), .A2(new_n660), .A3(new_n679), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n671), .A2(new_n650), .A3(new_n657), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n413), .A3(new_n692), .A4(new_n674), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT52), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n711), .A3(new_n660), .A4(new_n679), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT113), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n597), .B(new_n694), .C1(new_n651), .C2(new_n603), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n591), .A2(new_n592), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n594), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n591), .A2(KEYINPUT85), .A3(new_n592), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n629), .B1(new_n300), .B2(new_n258), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n604), .A2(new_n832), .A3(new_n606), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n831), .A2(new_n833), .A3(new_n313), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n687), .A2(new_n690), .A3(new_n707), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n827), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n634), .A2(new_n639), .A3(new_n301), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n659), .A2(new_n837), .A3(new_n650), .A4(new_n677), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n771), .A2(new_n678), .A3(new_n717), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n713), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n735), .A2(new_n729), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n826), .A2(new_n836), .A3(KEYINPUT53), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT116), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n842), .A2(new_n827), .A3(new_n834), .A4(new_n835), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT53), .A4(new_n826), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n822), .A2(new_n823), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n822), .A2(new_n823), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT114), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n817), .A2(KEYINPUT52), .A3(new_n820), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n825), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n852), .A2(new_n836), .A3(new_n843), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n856), .A2(KEYINPUT115), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT115), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n816), .B(new_n849), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n846), .A2(new_n826), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n857), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n857), .B2(new_n856), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT117), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n860), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n790), .A2(new_n611), .A3(new_n685), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n815), .A2(new_n866), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n767), .A2(new_n629), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n870), .A2(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n592), .B1(new_n797), .B2(KEYINPUT49), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n749), .ZN(new_n874));
  INV_X1    g688(.A(new_n673), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n410), .B(new_n766), .C1(new_n797), .C2(KEYINPUT49), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n874), .A2(new_n600), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n877), .ZN(G75));
  NAND2_X1  g692(.A1(new_n856), .A2(new_n857), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n856), .A2(KEYINPUT115), .A3(new_n857), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n253), .B1(new_n883), .B2(new_n849), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(G210), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n562), .B(new_n567), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n885), .B2(new_n886), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n196), .A2(G952), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G51));
  AOI211_X1 g706(.A(new_n253), .B(new_n738), .C1(new_n883), .C2(new_n849), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n316), .B(KEYINPUT57), .Z(new_n894));
  AOI21_X1  g708(.A(new_n816), .B1(new_n883), .B2(new_n849), .ZN(new_n895));
  INV_X1    g709(.A(new_n860), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n897), .B2(new_n682), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n898), .B2(new_n891), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n900));
  INV_X1    g714(.A(new_n891), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n849), .B1(new_n858), .B2(new_n859), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n860), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n683), .B1(new_n904), .B2(new_n894), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n900), .B(new_n901), .C1(new_n905), .C2(new_n893), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n899), .A2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n638), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(new_n901), .ZN(G60));
  XNOR2_X1  g724(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n295), .A2(new_n253), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n911), .B(new_n912), .Z(new_n913));
  NAND3_X1  g727(.A1(new_n904), .A2(new_n622), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n913), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n866), .B2(new_n868), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n901), .B(new_n914), .C1(new_n916), .C2(new_n622), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(G63));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n883), .B2(new_n849), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n891), .B1(new_n923), .B2(new_n648), .ZN(new_n924));
  INV_X1    g738(.A(new_n922), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n456), .B1(new_n902), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n920), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n902), .A2(new_n648), .A3(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n901), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n930), .A2(KEYINPUT124), .A3(new_n926), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n919), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n924), .A2(new_n920), .A3(new_n927), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT124), .B1(new_n930), .B2(new_n926), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n935), .ZN(G66));
  OAI21_X1  g750(.A(G953), .B1(new_n303), .B2(new_n565), .ZN(new_n937));
  INV_X1    g751(.A(new_n196), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n836), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n588), .B(new_n556), .C1(G898), .C2(new_n196), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  AOI21_X1  g755(.A(new_n196), .B1(G227), .B2(G900), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n506), .B(new_n222), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(G900), .B2(new_n938), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n746), .A2(new_n697), .A3(new_n727), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n763), .A2(new_n729), .A3(new_n817), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n756), .A2(new_n945), .A3(new_n735), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n944), .B1(new_n947), .B2(new_n938), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n942), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n832), .A2(new_n713), .A3(new_n663), .A4(new_n541), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT126), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n951), .A2(KEYINPUT126), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n952), .B(new_n953), .C1(new_n747), .C2(new_n755), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n675), .A2(new_n817), .ZN(new_n955));
  AND2_X1   g769(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n956));
  NOR2_X1   g770(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n958), .B(new_n763), .C1(new_n955), .C2(new_n956), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n943), .B1(new_n960), .B2(new_n938), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n948), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n950), .B(new_n962), .Z(G72));
  NAND2_X1  g777(.A1(new_n530), .A2(new_n519), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n947), .A2(new_n497), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(new_n836), .C1(new_n507), .C2(new_n960), .ZN(new_n966));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  AOI21_X1  g782(.A(new_n964), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n863), .A2(new_n968), .A3(new_n964), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n891), .A3(new_n970), .ZN(G57));
endmodule


