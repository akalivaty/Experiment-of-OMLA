//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(G58), .A2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n229), .A2(G50), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n231), .A2(new_n204), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n206), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT0), .Z(new_n236));
  NOR3_X1   g0036(.A1(new_n226), .A2(new_n233), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n214), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n219), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n232), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n204), .A2(G1), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G77), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT15), .B(G87), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n204), .A2(G33), .ZN(new_n262));
  OR3_X1    g0062(.A1(new_n261), .A2(KEYINPUT69), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT8), .B(G58), .Z(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT69), .B1(new_n261), .B2(new_n262), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n257), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n255), .B(new_n260), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G238), .A2(G1698), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n272), .B(new_n273), .C1(new_n223), .C2(G1698), .ZN(new_n274));
  AND2_X1   g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n274), .B(new_n278), .C1(G107), .C2(new_n272), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT65), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n283), .A2(new_n284), .A3(new_n232), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT65), .B1(new_n275), .B2(new_n276), .ZN(new_n286));
  OAI211_X1 g0086(.A(G274), .B(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n283), .B2(new_n232), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n275), .A2(KEYINPUT65), .A3(new_n276), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n282), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n279), .B(new_n287), .C1(new_n220), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n271), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n271), .A2(KEYINPUT71), .A3(new_n294), .A4(new_n295), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n293), .A2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n270), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT67), .B1(new_n258), .B2(new_n217), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT67), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(G50), .C1(new_n204), .C2(G1), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n308), .A2(new_n269), .A3(new_n253), .A4(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(G50), .B2(new_n253), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT68), .ZN(new_n313));
  INV_X1    g0113(.A(new_n264), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n262), .ZN(new_n315));
  OAI21_X1  g0115(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n316));
  INV_X1    g0116(.A(G150), .ZN(new_n317));
  INV_X1    g0117(.A(new_n265), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n257), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT66), .A2(G223), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT66), .A2(G223), .ZN(new_n323));
  OAI21_X1  g0123(.A(G1698), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G222), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n272), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n278), .C1(G77), .C2(new_n272), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n287), .C1(new_n218), .C2(new_n292), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n304), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n321), .B(new_n330), .C1(G179), .C2(new_n329), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n321), .A2(KEYINPUT9), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n321), .A2(KEYINPUT9), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(G200), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n329), .A2(new_n299), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n335), .A2(KEYINPUT72), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT10), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n333), .B2(new_n334), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n336), .A4(new_n337), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n332), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G33), .ZN(new_n346));
  OR2_X1    g0146(.A1(G223), .A2(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G33), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n218), .A2(G1698), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n346), .A2(new_n347), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G87), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n278), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT82), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n277), .B1(new_n351), .B2(new_n352), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT82), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(G232), .B(new_n291), .C1(new_n285), .C2(new_n286), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n287), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT83), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT83), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n287), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n359), .A2(new_n299), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n287), .A2(new_n360), .A3(new_n363), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n363), .B1(new_n287), .B2(new_n360), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n366), .A2(new_n367), .A3(new_n356), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n365), .B1(new_n368), .B2(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n314), .A2(new_n253), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n259), .B2(new_n314), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  INV_X1    g0173(.A(G68), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT80), .ZN(new_n375));
  AOI21_X1  g0175(.A(G20), .B1(new_n346), .B2(new_n349), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT80), .B(new_n378), .C1(new_n272), .C2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT81), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n346), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n349), .B1(new_n346), .B2(new_n381), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT7), .B(new_n204), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n374), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n222), .A2(new_n374), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n227), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n265), .A2(G159), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n373), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n378), .B1(new_n272), .B2(G20), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n394), .B2(G68), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n269), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n372), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n369), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT84), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(KEYINPUT17), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n369), .B2(new_n397), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT85), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n402), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n391), .A2(new_n396), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n371), .ZN(new_n407));
  INV_X1    g0207(.A(G200), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n362), .A2(new_n364), .A3(new_n354), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n366), .A2(new_n367), .ZN(new_n410));
  AOI21_X1  g0210(.A(G190), .B1(new_n355), .B2(new_n358), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n405), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT85), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n369), .A2(new_n397), .A3(new_n399), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(G179), .B1(new_n355), .B2(new_n358), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n304), .A2(new_n409), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n407), .A2(KEYINPUT18), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(new_n417), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G169), .B2(new_n368), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n420), .B1(new_n422), .B2(new_n397), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n404), .A2(new_n416), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n318), .A2(new_n217), .B1(new_n204), .B2(G68), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n262), .A2(new_n219), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n257), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT11), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n253), .A2(KEYINPUT12), .A3(G68), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT12), .B1(new_n253), .B2(G68), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n431), .A2(new_n432), .B1(new_n259), .B2(G68), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT77), .ZN(new_n435));
  OAI211_X1 g0235(.A(G238), .B(new_n291), .C1(new_n285), .C2(new_n286), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n287), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n218), .A2(new_n325), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n223), .A2(G1698), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n272), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G97), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n277), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT13), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT74), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n278), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT13), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n287), .A4(new_n436), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT73), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n437), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT73), .A3(new_n447), .A4(new_n446), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT74), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(KEYINPUT13), .C1(new_n437), .C2(new_n442), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n444), .A2(new_n450), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT78), .A3(G169), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT14), .ZN(new_n457));
  INV_X1    g0257(.A(G179), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT76), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n443), .A2(new_n459), .A3(new_n448), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n451), .A2(KEYINPUT76), .A3(new_n447), .A4(new_n446), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n455), .A2(KEYINPUT78), .A3(new_n465), .A4(G169), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n457), .A2(new_n463), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n455), .A2(G200), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n468), .B(KEYINPUT75), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n299), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n435), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n435), .A2(new_n467), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n307), .A2(new_n344), .A3(new_n426), .A4(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n346), .A2(new_n349), .A3(G244), .A4(new_n325), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT86), .A2(KEYINPUT4), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n475), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n272), .A2(G244), .A3(new_n325), .A4(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(KEYINPUT86), .A2(KEYINPUT4), .B1(G33), .B2(G283), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n278), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n203), .A2(G45), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n288), .A2(new_n289), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G257), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n485), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(new_n290), .A3(G274), .A4(new_n282), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n482), .A2(new_n458), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT87), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n254), .A2(new_n209), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n203), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n253), .A2(new_n495), .A3(new_n232), .A4(new_n256), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G97), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n213), .B1(new_n380), .B2(new_n385), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n209), .A2(new_n213), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n204), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n318), .A2(new_n219), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n499), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n494), .B(new_n498), .C1(new_n508), .C2(new_n269), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n482), .A2(new_n487), .A3(new_n490), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n304), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n493), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n505), .A2(new_n204), .ZN(new_n513));
  INV_X1    g0313(.A(new_n507), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n345), .A2(G33), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(KEYINPUT81), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(G20), .B1(new_n517), .B2(new_n382), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(KEYINPUT7), .B1(new_n377), .B2(new_n379), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n513), .B(new_n514), .C1(new_n519), .C2(new_n213), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n257), .B1(G97), .B2(new_n497), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n510), .A2(G200), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n482), .A2(new_n487), .A3(new_n490), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G190), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n521), .A2(new_n494), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n512), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n346), .A2(new_n349), .A3(new_n204), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n272), .A2(new_n529), .A3(new_n204), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n204), .A2(G107), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n532), .B(KEYINPUT23), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n531), .A2(KEYINPUT24), .A3(new_n533), .A4(new_n534), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n257), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n497), .A2(G107), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n253), .A2(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT25), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n208), .A2(new_n325), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n210), .A2(G1698), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n272), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n278), .A2(new_n548), .B1(new_n486), .B2(G264), .ZN(new_n549));
  AOI21_X1  g0349(.A(G169), .B1(new_n549), .B2(new_n490), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n490), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n552), .B2(new_n458), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n543), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT21), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n253), .A2(G116), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n496), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(G33), .B2(G283), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G33), .B2(new_n209), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(G20), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n257), .A2(KEYINPUT91), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT91), .B1(new_n257), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT20), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(KEYINPUT20), .B(new_n560), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n556), .B(new_n558), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n486), .A2(G270), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n346), .A2(new_n349), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G264), .A2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n210), .B2(G1698), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n278), .C1(new_n570), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n490), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G169), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n555), .B1(new_n568), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n566), .A2(new_n567), .ZN(new_n579));
  INV_X1    g0379(.A(new_n556), .ZN(new_n580));
  INV_X1    g0380(.A(new_n558), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(KEYINPUT21), .A3(G169), .A4(new_n576), .ZN(new_n583));
  INV_X1    g0383(.A(new_n576), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G190), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n576), .A2(G200), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n568), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(G179), .A3(new_n584), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n578), .A2(new_n583), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n552), .A2(new_n408), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n551), .A2(new_n299), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n543), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n207), .A2(new_n209), .A3(new_n213), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n441), .A2(new_n204), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT19), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n346), .A2(new_n349), .A3(new_n204), .A4(G68), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n441), .B2(G20), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n257), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n261), .A2(new_n254), .ZN(new_n601));
  INV_X1    g0401(.A(new_n261), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT89), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n496), .B2(new_n261), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n600), .A2(new_n601), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n208), .A2(KEYINPUT88), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n485), .B1(new_n607), .B2(G274), .ZN(new_n608));
  OAI211_X1 g0408(.A(KEYINPUT88), .B(G250), .C1(new_n281), .C2(G1), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n608), .A2(new_n609), .B1(new_n288), .B2(new_n289), .ZN(new_n610));
  OR2_X1    g0410(.A1(G238), .A2(G1698), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n220), .A2(G1698), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n346), .A2(new_n611), .A3(new_n349), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G33), .A2(G116), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n277), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n304), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n615), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT88), .ZN(new_n618));
  AOI21_X1  g0418(.A(G274), .B1(new_n618), .B2(G250), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n609), .B1(new_n619), .B2(new_n484), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n290), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n458), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n606), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(G200), .B1(new_n610), .B2(new_n615), .ZN(new_n624));
  NOR2_X1   g0424(.A1(G238), .A2(G1698), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n220), .B2(G1698), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n272), .B1(G33), .B2(G116), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n621), .B(G190), .C1(new_n627), .C2(new_n277), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n599), .A2(new_n257), .B1(new_n261), .B2(new_n254), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n497), .A2(G87), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n624), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n623), .A2(new_n631), .A3(KEYINPUT90), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n589), .A2(new_n592), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n473), .A2(new_n526), .A3(new_n554), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g0438(.A(new_n638), .B(KEYINPUT92), .Z(G372));
  AND2_X1   g0439(.A1(new_n467), .A2(new_n435), .ZN(new_n640));
  INV_X1    g0440(.A(new_n306), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n469), .A2(new_n471), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n404), .A2(new_n416), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n424), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n339), .A2(new_n343), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n332), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT26), .B1(new_n512), .B2(new_n636), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n290), .A2(KEYINPUT93), .A3(new_n620), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT93), .B1(new_n290), .B2(new_n620), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n617), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n304), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n606), .A2(new_n622), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n554), .A2(new_n588), .A3(new_n583), .A4(new_n578), .ZN(new_n656));
  INV_X1    g0456(.A(new_n592), .ZN(new_n657));
  INV_X1    g0457(.A(new_n511), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n521), .B2(new_n494), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n656), .A2(new_n657), .B1(new_n659), .B2(new_n493), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n629), .A2(new_n630), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n610), .A2(new_n615), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(G190), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n652), .A2(G200), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n525), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n648), .B(new_n655), .C1(new_n660), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n473), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n647), .A2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n578), .A2(new_n583), .A3(new_n588), .ZN(new_n671));
  INV_X1    g0471(.A(G13), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G20), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n232), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT94), .ZN(new_n676));
  INV_X1    g0476(.A(G213), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(KEYINPUT94), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n568), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n671), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n589), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n554), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n543), .A2(new_n682), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n657), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n691), .B2(new_n554), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n671), .A2(new_n683), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n689), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n234), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n593), .A2(G116), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n231), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n656), .A2(new_n657), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n666), .A2(new_n655), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n512), .A2(new_n525), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n493), .A2(new_n509), .A3(new_n511), .A4(new_n666), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n623), .A2(new_n631), .A3(KEYINPUT90), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT90), .B1(new_n623), .B2(new_n631), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n659), .A2(new_n712), .A3(new_n661), .A4(new_n493), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n713), .A3(new_n655), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n683), .B1(new_n707), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT96), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n683), .C1(new_n707), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n668), .A2(new_n683), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT95), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT95), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n668), .A2(new_n724), .A3(new_n683), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n637), .A2(new_n526), .A3(new_n554), .A4(new_n683), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n584), .A2(G179), .A3(new_n549), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n482), .A2(new_n663), .A3(new_n487), .A4(new_n490), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n549), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n490), .A2(new_n569), .A3(new_n575), .A4(G179), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n523), .A3(KEYINPUT30), .A4(new_n663), .ZN(new_n736));
  AOI21_X1  g0536(.A(G179), .B1(new_n651), .B2(new_n617), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n510), .A3(new_n551), .A4(new_n576), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n682), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n728), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n727), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n703), .B1(new_n746), .B2(G1), .ZN(G364));
  NAND3_X1  g0547(.A1(new_n234), .A2(G355), .A3(new_n272), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n697), .A2(new_n272), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G45), .B2(new_n231), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n248), .A2(new_n281), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n748), .B1(G116), .B2(new_n234), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(G20), .B1(KEYINPUT97), .B2(G169), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(KEYINPUT97), .A2(G169), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n232), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n204), .A2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n408), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G283), .A2(new_n765), .B1(new_n768), .B2(G329), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n458), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G326), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n458), .A2(new_n408), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n204), .A2(new_n299), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n769), .B1(new_n770), .B2(new_n772), .C1(new_n773), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n763), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n272), .B(new_n777), .C1(G303), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n774), .A2(new_n762), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G317), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT33), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(KEYINPUT33), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n775), .A2(new_n771), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G322), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n766), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G294), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n780), .A2(new_n786), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n374), .A2(new_n781), .B1(new_n778), .B2(new_n207), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G97), .B2(new_n791), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n765), .A2(G107), .ZN(new_n796));
  INV_X1    g0596(.A(new_n776), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G50), .A2(new_n797), .B1(new_n788), .B2(G58), .ZN(new_n798));
  INV_X1    g0598(.A(new_n772), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n570), .B1(new_n799), .B2(G77), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n795), .A2(new_n796), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n768), .A2(G159), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n793), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT98), .Z(new_n805));
  AOI21_X1  g0605(.A(new_n761), .B1(new_n805), .B2(new_n756), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n673), .A2(G45), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n699), .A2(G1), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n759), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n806), .B(new_n809), .C1(new_n686), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n688), .A2(new_n809), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G330), .B2(new_n686), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NOR2_X1   g0615(.A1(new_n306), .A2(new_n682), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n270), .A2(new_n682), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n302), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n818), .B2(new_n306), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n722), .A2(new_n725), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n668), .A2(new_n307), .A3(new_n683), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT100), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n745), .B(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n809), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT100), .B1(new_n744), .B2(G330), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n820), .A2(new_n757), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n756), .A2(new_n757), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n219), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G50), .A2(new_n779), .B1(new_n765), .B2(G68), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT99), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G143), .A2(new_n788), .B1(new_n799), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(new_n836), .B2(new_n776), .C1(new_n317), .C2(new_n781), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n832), .A2(new_n833), .B1(G132), .B2(new_n768), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(new_n272), .A3(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n834), .B(new_n840), .C1(G58), .C2(new_n791), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n764), .A2(new_n207), .ZN(new_n842));
  INV_X1    g0642(.A(new_n791), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n570), .B1(new_n778), .B2(new_n213), .C1(new_n843), .C2(new_n209), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n842), .B(new_n844), .C1(G311), .C2(new_n768), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n797), .A2(G303), .B1(new_n799), .B2(G116), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(new_n846), .C1(new_n847), .C2(new_n781), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G294), .B2(new_n788), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n756), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n829), .A2(new_n809), .A3(new_n831), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n828), .A2(new_n851), .ZN(G384));
  NAND3_X1  g0652(.A1(new_n419), .A2(new_n423), .A3(new_n680), .ZN(new_n853));
  INV_X1    g0653(.A(new_n816), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n822), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n467), .A2(new_n435), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n435), .A2(new_n682), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n642), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n467), .A2(new_n435), .A3(new_n682), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT7), .B1(new_n570), .B2(new_n204), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n378), .B(G20), .C1(new_n346), .C2(new_n349), .ZN(new_n864));
  OAI21_X1  g0664(.A(G68), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n390), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(KEYINPUT16), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n257), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n519), .B2(new_n374), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n373), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n418), .B1(new_n870), .B2(new_n372), .ZN(new_n871));
  INV_X1    g0671(.A(new_n680), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n870), .B2(new_n372), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n369), .A2(new_n397), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n371), .B1(new_n868), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n418), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n872), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n874), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n880), .ZN(new_n883));
  AOI221_X4 g0683(.A(new_n862), .B1(new_n876), .B2(new_n882), .C1(new_n425), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n425), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n876), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT101), .B(new_n853), .C1(new_n861), .C2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n853), .B1(new_n861), .B2(new_n888), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n873), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n422), .A2(new_n397), .A3(new_n420), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT18), .B1(new_n407), .B2(new_n418), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n894), .A2(new_n895), .B1(new_n400), .B2(new_n403), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n893), .A2(new_n896), .B1(new_n898), .B2(new_n876), .ZN(new_n899));
  XNOR2_X1  g0699(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT103), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT103), .ZN(new_n903));
  INV_X1    g0703(.A(new_n900), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n898), .A2(new_n876), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n413), .A2(new_n415), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n873), .B1(new_n906), .B2(new_n424), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n901), .A2(new_n902), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT104), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT39), .B1(new_n884), .B2(new_n887), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT104), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n856), .A2(new_n682), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n889), .B(new_n892), .C1(new_n915), .C2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n720), .A2(new_n726), .A3(new_n473), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n647), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n740), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n739), .A2(KEYINPUT105), .A3(new_n682), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n741), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n728), .A2(new_n925), .A3(new_n743), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n473), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT106), .Z(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n819), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n472), .A2(new_n857), .B1(new_n640), .B2(new_n682), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n901), .A2(new_n902), .A3(new_n908), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n860), .A2(new_n929), .A3(new_n819), .A4(new_n926), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n888), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n928), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(G330), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n921), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n203), .B2(new_n673), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT35), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n204), .B(new_n232), .C1(new_n505), .C2(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n943), .B(G116), .C1(new_n942), .C2(new_n505), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT36), .ZN(new_n945));
  OAI21_X1  g0745(.A(G77), .B1(new_n222), .B2(new_n374), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n231), .A2(new_n946), .B1(G50), .B2(new_n374), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(G1), .A3(new_n672), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n941), .A2(new_n945), .A3(new_n948), .ZN(G367));
  INV_X1    g0749(.A(new_n749), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n760), .B1(new_n234), .B2(new_n261), .C1(new_n244), .C2(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n776), .A2(new_n770), .B1(new_n787), .B2(new_n571), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT113), .Z(new_n953));
  NAND2_X1  g0753(.A1(new_n779), .A2(G116), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT46), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n954), .A2(new_n955), .B1(new_n791), .B2(G107), .ZN(new_n956));
  INV_X1    g0756(.A(G294), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n953), .B(new_n956), .C1(new_n957), .C2(new_n781), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n570), .B1(new_n767), .B2(new_n783), .C1(new_n209), .C2(new_n764), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT114), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(new_n847), .C2(new_n772), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n954), .A2(new_n955), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n843), .A2(new_n374), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n772), .A2(new_n217), .B1(new_n767), .B2(new_n836), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n765), .A2(G77), .ZN(new_n966));
  INV_X1    g0766(.A(G159), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(new_n967), .B2(new_n781), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n965), .B(new_n968), .C1(G58), .C2(new_n779), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n570), .B1(new_n797), .B2(G143), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n317), .C2(new_n787), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT47), .Z(new_n973));
  INV_X1    g0773(.A(new_n756), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n809), .B(new_n951), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n682), .A2(new_n662), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT107), .Z(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(new_n654), .A3(new_n653), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT108), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n705), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n978), .B(new_n979), .C1(new_n981), .C2(new_n977), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n975), .B1(new_n759), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n692), .A2(new_n694), .ZN(new_n985));
  INV_X1    g0785(.A(new_n526), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n985), .A2(KEYINPUT42), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT42), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n526), .A2(new_n554), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n525), .A3(new_n683), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n983), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT109), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n980), .A2(new_n982), .A3(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n991), .A2(new_n993), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT110), .ZN(new_n999));
  INV_X1    g0799(.A(new_n693), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n509), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n526), .B1(new_n1001), .B2(new_n683), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n659), .A2(new_n493), .A3(new_n682), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n996), .A2(new_n999), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n998), .B(KEYINPUT110), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1006), .A2(new_n995), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n807), .A2(G1), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n692), .B(new_n694), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT112), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n688), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1000), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n695), .A2(new_n1004), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(KEYINPUT111), .B2(KEYINPUT44), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT111), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT44), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n695), .C2(new_n1004), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1018), .B(new_n1021), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n695), .A2(new_n1004), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT45), .Z(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n746), .A2(new_n1016), .A3(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1026), .A2(new_n746), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n698), .B(KEYINPUT41), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1011), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n984), .B1(new_n1009), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(G387));
  NOR2_X1   g0832(.A1(new_n746), .A2(new_n1016), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n746), .A2(new_n1016), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n698), .B(KEYINPUT115), .Z(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n772), .A2(new_n374), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n843), .A2(new_n261), .B1(new_n317), .B2(new_n767), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G50), .C2(new_n788), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n797), .A2(G159), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G77), .A2(new_n779), .B1(new_n765), .B2(G97), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n570), .B1(new_n782), .B2(new_n264), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G322), .A2(new_n797), .B1(new_n782), .B2(G311), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n571), .B2(new_n772), .C1(new_n783), .C2(new_n787), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT48), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n847), .B2(new_n843), .C1(new_n957), .C2(new_n778), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT49), .Z(new_n1050));
  OAI221_X1 g0850(.A(new_n570), .B1(new_n767), .B2(new_n773), .C1(new_n557), .C2(new_n764), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1045), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n756), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n809), .C1(new_n692), .C2(new_n810), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n264), .A2(new_n217), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT50), .Z(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n281), .C1(new_n374), .C2(new_n219), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n700), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n749), .B1(new_n241), .B2(new_n281), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n234), .A3(new_n272), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n234), .A2(G107), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n760), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1055), .A2(new_n1065), .B1(new_n1016), .B2(new_n1010), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1038), .A2(new_n1066), .ZN(G393));
  NAND2_X1  g0867(.A1(new_n1025), .A2(new_n1000), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1022), .A2(new_n1024), .A3(new_n693), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n1035), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n1026), .A3(new_n1037), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT116), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1026), .A3(new_n1074), .A4(new_n1037), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1002), .A2(new_n759), .A3(new_n1003), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n776), .A2(new_n783), .B1(new_n787), .B2(new_n770), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G303), .B2(new_n782), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n799), .A2(G294), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n768), .A2(G322), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n796), .B1(new_n847), .B2(new_n778), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n272), .B(new_n1082), .C1(G116), .C2(new_n791), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n776), .A2(new_n317), .B1(new_n787), .B2(new_n967), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  OAI22_X1  g0886(.A1(new_n314), .A2(new_n772), .B1(new_n374), .B2(new_n778), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1086), .A2(new_n842), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n782), .A2(G50), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n768), .A2(G143), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n570), .B1(new_n791), .B2(G77), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n974), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n749), .A2(new_n251), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n759), .B(new_n756), .C1(new_n697), .C2(G97), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n808), .B(new_n1093), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1073), .A2(new_n1075), .B1(new_n1076), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1068), .A2(new_n1010), .A3(new_n1069), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(G390));
  AND2_X1   g0899(.A1(new_n901), .A2(new_n902), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1100), .A2(KEYINPUT104), .A3(new_n909), .A4(new_n908), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n861), .A2(new_n917), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n885), .A2(new_n886), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n862), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n902), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n911), .B1(new_n1105), .B2(KEYINPUT39), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n910), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1101), .B(new_n1102), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n860), .A2(G330), .A3(new_n744), .A4(new_n819), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n716), .A2(new_n718), .A3(new_n854), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n818), .A2(new_n306), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n860), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n933), .A3(new_n917), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1108), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1110), .A2(new_n1111), .A3(new_n860), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n933), .A2(new_n917), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n915), .B2(new_n1102), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n860), .A2(G330), .A3(new_n819), .A4(new_n926), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n1011), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n915), .A2(new_n757), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT54), .B(G143), .Z(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n772), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n779), .A2(G150), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  INV_X1    g0927(.A(G132), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n272), .B1(new_n781), .B2(new_n836), .C1(new_n1128), .C2(new_n787), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G50), .A2(new_n765), .B1(new_n768), .B2(G125), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n967), .C2(new_n843), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1125), .B(new_n1132), .C1(G128), .C2(new_n797), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n772), .A2(new_n209), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G87), .A2(new_n779), .B1(new_n765), .B2(G68), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n797), .A2(G283), .B1(new_n768), .B2(G294), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n782), .A2(G107), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n272), .B1(new_n791), .B2(G77), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1134), .B(new_n1139), .C1(G116), .C2(new_n788), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n756), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1122), .A2(new_n809), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n314), .B2(new_n830), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1121), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n473), .A2(G330), .A3(new_n926), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n919), .A2(new_n647), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n926), .A2(G330), .A3(new_n819), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1110), .A2(new_n1111), .B1(new_n931), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1109), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n931), .B1(new_n745), .B2(new_n820), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1119), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n855), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1120), .A2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1109), .A2(new_n1149), .B1(new_n1152), .B2(new_n855), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n1146), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1114), .B(new_n1158), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n1037), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1144), .A2(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(KEYINPUT120), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1101), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n916), .B1(new_n891), .B2(new_n890), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n344), .A2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n332), .B(new_n1165), .C1(new_n339), .C2(new_n343), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n321), .A2(new_n872), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n344), .A2(new_n1166), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1170), .B1(new_n1173), .B2(new_n1168), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(G330), .C1(new_n934), .C2(new_n936), .ZN(new_n1176));
  OAI21_X1  g0976(.A(G330), .B1(new_n934), .B2(new_n936), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1164), .A2(new_n889), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1176), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n918), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1147), .A2(new_n1159), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1162), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1159), .A2(new_n1147), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(KEYINPUT120), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1180), .A2(new_n1182), .A3(KEYINPUT119), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT119), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1181), .A2(new_n918), .A3(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n1185), .A3(KEYINPUT57), .A4(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1184), .A2(new_n1189), .A3(new_n1037), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n830), .A2(new_n217), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G41), .B(new_n272), .C1(new_n765), .C2(G58), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n219), .B2(new_n778), .C1(new_n847), .C2(new_n767), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT117), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n772), .A2(new_n261), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n787), .A2(new_n213), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT118), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1198), .A2(new_n964), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n209), .B2(new_n781), .C1(new_n557), .C2(new_n776), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT58), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n772), .A2(new_n836), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n843), .A2(new_n317), .B1(new_n1124), .B2(new_n778), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G128), .C2(new_n788), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n797), .A2(G125), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n1128), .C2(new_n781), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT59), .Z(new_n1210));
  INV_X1    g1010(.A(G124), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n348), .B(new_n280), .C1(new_n767), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G159), .B2(new_n765), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n280), .B1(new_n345), .B2(new_n348), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1210), .A2(new_n1213), .B1(new_n217), .B2(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1204), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n809), .B(new_n1195), .C1(new_n1216), .C2(new_n974), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1178), .B2(new_n757), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1186), .B2(new_n1010), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1194), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1157), .A2(new_n1146), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT121), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT121), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1157), .A2(new_n1146), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n1028), .A3(new_n1155), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1010), .B(KEYINPUT122), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n931), .A2(new_n757), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G159), .A2(new_n779), .B1(new_n765), .B2(G58), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n1128), .B2(new_n776), .C1(new_n317), .C2(new_n772), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n570), .B(new_n1230), .C1(G128), .C2(new_n768), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n217), .B2(new_n843), .C1(new_n781), .C2(new_n1124), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G137), .B2(new_n788), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n966), .B1(new_n213), .B2(new_n772), .C1(new_n557), .C2(new_n781), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G283), .B2(new_n788), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n843), .A2(new_n261), .B1(new_n778), .B2(new_n209), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n272), .B(new_n1236), .C1(G294), .C2(new_n797), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1235), .B(new_n1237), .C1(new_n571), .C2(new_n767), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT123), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n756), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n830), .A2(new_n374), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1228), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1154), .A2(new_n1227), .B1(new_n809), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1226), .A2(new_n1243), .ZN(G381));
  NOR2_X1   g1044(.A1(G375), .A2(G378), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(G381), .A2(G384), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1097), .A2(new_n1031), .A3(new_n1098), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(G407));
  AOI21_X1  g1049(.A(new_n677), .B1(new_n1245), .B2(new_n681), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(G407), .ZN(G409));
  AOI21_X1  g1051(.A(new_n814), .B1(new_n1038), .B2(new_n1066), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1031), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1247), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G390), .A2(G387), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1253), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1097), .A2(new_n1031), .A3(new_n1098), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1222), .A2(new_n1224), .B1(new_n1155), .B2(KEYINPUT60), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1037), .B1(new_n1221), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1243), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(G384), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G384), .B(new_n1243), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n677), .A2(G343), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT124), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(G2897), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1266), .A2(new_n1271), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1273), .A2(KEYINPUT125), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT125), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1194), .A2(G378), .A3(new_n1219), .ZN(new_n1278));
  INV_X1    g1078(.A(G378), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1190), .A2(new_n1192), .A3(new_n1227), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1187), .B2(new_n1029), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1279), .B1(new_n1281), .B2(new_n1218), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1268), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1260), .B1(new_n1277), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1268), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1286), .B(new_n1287), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1288), .A2(new_n1295), .A3(new_n1291), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1287), .B1(new_n1288), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1296), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1260), .B(KEYINPUT126), .Z(new_n1301));
  OAI21_X1  g1101(.A(new_n1294), .B1(new_n1300), .B2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1279), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1278), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(G375), .A2(KEYINPUT127), .A3(new_n1279), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1305), .A2(new_n1260), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1260), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1290), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1260), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1278), .A2(new_n1304), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G378), .B1(new_n1194), .B2(new_n1219), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1306), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1310), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1305), .A2(new_n1260), .A3(new_n1306), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1291), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1309), .A2(new_n1317), .ZN(G402));
endmodule


