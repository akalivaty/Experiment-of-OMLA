//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G141gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n214));
  OAI211_X1 g013(.A(KEYINPUT74), .B(new_n208), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n208), .A2(KEYINPUT74), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT74), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n206), .A2(new_n217), .A3(new_n207), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n210), .A2(new_n212), .B1(KEYINPUT2), .B2(new_n207), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222));
  XNOR2_X1  g021(.A(G211gat), .B(G218gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT71), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT69), .B(G211gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT70), .B(G218gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G197gat), .B(G204gat), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n226), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT22), .B1(new_n227), .B2(new_n228), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n235), .A2(new_n225), .A3(new_n232), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n222), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT75), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(new_n226), .A3(new_n233), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n225), .B1(new_n235), .B2(new_n232), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT29), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT75), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n221), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n234), .A2(new_n236), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G228gat), .ZN(new_n251));
  INV_X1    g050(.A(G233gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT76), .B1(new_n244), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n221), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n237), .A2(new_n238), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n245), .B1(new_n242), .B2(KEYINPUT75), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n250), .A2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT76), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n223), .B1(new_n235), .B2(new_n232), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n247), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n235), .A2(new_n223), .A3(new_n232), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n245), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n256), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n253), .B1(new_n268), .B2(new_n250), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n203), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  AOI211_X1 g070(.A(G22gat), .B(new_n269), .C1(new_n255), .C2(new_n262), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n244), .A2(KEYINPUT76), .A3(new_n254), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n261), .B1(new_n259), .B2(new_n260), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G22gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n263), .A2(new_n203), .A3(new_n270), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G78gat), .B(G106gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT31), .B(G50gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n278), .A4(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G113gat), .B2(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(G113gat), .A2(G120gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G127gat), .ZN(new_n293));
  INV_X1    g092(.A(G127gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n287), .B(new_n294), .C1(new_n289), .C2(new_n291), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(G134gat), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(G134gat), .B1(new_n293), .B2(new_n295), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n221), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n215), .A2(new_n220), .A3(KEYINPUT3), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n246), .A3(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n298), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n307), .A2(new_n296), .B1(new_n215), .B2(new_n220), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT4), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n305), .A2(KEYINPUT5), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n306), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n297), .A2(new_n221), .A3(new_n298), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT5), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n309), .A2(new_n301), .A3(new_n304), .A4(new_n306), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT0), .ZN(new_n319));
  XNOR2_X1  g118(.A(G57gat), .B(G85gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  AOI21_X1  g120(.A(KEYINPUT6), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n310), .A2(new_n316), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n310), .A2(new_n316), .A3(KEYINPUT6), .A4(new_n323), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT27), .B(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n334));
  OR2_X1    g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n334), .ZN(new_n336));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(G169gat), .ZN(new_n338));
  INV_X1    g137(.A(G176gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n340), .A2(KEYINPUT26), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(KEYINPUT26), .ZN(new_n342));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n337), .ZN(new_n347));
  NAND3_X1  g146(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n343), .A2(KEYINPUT23), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n340), .ZN(new_n351));
  OR2_X1    g150(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n349), .B(new_n351), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT66), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n355), .A2(G176gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n357), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n348), .B(KEYINPUT65), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n346), .A2(new_n337), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n361), .B(new_n351), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n358), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n359), .B1(new_n358), .B2(new_n364), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n330), .B(new_n345), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(new_n364), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n345), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n222), .A3(new_n329), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n249), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n330), .A3(new_n345), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n345), .B1(new_n365), .B2(new_n366), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n247), .A2(new_n329), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n371), .B1(new_n249), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  OAI21_X1  g180(.A(new_n328), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n371), .ZN(new_n383));
  INV_X1    g182(.A(new_n345), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n368), .A2(KEYINPUT66), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n359), .A3(new_n364), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n249), .B(new_n372), .C1(new_n387), .C2(new_n375), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n381), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n378), .A2(new_n392), .A3(new_n381), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n383), .A2(new_n388), .A3(new_n381), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT30), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n382), .A2(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n327), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n286), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT38), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT37), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n372), .B1(new_n387), .B2(new_n375), .ZN(new_n401));
  INV_X1    g200(.A(new_n249), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT79), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n367), .A2(new_n249), .A3(new_n370), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(KEYINPUT79), .A3(new_n402), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n400), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n390), .B1(new_n389), .B2(KEYINPUT37), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n399), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n400), .B1(new_n383), .B2(new_n388), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT80), .B1(new_n410), .B2(new_n381), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n412), .B(new_n390), .C1(new_n378), .C2(new_n400), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n399), .B1(new_n378), .B2(new_n400), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n325), .A2(new_n326), .A3(new_n394), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT78), .B(KEYINPUT39), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n301), .A2(new_n304), .ZN(new_n419));
  INV_X1    g218(.A(new_n309), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n311), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n306), .B1(new_n305), .B2(new_n309), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n308), .A2(new_n312), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT39), .B1(new_n423), .B2(new_n311), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n421), .B(new_n321), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT40), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n427), .A2(new_n324), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n396), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n416), .A2(new_n417), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n284), .A2(new_n285), .ZN(new_n432));
  INV_X1    g231(.A(new_n302), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n374), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G227gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n252), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n302), .B(new_n345), .C1(new_n365), .C2(new_n366), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n438), .A2(KEYINPUT32), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G15gat), .B(G43gat), .Z(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n436), .B1(new_n434), .B2(new_n437), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT34), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI211_X1 g247(.A(KEYINPUT34), .B(new_n436), .C1(new_n434), .C2(new_n437), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n444), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n438), .B2(new_n440), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n446), .A2(new_n447), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n449), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n439), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n451), .A2(new_n439), .A3(new_n455), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(KEYINPUT36), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n451), .A2(new_n439), .A3(new_n455), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n431), .A2(new_n432), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n327), .A2(new_n396), .A3(KEYINPUT81), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n461), .A2(new_n456), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n285), .A4(new_n284), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n432), .A2(new_n468), .A3(new_n465), .A4(new_n464), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n398), .A2(new_n463), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G113gat), .B(G141gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G197gat), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT11), .B(G169gat), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n474), .B(KEYINPUT12), .Z(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G8gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT16), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(G1gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n479), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT82), .B(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT83), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n488), .B(G36gat), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(G29gat), .A2(G36gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT14), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497));
  INV_X1    g296(.A(G50gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(G43gat), .ZN(new_n499));
  INV_X1    g298(.A(G43gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT84), .B1(new_n500), .B2(G50gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n498), .A2(G43gat), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n496), .B(new_n499), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n492), .A3(new_n495), .A4(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n500), .A2(G50gat), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n502), .A2(new_n505), .A3(new_n496), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n487), .A2(new_n506), .A3(new_n492), .A4(new_n495), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n508), .A2(KEYINPUT17), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT17), .B1(new_n508), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n484), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n479), .B(new_n482), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n509), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n512), .A2(KEYINPUT18), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n512), .A2(new_n517), .A3(new_n516), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n484), .A2(new_n514), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n516), .A3(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n517), .B(KEYINPUT13), .Z(new_n527));
  NAND3_X1  g326(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n514), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n475), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n518), .B(KEYINPUT86), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n523), .A2(new_n529), .ZN(new_n533));
  INV_X1    g332(.A(new_n475), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n470), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G190gat), .B(G218gat), .Z(new_n539));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT8), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(G85gat), .B2(G92gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n546));
  NOR2_X1   g345(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n544), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n548), .A2(KEYINPUT94), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT94), .B1(new_n548), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n543), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G99gat), .B(G106gat), .Z(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558));
  NAND2_X1  g357(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n544), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n547), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n548), .A2(KEYINPUT94), .A3(new_n552), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n556), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n565), .A3(new_n543), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n557), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n510), .B2(new_n511), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT95), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n567), .B(new_n570), .C1(new_n510), .C2(new_n511), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n567), .B2(new_n514), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n539), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT92), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n576), .B1(new_n569), .B2(new_n571), .ZN(new_n582));
  INV_X1    g381(.A(new_n539), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n587), .B(new_n586), .C1(new_n590), .C2(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(KEYINPUT91), .A3(new_n594), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT21), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n484), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n484), .ZN(new_n605));
  INV_X1    g404(.A(new_n597), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n596), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT20), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT89), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n604), .A2(new_n608), .A3(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n581), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n582), .A2(new_n583), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n539), .B(new_n576), .C1(new_n569), .C2(new_n571), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n585), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n585), .A2(new_n620), .A3(new_n624), .A4(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n565), .B1(new_n564), .B2(new_n543), .ZN(new_n630));
  AOI211_X1 g429(.A(new_n556), .B(new_n542), .C1(new_n562), .C2(new_n563), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT97), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n557), .A2(new_n633), .A3(new_n566), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n634), .A3(new_n595), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n630), .A2(new_n631), .ZN(new_n636));
  INV_X1    g435(.A(new_n595), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT10), .B1(new_n635), .B2(new_n638), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT98), .B1(new_n647), .B2(new_n643), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n639), .A2(new_n646), .ZN(new_n650));
  XOR2_X1   g449(.A(G120gat), .B(G148gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT99), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n647), .A2(new_n643), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n646), .B(KEYINPUT100), .Z(new_n660));
  OAI21_X1  g459(.A(new_n650), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n654), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n658), .B1(new_n657), .B2(new_n662), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n629), .A2(KEYINPUT102), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n657), .A2(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT101), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n626), .A2(new_n668), .A3(new_n628), .A4(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n538), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n327), .B(KEYINPUT103), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n430), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT16), .B(G8gat), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(G8gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n682), .A2(KEYINPUT104), .A3(new_n683), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(new_n674), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n459), .A2(new_n462), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n465), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n690), .B2(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n674), .A2(new_n286), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n620), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n585), .A2(new_n624), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AND4_X1   g500(.A1(new_n538), .A2(new_n699), .A3(new_n701), .A4(new_n665), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n485), .A3(new_n676), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n467), .A2(new_n469), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n431), .A2(new_n432), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n398), .A3(new_n691), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n700), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT106), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n711), .B(KEYINPUT44), .C1(new_n470), .C2(new_n700), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n286), .A2(new_n713), .A3(new_n397), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n398), .A2(KEYINPUT107), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n463), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n705), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n709), .A3(new_n701), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n710), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n536), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n531), .A2(KEYINPUT105), .A3(new_n535), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n668), .A2(new_n669), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n724), .A2(new_n620), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n719), .A2(new_n676), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n704), .B1(new_n485), .B2(new_n727), .ZN(G1328gat));
  NAND3_X1  g527(.A1(new_n702), .A2(new_n486), .A3(new_n430), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n719), .A2(new_n430), .A3(new_n726), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n486), .B2(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(new_n691), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n734), .A3(new_n726), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n702), .A2(new_n500), .A3(new_n465), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT47), .B1(new_n738), .B2(KEYINPUT109), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n740), .B(new_n741), .C1(new_n736), .C2(new_n737), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n739), .A2(new_n742), .ZN(G1330gat));
  NAND3_X1  g542(.A1(new_n702), .A2(new_n498), .A3(new_n286), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n719), .A2(new_n286), .A3(new_n726), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n498), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1331gat));
  AND4_X1   g547(.A1(new_n629), .A2(new_n717), .A3(new_n725), .A4(new_n724), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n676), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT110), .B(G57gat), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1332gat));
  AOI21_X1  g551(.A(new_n396), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT111), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1333gat));
  NAND2_X1  g556(.A1(new_n749), .A2(new_n734), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n693), .A2(G71gat), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n758), .A2(G71gat), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n749), .A2(new_n286), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n723), .A2(new_n620), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n717), .A2(new_n701), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n717), .A2(KEYINPUT51), .A3(new_n701), .A4(new_n764), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n665), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(G85gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n770), .A3(new_n676), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n723), .A2(new_n665), .A3(new_n620), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n719), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n676), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(new_n770), .ZN(G1336gat));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n430), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n396), .A2(G92gat), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(new_n769), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n767), .A2(KEYINPUT112), .A3(new_n768), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n782), .A3(new_n766), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n725), .A2(new_n778), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n776), .A2(G92gat), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n780), .B1(new_n786), .B2(new_n787), .ZN(G1337gat));
  AOI21_X1  g587(.A(G99gat), .B1(new_n769), .B2(new_n465), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n734), .A2(G99gat), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n773), .B2(new_n790), .ZN(G1338gat));
  NAND2_X1  g590(.A1(new_n767), .A2(new_n768), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n432), .A2(G106gat), .A3(new_n665), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT53), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n719), .A2(new_n286), .A3(new_n772), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G106gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n795), .A2(new_n801), .A3(G106gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n795), .B2(G106gat), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n781), .A2(new_n783), .A3(new_n793), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(G1339gat));
  NOR2_X1   g606(.A1(new_n670), .A2(new_n723), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n659), .B2(new_n660), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n649), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n660), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n809), .B(new_n812), .C1(new_n647), .C2(new_n643), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n654), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n657), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n814), .B1(new_n649), .B2(new_n810), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(KEYINPUT55), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n818), .A2(KEYINPUT55), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n818), .A2(KEYINPUT55), .B1(new_n649), .B2(new_n656), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n820), .A2(new_n824), .A3(new_n723), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n517), .B1(new_n512), .B2(new_n516), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n474), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n535), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n663), .B2(new_n664), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT116), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n725), .A2(new_n833), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n700), .B1(new_n825), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n820), .A2(new_n824), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n700), .A2(new_n829), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n808), .B1(new_n840), .B2(new_n699), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n675), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n693), .A2(new_n286), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n842), .A2(new_n396), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n723), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n841), .A2(new_n286), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n675), .A2(new_n430), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n465), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(G113gat), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(new_n537), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n845), .A2(new_n850), .ZN(G1340gat));
  AOI21_X1  g650(.A(G120gat), .B1(new_n844), .B2(new_n725), .ZN(new_n852));
  INV_X1    g651(.A(G120gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n848), .A2(new_n853), .A3(new_n665), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n852), .A2(new_n854), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n844), .A2(new_n294), .A3(new_n620), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n848), .B2(new_n699), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  INV_X1    g657(.A(G134gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n430), .A2(new_n700), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n842), .A2(new_n859), .A3(new_n843), .A4(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n848), .B2(new_n700), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(KEYINPUT117), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(KEYINPUT117), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n862), .B(new_n863), .C1(new_n865), .C2(new_n866), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n847), .A2(new_n691), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n808), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n820), .A2(new_n824), .A3(new_n723), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n832), .A3(new_n834), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n873), .A2(new_n700), .B1(new_n838), .B2(new_n837), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n874), .B2(new_n620), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n286), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n432), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n839), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n818), .B2(new_n882), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT119), .B(new_n814), .C1(new_n649), .C2(new_n810), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n536), .A2(new_n816), .A3(new_n657), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n831), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n700), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n699), .B1(new_n880), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n879), .B1(new_n889), .B2(new_n871), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n870), .B1(new_n876), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G141gat), .B1(new_n891), .B2(new_n537), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n691), .A2(new_n286), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT120), .Z(new_n895));
  NAND3_X1  g694(.A1(new_n842), .A2(new_n396), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n536), .A2(new_n209), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n676), .A3(new_n895), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n430), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n900), .A2(KEYINPUT122), .A3(new_n209), .A4(new_n536), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n892), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  OR4_X1    g702(.A1(KEYINPUT121), .A2(new_n899), .A3(new_n430), .A4(new_n897), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT121), .B1(new_n896), .B2(new_n897), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n723), .B(new_n870), .C1(new_n876), .C2(new_n890), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n907), .B2(G141gat), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n902), .A2(new_n903), .B1(new_n906), .B2(new_n908), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n211), .A2(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n900), .B2(new_n725), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n891), .A2(KEYINPUT59), .A3(new_n665), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n211), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n841), .B2(new_n879), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n666), .A2(new_n537), .A3(new_n672), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n838), .A2(new_n822), .A3(new_n821), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n887), .B2(new_n700), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n918), .B2(new_n620), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT125), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n916), .B(new_n921), .C1(new_n918), .C2(new_n620), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n286), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n877), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n875), .A2(KEYINPUT124), .A3(new_n878), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n915), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n870), .A2(KEYINPUT123), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n870), .A2(KEYINPUT123), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n725), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT59), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n911), .B1(new_n913), .B2(new_n931), .ZN(G1345gat));
  OAI21_X1  g731(.A(G155gat), .B1(new_n891), .B2(new_n699), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n900), .A2(new_n204), .A3(new_n620), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n891), .B2(new_n700), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n860), .A2(new_n205), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n899), .B2(new_n937), .ZN(G1347gat));
  NAND2_X1  g737(.A1(new_n675), .A2(new_n430), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n693), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n846), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(new_n338), .A3(new_n537), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n875), .A2(new_n430), .A3(new_n843), .A4(new_n675), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n723), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n942), .B1(new_n946), .B2(new_n338), .ZN(G1348gat));
  AOI211_X1 g746(.A(new_n665), .B(new_n941), .C1(new_n352), .C2(new_n353), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n725), .A3(new_n945), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n339), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n941), .B2(new_n699), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n620), .A2(new_n331), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n943), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT60), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n951), .B(new_n955), .C1(new_n943), .C2(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1350gat));
  NAND4_X1  g756(.A1(new_n875), .A2(new_n432), .A3(new_n701), .A4(new_n940), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G190gat), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(KEYINPUT61), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n944), .A2(new_n332), .A3(new_n701), .A4(new_n945), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n962), .B(new_n963), .C1(KEYINPUT61), .C2(new_n961), .ZN(G1351gat));
  NOR2_X1   g763(.A1(new_n841), .A2(new_n676), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n894), .A2(new_n396), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n723), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n734), .A2(new_n939), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n926), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n536), .A2(G197gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1352gat));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n725), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G204gat), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n665), .A2(G204gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n965), .A2(new_n966), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  NAND2_X1  g777(.A1(new_n975), .A2(new_n978), .ZN(G1353gat));
  OR3_X1    g778(.A1(new_n967), .A2(new_n227), .A3(new_n699), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n926), .A2(new_n620), .A3(new_n970), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  AOI21_X1  g783(.A(G218gat), .B1(new_n968), .B2(new_n701), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n701), .A2(new_n228), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n971), .B2(new_n986), .ZN(G1355gat));
endmodule


